magic
tech sky130A
magscale 1 2
timestamp 1606473343
<< locali >>
rect 7573 17731 7607 17901
rect 9505 17799 9539 18105
rect 9505 12087 9539 12189
rect 9413 7735 9447 7837
rect 9505 7803 9539 8041
rect 9505 6715 9539 6953
rect 13461 6103 13495 6341
rect 9137 2839 9171 2941
rect 9781 1547 9815 1989
<< viali >>
rect 9505 18105 9539 18139
rect 7573 17901 7607 17935
rect 9505 17765 9539 17799
rect 7573 17697 7607 17731
rect 11897 17289 11931 17323
rect 12817 17289 12851 17323
rect 5089 17153 5123 17187
rect 6285 17153 6319 17187
rect 7849 17153 7883 17187
rect 8953 17153 8987 17187
rect 10241 17153 10275 17187
rect 10425 17153 10459 17187
rect 13553 17153 13587 17187
rect 13829 17153 13863 17187
rect 1869 17085 1903 17119
rect 2789 17085 2823 17119
rect 8861 17085 8895 17119
rect 10977 17085 11011 17119
rect 11713 17085 11747 17119
rect 12633 17085 12667 17119
rect 2145 17017 2179 17051
rect 3065 17017 3099 17051
rect 4905 17017 4939 17051
rect 6009 17017 6043 17051
rect 7573 17017 7607 17051
rect 7665 17017 7699 17051
rect 8769 17017 8803 17051
rect 13645 17017 13679 17051
rect 4445 16949 4479 16983
rect 4813 16949 4847 16983
rect 5641 16949 5675 16983
rect 6101 16949 6135 16983
rect 7205 16949 7239 16983
rect 8401 16949 8435 16983
rect 9781 16949 9815 16983
rect 10149 16949 10183 16983
rect 11161 16949 11195 16983
rect 6929 16745 6963 16779
rect 7297 16745 7331 16779
rect 8585 16745 8619 16779
rect 11069 16745 11103 16779
rect 11805 16745 11839 16779
rect 12541 16745 12575 16779
rect 13277 16745 13311 16779
rect 1593 16609 1627 16643
rect 1869 16609 1903 16643
rect 2513 16609 2547 16643
rect 2789 16609 2823 16643
rect 3617 16609 3651 16643
rect 4353 16609 4387 16643
rect 4620 16609 4654 16643
rect 6193 16609 6227 16643
rect 7389 16609 7423 16643
rect 8493 16609 8527 16643
rect 10057 16609 10091 16643
rect 10885 16609 10919 16643
rect 11621 16609 11655 16643
rect 12357 16609 12391 16643
rect 13093 16609 13127 16643
rect 13829 16609 13863 16643
rect 7573 16541 7607 16575
rect 8769 16541 8803 16575
rect 10149 16541 10183 16575
rect 10333 16541 10367 16575
rect 14565 16541 14599 16575
rect 3433 16473 3467 16507
rect 6377 16473 6411 16507
rect 5733 16405 5767 16439
rect 8125 16405 8159 16439
rect 9689 16405 9723 16439
rect 14013 16405 14047 16439
rect 1593 16201 1627 16235
rect 3157 16201 3191 16235
rect 6929 16201 6963 16235
rect 4353 16133 4387 16167
rect 8309 16133 8343 16167
rect 11805 16133 11839 16167
rect 13829 16133 13863 16167
rect 2513 16065 2547 16099
rect 3617 16065 3651 16099
rect 3801 16065 3835 16099
rect 4813 16065 4847 16099
rect 4997 16065 5031 16099
rect 6193 16065 6227 16099
rect 7573 16065 7607 16099
rect 9781 16065 9815 16099
rect 10977 16065 11011 16099
rect 14933 16065 14967 16099
rect 1409 15997 1443 16031
rect 2237 15997 2271 16031
rect 6009 15997 6043 16031
rect 8125 15997 8159 16031
rect 9597 15997 9631 16031
rect 11621 15997 11655 16031
rect 12449 15997 12483 16031
rect 12817 15997 12851 16031
rect 13645 15997 13679 16031
rect 14657 15997 14691 16031
rect 5917 15929 5951 15963
rect 10885 15929 10919 15963
rect 13277 15929 13311 15963
rect 3525 15861 3559 15895
rect 4721 15861 4755 15895
rect 5549 15861 5583 15895
rect 7297 15861 7331 15895
rect 7389 15861 7423 15895
rect 9229 15861 9263 15895
rect 9689 15861 9723 15895
rect 10425 15861 10459 15895
rect 10793 15861 10827 15895
rect 12909 15861 12943 15895
rect 3157 15657 3191 15691
rect 5365 15657 5399 15691
rect 6929 15657 6963 15691
rect 8125 15657 8159 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 13461 15657 13495 15691
rect 14197 15657 14231 15691
rect 11345 15589 11379 15623
rect 1869 15521 1903 15555
rect 3249 15521 3283 15555
rect 4537 15521 4571 15555
rect 4629 15521 4663 15555
rect 5733 15521 5767 15555
rect 7021 15521 7055 15555
rect 8217 15521 8251 15555
rect 10057 15521 10091 15555
rect 11253 15521 11287 15555
rect 12449 15521 12483 15555
rect 13277 15521 13311 15555
rect 14013 15521 14047 15555
rect 2145 15453 2179 15487
rect 3433 15453 3467 15487
rect 4813 15453 4847 15487
rect 5825 15453 5859 15487
rect 6009 15453 6043 15487
rect 7205 15453 7239 15487
rect 8309 15453 8343 15487
rect 8953 15453 8987 15487
rect 10241 15453 10275 15487
rect 11437 15453 11471 15487
rect 12541 15453 12575 15487
rect 12633 15453 12667 15487
rect 7757 15385 7791 15419
rect 2789 15317 2823 15351
rect 4169 15317 4203 15351
rect 6561 15317 6595 15351
rect 10885 15317 10919 15351
rect 12081 15317 12115 15351
rect 6837 15113 6871 15147
rect 13369 15113 13403 15147
rect 3157 15045 3191 15079
rect 9873 15045 9907 15079
rect 12633 15045 12667 15079
rect 14105 15045 14139 15079
rect 2605 14977 2639 15011
rect 3801 14977 3835 15011
rect 4997 14977 5031 15011
rect 6009 14977 6043 15011
rect 6101 14977 6135 15011
rect 7481 14977 7515 15011
rect 9229 14977 9263 15011
rect 10333 14977 10367 15011
rect 10425 14977 10459 15011
rect 5917 14909 5951 14943
rect 7205 14909 7239 14943
rect 11069 14909 11103 14943
rect 12449 14909 12483 14943
rect 13185 14909 13219 14943
rect 13921 14909 13955 14943
rect 2421 14841 2455 14875
rect 3617 14841 3651 14875
rect 4721 14841 4755 14875
rect 1961 14773 1995 14807
rect 2329 14773 2363 14807
rect 3525 14773 3559 14807
rect 4353 14773 4387 14807
rect 4813 14773 4847 14807
rect 5549 14773 5583 14807
rect 7297 14773 7331 14807
rect 8033 14773 8067 14807
rect 8677 14773 8711 14807
rect 9045 14773 9079 14807
rect 9137 14773 9171 14807
rect 10241 14773 10275 14807
rect 11253 14773 11287 14807
rect 1593 14569 1627 14603
rect 4169 14569 4203 14603
rect 4537 14569 4571 14603
rect 12081 14569 12115 14603
rect 13277 14569 13311 14603
rect 1961 14501 1995 14535
rect 12541 14501 12575 14535
rect 13645 14501 13679 14535
rect 3157 14433 3191 14467
rect 4629 14433 4663 14467
rect 5632 14433 5666 14467
rect 7472 14433 7506 14467
rect 9229 14433 9263 14467
rect 10057 14433 10091 14467
rect 11253 14433 11287 14467
rect 12449 14433 12483 14467
rect 13737 14433 13771 14467
rect 2053 14365 2087 14399
rect 2145 14365 2179 14399
rect 3249 14365 3283 14399
rect 3433 14365 3467 14399
rect 4813 14365 4847 14399
rect 5365 14365 5399 14399
rect 7205 14365 7239 14399
rect 10149 14365 10183 14399
rect 10241 14365 10275 14399
rect 11345 14365 11379 14399
rect 11529 14365 11563 14399
rect 12633 14365 12667 14399
rect 13829 14365 13863 14399
rect 8585 14297 8619 14331
rect 9689 14297 9723 14331
rect 2789 14229 2823 14263
rect 6745 14229 6779 14263
rect 9045 14229 9079 14263
rect 10885 14229 10919 14263
rect 2513 14025 2547 14059
rect 10517 14025 10551 14059
rect 11713 14025 11747 14059
rect 3709 13957 3743 13991
rect 6285 13957 6319 13991
rect 8217 13957 8251 13991
rect 10057 13957 10091 13991
rect 3157 13889 3191 13923
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 8677 13889 8711 13923
rect 11161 13889 11195 13923
rect 13001 13889 13035 13923
rect 1593 13821 1627 13855
rect 1869 13821 1903 13855
rect 2973 13821 3007 13855
rect 4905 13821 4939 13855
rect 6837 13821 6871 13855
rect 11897 13821 11931 13855
rect 12817 13821 12851 13855
rect 12909 13821 12943 13855
rect 13956 13821 13990 13855
rect 5172 13753 5206 13787
rect 7104 13753 7138 13787
rect 8922 13753 8956 13787
rect 2881 13685 2915 13719
rect 4077 13685 4111 13719
rect 10885 13685 10919 13719
rect 10977 13685 11011 13719
rect 12449 13685 12483 13719
rect 14059 13685 14093 13719
rect 1961 13481 1995 13515
rect 3249 13481 3283 13515
rect 6377 13481 6411 13515
rect 8217 13481 8251 13515
rect 11897 13481 11931 13515
rect 12725 13481 12759 13515
rect 2053 13413 2087 13447
rect 13829 13413 13863 13447
rect 3157 13345 3191 13379
rect 4077 13345 4111 13379
rect 5253 13345 5287 13379
rect 7104 13345 7138 13379
rect 8677 13345 8711 13379
rect 9689 13345 9723 13379
rect 9945 13345 9979 13379
rect 11989 13345 12023 13379
rect 12909 13345 12943 13379
rect 2145 13277 2179 13311
rect 3433 13277 3467 13311
rect 4261 13277 4295 13311
rect 4997 13277 5031 13311
rect 6837 13277 6871 13311
rect 8861 13277 8895 13311
rect 12081 13277 12115 13311
rect 13737 13277 13771 13311
rect 14013 13277 14047 13311
rect 1593 13209 1627 13243
rect 2789 13209 2823 13243
rect 11069 13209 11103 13243
rect 11529 13141 11563 13175
rect 1869 12937 1903 12971
rect 4445 12937 4479 12971
rect 6837 12937 6871 12971
rect 10609 12937 10643 12971
rect 13645 12937 13679 12971
rect 12449 12869 12483 12903
rect 2513 12801 2547 12835
rect 3065 12801 3099 12835
rect 4905 12801 4939 12835
rect 7481 12801 7515 12835
rect 9045 12801 9079 12835
rect 11161 12801 11195 12835
rect 12909 12801 12943 12835
rect 13001 12801 13035 12835
rect 14197 12801 14231 12835
rect 5161 12733 5195 12767
rect 7205 12733 7239 12767
rect 8309 12733 8343 12767
rect 8401 12733 8435 12767
rect 10517 12733 10551 12767
rect 10977 12733 11011 12767
rect 11989 12733 12023 12767
rect 12817 12733 12851 12767
rect 3332 12665 3366 12699
rect 7297 12665 7331 12699
rect 11069 12665 11103 12699
rect 14105 12665 14139 12699
rect 2237 12597 2271 12631
rect 2329 12597 2363 12631
rect 6285 12597 6319 12631
rect 8125 12597 8159 12631
rect 9689 12597 9723 12631
rect 10333 12597 10367 12631
rect 11805 12597 11839 12631
rect 14013 12597 14047 12631
rect 1685 12393 1719 12427
rect 2053 12393 2087 12427
rect 6101 12393 6135 12427
rect 6561 12393 6595 12427
rect 7481 12393 7515 12427
rect 8769 12393 8803 12427
rect 9689 12393 9723 12427
rect 10885 12393 10919 12427
rect 11253 12393 11287 12427
rect 4077 12325 4111 12359
rect 4353 12325 4387 12359
rect 8677 12325 8711 12359
rect 13645 12325 13679 12359
rect 2697 12257 2731 12291
rect 4721 12257 4755 12291
rect 4988 12257 5022 12291
rect 6745 12257 6779 12291
rect 10425 12257 10459 12291
rect 10793 12257 10827 12291
rect 11345 12257 11379 12291
rect 12449 12257 12483 12291
rect 12541 12257 12575 12291
rect 2145 12189 2179 12223
rect 2329 12189 2363 12223
rect 3341 12189 3375 12223
rect 7573 12189 7607 12223
rect 7757 12189 7791 12223
rect 8953 12189 8987 12223
rect 9505 12189 9539 12223
rect 11437 12189 11471 12223
rect 12633 12189 12667 12223
rect 13737 12189 13771 12223
rect 13829 12189 13863 12223
rect 7113 12121 7147 12155
rect 10241 12121 10275 12155
rect 13277 12121 13311 12155
rect 8309 12053 8343 12087
rect 9505 12053 9539 12087
rect 12081 12053 12115 12087
rect 4445 11849 4479 11883
rect 12449 11849 12483 11883
rect 2513 11713 2547 11747
rect 3065 11713 3099 11747
rect 4905 11713 4939 11747
rect 6837 11713 6871 11747
rect 11069 11713 11103 11747
rect 13001 11713 13035 11747
rect 14197 11713 14231 11747
rect 3332 11645 3366 11679
rect 7093 11645 7127 11679
rect 8677 11645 8711 11679
rect 8933 11645 8967 11679
rect 10885 11645 10919 11679
rect 12817 11645 12851 11679
rect 14841 11645 14875 11679
rect 2329 11577 2363 11611
rect 5172 11577 5206 11611
rect 11713 11577 11747 11611
rect 12909 11577 12943 11611
rect 14013 11577 14047 11611
rect 1869 11509 1903 11543
rect 2237 11509 2271 11543
rect 6285 11509 6319 11543
rect 8217 11509 8251 11543
rect 10057 11509 10091 11543
rect 10517 11509 10551 11543
rect 10977 11509 11011 11543
rect 13645 11509 13679 11543
rect 14105 11509 14139 11543
rect 15025 11509 15059 11543
rect 11529 11305 11563 11339
rect 11989 11305 12023 11339
rect 12725 11305 12759 11339
rect 13921 11305 13955 11339
rect 1869 11237 1903 11271
rect 6285 11237 6319 11271
rect 7196 11237 7230 11271
rect 9934 11237 9968 11271
rect 14381 11237 14415 11271
rect 1593 11169 1627 11203
rect 2145 11169 2179 11203
rect 2412 11169 2446 11203
rect 4077 11169 4111 11203
rect 4344 11169 4378 11203
rect 6101 11169 6135 11203
rect 11897 11169 11931 11203
rect 13093 11169 13127 11203
rect 14289 11169 14323 11203
rect 6929 11101 6963 11135
rect 8769 11101 8803 11135
rect 9689 11101 9723 11135
rect 12081 11101 12115 11135
rect 13185 11101 13219 11135
rect 13277 11101 13311 11135
rect 14565 11101 14599 11135
rect 3525 11033 3559 11067
rect 5457 11033 5491 11067
rect 5917 11033 5951 11067
rect 8309 11033 8343 11067
rect 11069 11033 11103 11067
rect 1593 10761 1627 10795
rect 1869 10761 1903 10795
rect 6285 10761 6319 10795
rect 13645 10761 13679 10795
rect 8217 10693 8251 10727
rect 11897 10693 11931 10727
rect 2513 10625 2547 10659
rect 4905 10625 4939 10659
rect 6837 10625 6871 10659
rect 10517 10625 10551 10659
rect 13001 10625 13035 10659
rect 14197 10625 14231 10659
rect 1409 10557 1443 10591
rect 3065 10557 3099 10591
rect 7104 10557 7138 10591
rect 8677 10557 8711 10591
rect 12817 10557 12851 10591
rect 12909 10557 12943 10591
rect 14841 10557 14875 10591
rect 2329 10489 2363 10523
rect 3332 10489 3366 10523
rect 5150 10489 5184 10523
rect 8922 10489 8956 10523
rect 10784 10489 10818 10523
rect 2237 10421 2271 10455
rect 4445 10421 4479 10455
rect 10057 10421 10091 10455
rect 12449 10421 12483 10455
rect 14013 10421 14047 10455
rect 14105 10421 14139 10455
rect 15025 10421 15059 10455
rect 7297 10217 7331 10251
rect 9137 10217 9171 10251
rect 11897 10217 11931 10251
rect 13185 10217 13219 10251
rect 13921 10217 13955 10251
rect 2412 10149 2446 10183
rect 6184 10149 6218 10183
rect 8002 10149 8036 10183
rect 14289 10149 14323 10183
rect 1409 10081 1443 10115
rect 2145 10081 2179 10115
rect 4077 10081 4111 10115
rect 4344 10081 4378 10115
rect 7757 10081 7791 10115
rect 9945 10081 9979 10115
rect 13093 10081 13127 10115
rect 5917 10013 5951 10047
rect 9689 10013 9723 10047
rect 11989 10013 12023 10047
rect 12081 10013 12115 10047
rect 13277 10013 13311 10047
rect 14381 10013 14415 10047
rect 14473 10013 14507 10047
rect 5457 9945 5491 9979
rect 11069 9945 11103 9979
rect 12725 9945 12759 9979
rect 1593 9877 1627 9911
rect 3525 9877 3559 9911
rect 11529 9877 11563 9911
rect 1869 9673 1903 9707
rect 4445 9673 4479 9707
rect 12449 9673 12483 9707
rect 15025 9673 15059 9707
rect 4997 9605 5031 9639
rect 10425 9605 10459 9639
rect 2513 9537 2547 9571
rect 5273 9537 5307 9571
rect 13093 9537 13127 9571
rect 14197 9537 14231 9571
rect 3065 9469 3099 9503
rect 5181 9469 5215 9503
rect 8769 9469 8803 9503
rect 9045 9469 9079 9503
rect 10517 9469 10551 9503
rect 12817 9469 12851 9503
rect 12909 9469 12943 9503
rect 14841 9469 14875 9503
rect 2237 9401 2271 9435
rect 3332 9401 3366 9435
rect 5540 9401 5574 9435
rect 7205 9401 7239 9435
rect 9312 9401 9346 9435
rect 10784 9401 10818 9435
rect 14105 9401 14139 9435
rect 2329 9333 2363 9367
rect 6653 9333 6687 9367
rect 11897 9333 11931 9367
rect 13645 9333 13679 9367
rect 14013 9333 14047 9367
rect 13829 9129 13863 9163
rect 9934 9061 9968 9095
rect 1409 8993 1443 9027
rect 2145 8993 2179 9027
rect 2412 8993 2446 9027
rect 4528 8993 4562 9027
rect 5733 8993 5767 9027
rect 6000 8993 6034 9027
rect 7573 8993 7607 9027
rect 7840 8993 7874 9027
rect 11785 8993 11819 9027
rect 13737 8993 13771 9027
rect 4261 8925 4295 8959
rect 9689 8925 9723 8959
rect 11529 8925 11563 8959
rect 13921 8925 13955 8959
rect 14565 8925 14599 8959
rect 3525 8857 3559 8891
rect 5641 8857 5675 8891
rect 8953 8857 8987 8891
rect 13369 8857 13403 8891
rect 1593 8789 1627 8823
rect 7113 8789 7147 8823
rect 11069 8789 11103 8823
rect 12909 8789 12943 8823
rect 8217 8585 8251 8619
rect 11897 8585 11931 8619
rect 12449 8585 12483 8619
rect 13645 8585 13679 8619
rect 4445 8517 4479 8551
rect 6285 8517 6319 8551
rect 10057 8517 10091 8551
rect 15025 8517 15059 8551
rect 2053 8449 2087 8483
rect 2237 8449 2271 8483
rect 3065 8449 3099 8483
rect 8677 8449 8711 8483
rect 13001 8449 13035 8483
rect 14289 8449 14323 8483
rect 1961 8381 1995 8415
rect 2973 8381 3007 8415
rect 4905 8381 4939 8415
rect 6837 8381 6871 8415
rect 8933 8381 8967 8415
rect 10517 8381 10551 8415
rect 12909 8381 12943 8415
rect 14841 8381 14875 8415
rect 3310 8313 3344 8347
rect 5172 8313 5206 8347
rect 7082 8313 7116 8347
rect 10762 8313 10796 8347
rect 12817 8313 12851 8347
rect 14105 8313 14139 8347
rect 1593 8245 1627 8279
rect 2789 8245 2823 8279
rect 14013 8245 14047 8279
rect 4905 8041 4939 8075
rect 7113 8041 7147 8075
rect 7941 8041 7975 8075
rect 8033 8041 8067 8075
rect 8769 8041 8803 8075
rect 9505 8041 9539 8075
rect 11529 8041 11563 8075
rect 11897 8041 11931 8075
rect 13921 8041 13955 8075
rect 6000 7973 6034 8007
rect 8677 7973 8711 8007
rect 9137 7973 9171 8007
rect 1409 7905 1443 7939
rect 2412 7905 2446 7939
rect 4997 7905 5031 7939
rect 2145 7837 2179 7871
rect 5181 7837 5215 7871
rect 5733 7837 5767 7871
rect 8861 7837 8895 7871
rect 9413 7837 9447 7871
rect 3525 7769 3559 7803
rect 14289 7973 14323 8007
rect 9689 7905 9723 7939
rect 9945 7905 9979 7939
rect 11989 7905 12023 7939
rect 13093 7905 13127 7939
rect 12081 7837 12115 7871
rect 13185 7837 13219 7871
rect 13277 7837 13311 7871
rect 14381 7837 14415 7871
rect 14473 7837 14507 7871
rect 9505 7769 9539 7803
rect 1593 7701 1627 7735
rect 4537 7701 4571 7735
rect 8309 7701 8343 7735
rect 9413 7701 9447 7735
rect 11069 7701 11103 7735
rect 12725 7701 12759 7735
rect 4445 7497 4479 7531
rect 12449 7497 12483 7531
rect 13645 7497 13679 7531
rect 1869 7429 1903 7463
rect 8217 7429 8251 7463
rect 2513 7361 2547 7395
rect 3065 7361 3099 7395
rect 4905 7361 4939 7395
rect 8677 7361 8711 7395
rect 11069 7361 11103 7395
rect 13001 7361 13035 7395
rect 14197 7361 14231 7395
rect 6844 7293 6878 7327
rect 8309 7293 8343 7327
rect 10977 7293 11011 7327
rect 12817 7293 12851 7327
rect 14841 7293 14875 7327
rect 3332 7225 3366 7259
rect 5172 7225 5206 7259
rect 7104 7225 7138 7259
rect 8944 7225 8978 7259
rect 10885 7225 10919 7259
rect 14105 7225 14139 7259
rect 2237 7157 2271 7191
rect 2329 7157 2363 7191
rect 6285 7157 6319 7191
rect 10057 7157 10091 7191
rect 10517 7157 10551 7191
rect 11713 7157 11747 7191
rect 12909 7157 12943 7191
rect 14013 7157 14047 7191
rect 15025 7157 15059 7191
rect 7205 6953 7239 6987
rect 9505 6953 9539 6987
rect 10057 6953 10091 6987
rect 12449 6953 12483 6987
rect 14657 6953 14691 6987
rect 4905 6885 4939 6919
rect 1409 6817 1443 6851
rect 2145 6817 2179 6851
rect 2412 6817 2446 6851
rect 6081 6817 6115 6851
rect 7932 6817 7966 6851
rect 4997 6749 5031 6783
rect 5181 6749 5215 6783
rect 5825 6749 5859 6783
rect 7665 6749 7699 6783
rect 11253 6885 11287 6919
rect 10149 6817 10183 6851
rect 12541 6817 12575 6851
rect 13645 6817 13679 6851
rect 14473 6817 14507 6851
rect 10241 6749 10275 6783
rect 11345 6749 11379 6783
rect 11529 6749 11563 6783
rect 12633 6749 12667 6783
rect 13737 6749 13771 6783
rect 13921 6749 13955 6783
rect 3525 6681 3559 6715
rect 9045 6681 9079 6715
rect 9505 6681 9539 6715
rect 9689 6681 9723 6715
rect 1593 6613 1627 6647
rect 4537 6613 4571 6647
rect 10885 6613 10919 6647
rect 12081 6613 12115 6647
rect 13277 6613 13311 6647
rect 1869 6409 1903 6443
rect 4445 6409 4479 6443
rect 8217 6409 8251 6443
rect 10057 6409 10091 6443
rect 10517 6409 10551 6443
rect 12449 6409 12483 6443
rect 13461 6341 13495 6375
rect 2421 6273 2455 6307
rect 10977 6273 11011 6307
rect 11161 6273 11195 6307
rect 11713 6273 11747 6307
rect 13001 6273 13035 6307
rect 2237 6205 2271 6239
rect 3065 6205 3099 6239
rect 3321 6205 3355 6239
rect 4905 6205 4939 6239
rect 6837 6205 6871 6239
rect 7093 6205 7127 6239
rect 8677 6205 8711 6239
rect 12817 6205 12851 6239
rect 13277 6205 13311 6239
rect 5172 6137 5206 6171
rect 8922 6137 8956 6171
rect 14197 6273 14231 6307
rect 14841 6205 14875 6239
rect 14105 6137 14139 6171
rect 2329 6069 2363 6103
rect 6285 6069 6319 6103
rect 10885 6069 10919 6103
rect 12909 6069 12943 6103
rect 13461 6069 13495 6103
rect 13645 6069 13679 6103
rect 14013 6069 14047 6103
rect 15025 6069 15059 6103
rect 1409 5865 1443 5899
rect 3157 5865 3191 5899
rect 4905 5865 4939 5899
rect 9689 5865 9723 5899
rect 11253 5865 11287 5899
rect 14657 5865 14691 5899
rect 1777 5797 1811 5831
rect 2513 5797 2547 5831
rect 7932 5797 7966 5831
rect 10057 5797 10091 5831
rect 12449 5797 12483 5831
rect 13737 5797 13771 5831
rect 2237 5729 2271 5763
rect 3249 5729 3283 5763
rect 5989 5729 6023 5763
rect 10149 5729 10183 5763
rect 11345 5729 11379 5763
rect 13645 5729 13679 5763
rect 14473 5729 14507 5763
rect 1869 5661 1903 5695
rect 2053 5661 2087 5695
rect 3433 5661 3467 5695
rect 4997 5661 5031 5695
rect 5181 5661 5215 5695
rect 5733 5661 5767 5695
rect 7665 5661 7699 5695
rect 10333 5661 10367 5695
rect 11529 5661 11563 5695
rect 12541 5661 12575 5695
rect 12633 5661 12667 5695
rect 13829 5661 13863 5695
rect 4537 5593 4571 5627
rect 10885 5593 10919 5627
rect 2789 5525 2823 5559
rect 7113 5525 7147 5559
rect 9045 5525 9079 5559
rect 12081 5525 12115 5559
rect 13277 5525 13311 5559
rect 6285 5321 6319 5355
rect 9229 5321 9263 5355
rect 10425 5321 10459 5355
rect 11253 5321 11287 5355
rect 3525 5253 3559 5287
rect 8769 5253 8803 5287
rect 1869 5185 1903 5219
rect 1961 5185 1995 5219
rect 2973 5185 3007 5219
rect 3157 5185 3191 5219
rect 4353 5185 4387 5219
rect 7389 5185 7423 5219
rect 9781 5185 9815 5219
rect 10977 5185 11011 5219
rect 11897 5185 11931 5219
rect 13001 5185 13035 5219
rect 14197 5185 14231 5219
rect 3341 5117 3375 5151
rect 4905 5117 4939 5151
rect 10793 5117 10827 5151
rect 11713 5117 11747 5151
rect 12909 5117 12943 5151
rect 14013 5117 14047 5151
rect 14841 5117 14875 5151
rect 1777 5049 1811 5083
rect 2881 5049 2915 5083
rect 4077 5049 4111 5083
rect 5172 5049 5206 5083
rect 7656 5049 7690 5083
rect 9597 5049 9631 5083
rect 10885 5049 10919 5083
rect 12817 5049 12851 5083
rect 1409 4981 1443 5015
rect 2513 4981 2547 5015
rect 3709 4981 3743 5015
rect 4169 4981 4203 5015
rect 9689 4981 9723 5015
rect 11621 4981 11655 5015
rect 12449 4981 12483 5015
rect 13645 4981 13679 5015
rect 14105 4981 14139 5015
rect 15025 4981 15059 5015
rect 2789 4777 2823 4811
rect 3249 4777 3283 4811
rect 4537 4777 4571 4811
rect 5273 4777 5307 4811
rect 8309 4777 8343 4811
rect 8769 4777 8803 4811
rect 9689 4777 9723 4811
rect 11345 4777 11379 4811
rect 11897 4777 11931 4811
rect 13645 4777 13679 4811
rect 1676 4709 1710 4743
rect 4445 4709 4479 4743
rect 6736 4709 6770 4743
rect 8677 4709 8711 4743
rect 11253 4709 11287 4743
rect 12449 4709 12483 4743
rect 13737 4709 13771 4743
rect 5641 4641 5675 4675
rect 6469 4641 6503 4675
rect 10057 4641 10091 4675
rect 11713 4641 11747 4675
rect 14473 4641 14507 4675
rect 3341 4573 3375 4607
rect 3525 4573 3559 4607
rect 4629 4573 4663 4607
rect 5733 4573 5767 4607
rect 5917 4573 5951 4607
rect 8953 4573 8987 4607
rect 10149 4573 10183 4607
rect 10241 4573 10275 4607
rect 11529 4573 11563 4607
rect 12541 4573 12575 4607
rect 12633 4573 12667 4607
rect 13829 4573 13863 4607
rect 2881 4505 2915 4539
rect 10885 4505 10919 4539
rect 4077 4437 4111 4471
rect 7849 4437 7883 4471
rect 12081 4437 12115 4471
rect 13277 4437 13311 4471
rect 14657 4437 14691 4471
rect 3985 4233 4019 4267
rect 5549 4233 5583 4267
rect 6837 4233 6871 4267
rect 4077 4165 4111 4199
rect 8861 4165 8895 4199
rect 11253 4165 11287 4199
rect 12449 4165 12483 4199
rect 13645 4165 13679 4199
rect 2237 4097 2271 4131
rect 4721 4097 4755 4131
rect 6193 4097 6227 4131
rect 7389 4097 7423 4131
rect 8585 4097 8619 4131
rect 9321 4097 9355 4131
rect 9505 4097 9539 4131
rect 10977 4097 11011 4131
rect 11851 4097 11885 4131
rect 13001 4097 13035 4131
rect 14197 4097 14231 4131
rect 2605 4029 2639 4063
rect 4905 4029 4939 4063
rect 8493 4029 8527 4063
rect 10241 4029 10275 4063
rect 10793 4029 10827 4063
rect 11621 4029 11655 4063
rect 14841 4029 14875 4063
rect 2850 3961 2884 3995
rect 5181 3961 5215 3995
rect 5917 3961 5951 3995
rect 6009 3961 6043 3995
rect 7297 3961 7331 3995
rect 8401 3961 8435 3995
rect 9229 3961 9263 3995
rect 10885 3961 10919 3995
rect 11713 3961 11747 3995
rect 13553 3961 13587 3995
rect 14013 3961 14047 3995
rect 14105 3961 14139 3995
rect 1593 3893 1627 3927
rect 1961 3893 1995 3927
rect 2053 3893 2087 3927
rect 4445 3893 4479 3927
rect 4537 3893 4571 3927
rect 7205 3893 7239 3927
rect 8033 3893 8067 3927
rect 10057 3893 10091 3927
rect 10425 3893 10459 3927
rect 12817 3893 12851 3927
rect 12909 3893 12943 3927
rect 15025 3893 15059 3927
rect 1869 3689 1903 3723
rect 2881 3689 2915 3723
rect 4445 3689 4479 3723
rect 6193 3689 6227 3723
rect 7389 3689 7423 3723
rect 8217 3689 8251 3723
rect 13277 3689 13311 3723
rect 13737 3689 13771 3723
rect 4537 3621 4571 3655
rect 6561 3621 6595 3655
rect 7757 3621 7791 3655
rect 8677 3621 8711 3655
rect 10149 3621 10183 3655
rect 11253 3621 11287 3655
rect 12449 3621 12483 3655
rect 12541 3621 12575 3655
rect 1777 3553 1811 3587
rect 2789 3553 2823 3587
rect 3249 3553 3283 3587
rect 3341 3553 3375 3587
rect 5365 3553 5399 3587
rect 5457 3553 5491 3587
rect 7849 3553 7883 3587
rect 8585 3553 8619 3587
rect 9045 3553 9079 3587
rect 10057 3553 10091 3587
rect 11345 3553 11379 3587
rect 11713 3553 11747 3587
rect 13645 3553 13679 3587
rect 14473 3553 14507 3587
rect 2053 3485 2087 3519
rect 3525 3485 3559 3519
rect 4721 3485 4755 3519
rect 5641 3485 5675 3519
rect 6653 3485 6687 3519
rect 6837 3485 6871 3519
rect 7941 3485 7975 3519
rect 8861 3485 8895 3519
rect 9229 3485 9263 3519
rect 10333 3485 10367 3519
rect 11437 3485 11471 3519
rect 12633 3485 12667 3519
rect 13921 3485 13955 3519
rect 1409 3417 1443 3451
rect 4997 3417 5031 3451
rect 10885 3417 10919 3451
rect 4077 3349 4111 3383
rect 9689 3349 9723 3383
rect 11897 3349 11931 3383
rect 12081 3349 12115 3383
rect 14657 3349 14691 3383
rect 2789 3145 2823 3179
rect 5549 3145 5583 3179
rect 6837 3145 6871 3179
rect 7665 3145 7699 3179
rect 9229 3145 9263 3179
rect 11253 3145 11287 3179
rect 13277 3145 13311 3179
rect 4353 3077 4387 3111
rect 8861 3077 8895 3111
rect 10241 3077 10275 3111
rect 2881 3009 2915 3043
rect 4997 3009 5031 3043
rect 6009 3009 6043 3043
rect 6193 3009 6227 3043
rect 7297 3009 7331 3043
rect 7481 3009 7515 3043
rect 8125 3009 8159 3043
rect 8309 3009 8343 3043
rect 9781 3009 9815 3043
rect 10977 3009 11011 3043
rect 11805 3009 11839 3043
rect 13001 3009 13035 3043
rect 13829 3009 13863 3043
rect 14381 3009 14415 3043
rect 3148 2941 3182 2975
rect 4721 2941 4755 2975
rect 4813 2941 4847 2975
rect 5917 2941 5951 2975
rect 7205 2941 7239 2975
rect 9045 2941 9079 2975
rect 9137 2941 9171 2975
rect 9597 2941 9631 2975
rect 9689 2941 9723 2975
rect 10057 2941 10091 2975
rect 10793 2941 10827 2975
rect 11621 2941 11655 2975
rect 11713 2941 11747 2975
rect 14105 2941 14139 2975
rect 14657 2941 14691 2975
rect 1676 2873 1710 2907
rect 12817 2873 12851 2907
rect 13737 2873 13771 2907
rect 4261 2805 4295 2839
rect 8033 2805 8067 2839
rect 9137 2805 9171 2839
rect 10425 2805 10459 2839
rect 10885 2805 10919 2839
rect 12449 2805 12483 2839
rect 12909 2805 12943 2839
rect 13645 2805 13679 2839
rect 14841 2805 14875 2839
rect 2881 2601 2915 2635
rect 3249 2601 3283 2635
rect 5457 2601 5491 2635
rect 5917 2601 5951 2635
rect 6929 2601 6963 2635
rect 8585 2601 8619 2635
rect 8677 2601 8711 2635
rect 10241 2601 10275 2635
rect 11437 2601 11471 2635
rect 12633 2601 12667 2635
rect 13921 2601 13955 2635
rect 6561 2533 6595 2567
rect 7297 2533 7331 2567
rect 10149 2533 10183 2567
rect 11345 2533 11379 2567
rect 15117 2533 15151 2567
rect 1409 2465 1443 2499
rect 1676 2465 1710 2499
rect 4629 2465 4663 2499
rect 4721 2465 4755 2499
rect 5825 2465 5859 2499
rect 6285 2465 6319 2499
rect 11989 2465 12023 2499
rect 13001 2465 13035 2499
rect 13829 2465 13863 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 3341 2397 3375 2431
rect 3525 2397 3559 2431
rect 4905 2397 4939 2431
rect 6101 2397 6135 2431
rect 7389 2397 7423 2431
rect 7481 2397 7515 2431
rect 8861 2397 8895 2431
rect 10333 2397 10367 2431
rect 11529 2397 11563 2431
rect 12173 2397 12207 2431
rect 13093 2397 13127 2431
rect 13277 2397 13311 2431
rect 14105 2397 14139 2431
rect 14473 2397 14507 2431
rect 8217 2329 8251 2363
rect 13461 2329 13495 2363
rect 2789 2261 2823 2295
rect 4261 2261 4295 2295
rect 9781 2261 9815 2295
rect 10977 2261 11011 2295
rect 9781 1989 9815 2023
rect 9781 1513 9815 1547
<< metal1 >>
rect 566 18368 572 18420
rect 624 18408 630 18420
rect 9122 18408 9128 18420
rect 624 18380 9128 18408
rect 624 18368 630 18380
rect 9122 18368 9128 18380
rect 9180 18368 9186 18420
rect 8202 18164 8208 18216
rect 8260 18204 8266 18216
rect 8754 18204 8760 18216
rect 8260 18176 8760 18204
rect 8260 18164 8266 18176
rect 8754 18164 8760 18176
rect 8812 18164 8818 18216
rect 1762 18096 1768 18148
rect 1820 18136 1826 18148
rect 9493 18139 9551 18145
rect 9493 18136 9505 18139
rect 1820 18108 9505 18136
rect 1820 18096 1826 18108
rect 9493 18105 9505 18108
rect 9539 18105 9551 18139
rect 9493 18099 9551 18105
rect 9674 18096 9680 18148
rect 9732 18136 9738 18148
rect 11054 18136 11060 18148
rect 9732 18108 11060 18136
rect 9732 18096 9738 18108
rect 11054 18096 11060 18108
rect 11112 18096 11118 18148
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 10594 18068 10600 18080
rect 7524 18040 10600 18068
rect 7524 18028 7530 18040
rect 10594 18028 10600 18040
rect 10652 18028 10658 18080
rect 4062 17960 4068 18012
rect 4120 18000 4126 18012
rect 12986 18000 12992 18012
rect 4120 17972 12992 18000
rect 4120 17960 4126 17972
rect 12986 17960 12992 17972
rect 13044 17960 13050 18012
rect 7561 17935 7619 17941
rect 7561 17901 7573 17935
rect 7607 17932 7619 17935
rect 12802 17932 12808 17944
rect 7607 17904 12808 17932
rect 7607 17901 7619 17904
rect 7561 17895 7619 17901
rect 12802 17892 12808 17904
rect 12860 17892 12866 17944
rect 7834 17824 7840 17876
rect 7892 17864 7898 17876
rect 12618 17864 12624 17876
rect 7892 17836 12624 17864
rect 7892 17824 7898 17836
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 3418 17756 3424 17808
rect 3476 17796 3482 17808
rect 9398 17796 9404 17808
rect 3476 17768 9404 17796
rect 3476 17756 3482 17768
rect 9398 17756 9404 17768
rect 9456 17756 9462 17808
rect 9493 17799 9551 17805
rect 9493 17765 9505 17799
rect 9539 17796 9551 17799
rect 12526 17796 12532 17808
rect 9539 17768 12532 17796
rect 9539 17765 9551 17768
rect 9493 17759 9551 17765
rect 12526 17756 12532 17768
rect 12584 17756 12590 17808
rect 2222 17688 2228 17740
rect 2280 17728 2286 17740
rect 7561 17731 7619 17737
rect 7561 17728 7573 17731
rect 2280 17700 7573 17728
rect 2280 17688 2286 17700
rect 7561 17697 7573 17700
rect 7607 17697 7619 17731
rect 7561 17691 7619 17697
rect 8294 17688 8300 17740
rect 8352 17728 8358 17740
rect 8938 17728 8944 17740
rect 8352 17700 8944 17728
rect 8352 17688 8358 17700
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 7006 17620 7012 17672
rect 7064 17660 7070 17672
rect 12158 17660 12164 17672
rect 7064 17632 12164 17660
rect 7064 17620 7070 17632
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 13538 17620 13544 17672
rect 13596 17660 13602 17672
rect 14458 17660 14464 17672
rect 13596 17632 14464 17660
rect 13596 17620 13602 17632
rect 14458 17620 14464 17632
rect 14516 17620 14522 17672
rect 1302 17552 1308 17604
rect 1360 17592 1366 17604
rect 5442 17592 5448 17604
rect 1360 17564 5448 17592
rect 1360 17552 1366 17564
rect 5442 17552 5448 17564
rect 5500 17552 5506 17604
rect 8662 17552 8668 17604
rect 8720 17592 8726 17604
rect 15194 17592 15200 17604
rect 8720 17564 15200 17592
rect 8720 17552 8726 17564
rect 15194 17552 15200 17564
rect 15252 17592 15258 17604
rect 15930 17592 15936 17604
rect 15252 17564 15936 17592
rect 15252 17552 15258 17564
rect 15930 17552 15936 17564
rect 15988 17552 15994 17604
rect 1394 17484 1400 17536
rect 1452 17524 1458 17536
rect 7282 17524 7288 17536
rect 1452 17496 7288 17524
rect 1452 17484 1458 17496
rect 7282 17484 7288 17496
rect 7340 17484 7346 17536
rect 7558 17484 7564 17536
rect 7616 17524 7622 17536
rect 10318 17524 10324 17536
rect 7616 17496 10324 17524
rect 7616 17484 7622 17496
rect 10318 17484 10324 17496
rect 10376 17484 10382 17536
rect 10778 17484 10784 17536
rect 10836 17524 10842 17536
rect 11238 17524 11244 17536
rect 10836 17496 11244 17524
rect 10836 17484 10842 17496
rect 11238 17484 11244 17496
rect 11296 17484 11302 17536
rect 1104 17434 15824 17456
rect 1104 17382 3447 17434
rect 3499 17382 3511 17434
rect 3563 17382 3575 17434
rect 3627 17382 3639 17434
rect 3691 17382 8378 17434
rect 8430 17382 8442 17434
rect 8494 17382 8506 17434
rect 8558 17382 8570 17434
rect 8622 17382 13308 17434
rect 13360 17382 13372 17434
rect 13424 17382 13436 17434
rect 13488 17382 13500 17434
rect 13552 17382 15824 17434
rect 1104 17360 15824 17382
rect 7282 17280 7288 17332
rect 7340 17320 7346 17332
rect 10778 17320 10784 17332
rect 7340 17292 10784 17320
rect 7340 17280 7346 17292
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 11238 17280 11244 17332
rect 11296 17320 11302 17332
rect 11885 17323 11943 17329
rect 11885 17320 11897 17323
rect 11296 17292 11897 17320
rect 11296 17280 11302 17292
rect 11885 17289 11897 17292
rect 11931 17289 11943 17323
rect 11885 17283 11943 17289
rect 12618 17280 12624 17332
rect 12676 17320 12682 17332
rect 12805 17323 12863 17329
rect 12805 17320 12817 17323
rect 12676 17292 12817 17320
rect 12676 17280 12682 17292
rect 12805 17289 12817 17292
rect 12851 17289 12863 17323
rect 12805 17283 12863 17289
rect 5534 17252 5540 17264
rect 5000 17224 5540 17252
rect 3602 17144 3608 17196
rect 3660 17184 3666 17196
rect 5000 17184 5028 17224
rect 5534 17212 5540 17224
rect 5592 17212 5598 17264
rect 7374 17212 7380 17264
rect 7432 17252 7438 17264
rect 7432 17224 7880 17252
rect 7432 17212 7438 17224
rect 3660 17156 5028 17184
rect 5077 17187 5135 17193
rect 3660 17144 3666 17156
rect 5077 17153 5089 17187
rect 5123 17184 5135 17187
rect 6273 17187 6331 17193
rect 5123 17156 6224 17184
rect 5123 17153 5135 17156
rect 5077 17147 5135 17153
rect 1857 17119 1915 17125
rect 1857 17085 1869 17119
rect 1903 17116 1915 17119
rect 2777 17119 2835 17125
rect 1903 17088 2360 17116
rect 1903 17085 1915 17088
rect 1857 17079 1915 17085
rect 2130 17048 2136 17060
rect 2091 17020 2136 17048
rect 2130 17008 2136 17020
rect 2188 17008 2194 17060
rect 2332 16980 2360 17088
rect 2777 17085 2789 17119
rect 2823 17116 2835 17119
rect 5350 17116 5356 17128
rect 2823 17088 5356 17116
rect 2823 17085 2835 17088
rect 2777 17079 2835 17085
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 6196 17116 6224 17156
rect 6273 17153 6285 17187
rect 6319 17184 6331 17187
rect 7650 17184 7656 17196
rect 6319 17156 7656 17184
rect 6319 17153 6331 17156
rect 6273 17147 6331 17153
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 7852 17193 7880 17224
rect 8110 17212 8116 17264
rect 8168 17252 8174 17264
rect 12066 17252 12072 17264
rect 8168 17224 8984 17252
rect 8168 17212 8174 17224
rect 8956 17193 8984 17224
rect 10428 17224 12072 17252
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 8941 17187 8999 17193
rect 8941 17153 8953 17187
rect 8987 17153 8999 17187
rect 10226 17184 10232 17196
rect 10187 17156 10232 17184
rect 8941 17147 8999 17153
rect 10226 17144 10232 17156
rect 10284 17144 10290 17196
rect 10428 17193 10456 17224
rect 12066 17212 12072 17224
rect 12124 17212 12130 17264
rect 10413 17187 10471 17193
rect 10413 17153 10425 17187
rect 10459 17153 10471 17187
rect 11974 17184 11980 17196
rect 10413 17147 10471 17153
rect 10980 17156 11980 17184
rect 6730 17116 6736 17128
rect 6196 17088 6736 17116
rect 6730 17076 6736 17088
rect 6788 17076 6794 17128
rect 7006 17076 7012 17128
rect 7064 17116 7070 17128
rect 8849 17119 8907 17125
rect 8849 17116 8861 17119
rect 7064 17088 8861 17116
rect 7064 17076 7070 17088
rect 8849 17085 8861 17088
rect 8895 17085 8907 17119
rect 8849 17079 8907 17085
rect 9122 17076 9128 17128
rect 9180 17116 9186 17128
rect 10502 17116 10508 17128
rect 9180 17088 10508 17116
rect 9180 17076 9186 17088
rect 10502 17076 10508 17088
rect 10560 17076 10566 17128
rect 10980 17125 11008 17156
rect 11974 17144 11980 17156
rect 12032 17144 12038 17196
rect 12986 17144 12992 17196
rect 13044 17184 13050 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 13044 17156 13553 17184
rect 13044 17144 13050 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 13722 17144 13728 17196
rect 13780 17184 13786 17196
rect 13817 17187 13875 17193
rect 13817 17184 13829 17187
rect 13780 17156 13829 17184
rect 13780 17144 13786 17156
rect 13817 17153 13829 17156
rect 13863 17153 13875 17187
rect 13817 17147 13875 17153
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 11701 17119 11759 17125
rect 11701 17085 11713 17119
rect 11747 17085 11759 17119
rect 11701 17079 11759 17085
rect 12621 17119 12679 17125
rect 12621 17085 12633 17119
rect 12667 17116 12679 17119
rect 13170 17116 13176 17128
rect 12667 17088 13176 17116
rect 12667 17085 12679 17088
rect 12621 17079 12679 17085
rect 3050 17048 3056 17060
rect 3011 17020 3056 17048
rect 3050 17008 3056 17020
rect 3108 17008 3114 17060
rect 4338 17008 4344 17060
rect 4396 17048 4402 17060
rect 4893 17051 4951 17057
rect 4893 17048 4905 17051
rect 4396 17020 4905 17048
rect 4396 17008 4402 17020
rect 4893 17017 4905 17020
rect 4939 17017 4951 17051
rect 4893 17011 4951 17017
rect 5997 17051 6055 17057
rect 5997 17017 6009 17051
rect 6043 17048 6055 17051
rect 6362 17048 6368 17060
rect 6043 17020 6368 17048
rect 6043 17017 6055 17020
rect 5997 17011 6055 17017
rect 6362 17008 6368 17020
rect 6420 17008 6426 17060
rect 7558 17048 7564 17060
rect 7519 17020 7564 17048
rect 7558 17008 7564 17020
rect 7616 17008 7622 17060
rect 7653 17051 7711 17057
rect 7653 17017 7665 17051
rect 7699 17048 7711 17051
rect 8757 17051 8815 17057
rect 7699 17020 8715 17048
rect 7699 17017 7711 17020
rect 7653 17011 7711 17017
rect 4433 16983 4491 16989
rect 4433 16980 4445 16983
rect 2332 16952 4445 16980
rect 4433 16949 4445 16952
rect 4479 16949 4491 16983
rect 4433 16943 4491 16949
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 4801 16983 4859 16989
rect 4801 16980 4813 16983
rect 4764 16952 4813 16980
rect 4764 16940 4770 16952
rect 4801 16949 4813 16952
rect 4847 16949 4859 16983
rect 5626 16980 5632 16992
rect 5587 16952 5632 16980
rect 4801 16943 4859 16949
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 6089 16983 6147 16989
rect 6089 16949 6101 16983
rect 6135 16980 6147 16983
rect 6546 16980 6552 16992
rect 6135 16952 6552 16980
rect 6135 16949 6147 16952
rect 6089 16943 6147 16949
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 7193 16983 7251 16989
rect 7193 16949 7205 16983
rect 7239 16980 7251 16983
rect 7926 16980 7932 16992
rect 7239 16952 7932 16980
rect 7239 16949 7251 16952
rect 7193 16943 7251 16949
rect 7926 16940 7932 16952
rect 7984 16940 7990 16992
rect 8386 16980 8392 16992
rect 8347 16952 8392 16980
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 8687 16980 8715 17020
rect 8757 17017 8769 17051
rect 8803 17048 8815 17051
rect 9858 17048 9864 17060
rect 8803 17020 9864 17048
rect 8803 17017 8815 17020
rect 8757 17011 8815 17017
rect 9858 17008 9864 17020
rect 9916 17008 9922 17060
rect 10042 17008 10048 17060
rect 10100 17048 10106 17060
rect 11716 17048 11744 17079
rect 13170 17076 13176 17088
rect 13228 17076 13234 17128
rect 13630 17048 13636 17060
rect 10100 17020 11744 17048
rect 13591 17020 13636 17048
rect 10100 17008 10106 17020
rect 13630 17008 13636 17020
rect 13688 17008 13694 17060
rect 9582 16980 9588 16992
rect 8687 16952 9588 16980
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 9766 16980 9772 16992
rect 9727 16952 9772 16980
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 10137 16983 10195 16989
rect 10137 16949 10149 16983
rect 10183 16980 10195 16983
rect 10410 16980 10416 16992
rect 10183 16952 10416 16980
rect 10183 16949 10195 16952
rect 10137 16943 10195 16949
rect 10410 16940 10416 16952
rect 10468 16940 10474 16992
rect 10594 16940 10600 16992
rect 10652 16980 10658 16992
rect 11149 16983 11207 16989
rect 11149 16980 11161 16983
rect 10652 16952 11161 16980
rect 10652 16940 10658 16952
rect 11149 16949 11161 16952
rect 11195 16949 11207 16983
rect 11149 16943 11207 16949
rect 1104 16890 15824 16912
rect 1104 16838 5912 16890
rect 5964 16838 5976 16890
rect 6028 16838 6040 16890
rect 6092 16838 6104 16890
rect 6156 16838 10843 16890
rect 10895 16838 10907 16890
rect 10959 16838 10971 16890
rect 11023 16838 11035 16890
rect 11087 16838 15824 16890
rect 1104 16816 15824 16838
rect 4614 16736 4620 16788
rect 4672 16776 4678 16788
rect 5258 16776 5264 16788
rect 4672 16748 5264 16776
rect 4672 16736 4678 16748
rect 5258 16736 5264 16748
rect 5316 16736 5322 16788
rect 6270 16736 6276 16788
rect 6328 16776 6334 16788
rect 6917 16779 6975 16785
rect 6917 16776 6929 16779
rect 6328 16748 6929 16776
rect 6328 16736 6334 16748
rect 6917 16745 6929 16748
rect 6963 16745 6975 16779
rect 7282 16776 7288 16788
rect 7243 16748 7288 16776
rect 6917 16739 6975 16745
rect 7282 16736 7288 16748
rect 7340 16736 7346 16788
rect 7558 16736 7564 16788
rect 7616 16776 7622 16788
rect 8386 16776 8392 16788
rect 7616 16748 8392 16776
rect 7616 16736 7622 16748
rect 8386 16736 8392 16748
rect 8444 16736 8450 16788
rect 8573 16779 8631 16785
rect 8573 16745 8585 16779
rect 8619 16776 8631 16779
rect 8662 16776 8668 16788
rect 8619 16748 8668 16776
rect 8619 16745 8631 16748
rect 8573 16739 8631 16745
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 8938 16736 8944 16788
rect 8996 16776 9002 16788
rect 11057 16779 11115 16785
rect 11057 16776 11069 16779
rect 8996 16748 11069 16776
rect 8996 16736 9002 16748
rect 11057 16745 11069 16748
rect 11103 16745 11115 16779
rect 11057 16739 11115 16745
rect 11793 16779 11851 16785
rect 11793 16745 11805 16779
rect 11839 16745 11851 16779
rect 12526 16776 12532 16788
rect 12487 16748 12532 16776
rect 11793 16739 11851 16745
rect 10502 16668 10508 16720
rect 10560 16708 10566 16720
rect 11808 16708 11836 16739
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 13265 16779 13323 16785
rect 13265 16776 13277 16779
rect 12860 16748 13277 16776
rect 12860 16736 12866 16748
rect 13265 16745 13277 16748
rect 13311 16745 13323 16779
rect 13265 16739 13323 16745
rect 10560 16680 11836 16708
rect 10560 16668 10566 16680
rect 1578 16640 1584 16652
rect 1539 16612 1584 16640
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 2498 16640 2504 16652
rect 2459 16612 2504 16640
rect 2498 16600 2504 16612
rect 2556 16600 2562 16652
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 3326 16640 3332 16652
rect 2823 16612 3332 16640
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 3326 16600 3332 16612
rect 3384 16600 3390 16652
rect 3602 16640 3608 16652
rect 3563 16612 3608 16640
rect 3602 16600 3608 16612
rect 3660 16600 3666 16652
rect 4341 16643 4399 16649
rect 4341 16609 4353 16643
rect 4387 16640 4399 16643
rect 4430 16640 4436 16652
rect 4387 16612 4436 16640
rect 4387 16609 4399 16612
rect 4341 16603 4399 16609
rect 4430 16600 4436 16612
rect 4488 16600 4494 16652
rect 4608 16643 4666 16649
rect 4608 16609 4620 16643
rect 4654 16640 4666 16643
rect 6181 16643 6239 16649
rect 4654 16612 6132 16640
rect 4654 16609 4666 16612
rect 4608 16603 4666 16609
rect 6104 16572 6132 16612
rect 6181 16609 6193 16643
rect 6227 16640 6239 16643
rect 7190 16640 7196 16652
rect 6227 16612 7196 16640
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 7377 16643 7435 16649
rect 7377 16609 7389 16643
rect 7423 16640 7435 16643
rect 8481 16643 8539 16649
rect 7423 16612 8432 16640
rect 7423 16609 7435 16612
rect 7377 16603 7435 16609
rect 6638 16572 6644 16584
rect 6104 16544 6644 16572
rect 6638 16532 6644 16544
rect 6696 16572 6702 16584
rect 7561 16575 7619 16581
rect 7561 16572 7573 16575
rect 6696 16544 7573 16572
rect 6696 16532 6702 16544
rect 7561 16541 7573 16544
rect 7607 16572 7619 16575
rect 8202 16572 8208 16584
rect 7607 16544 8208 16572
rect 7607 16541 7619 16544
rect 7561 16535 7619 16541
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 8404 16572 8432 16612
rect 8481 16609 8493 16643
rect 8527 16640 8539 16643
rect 9030 16640 9036 16652
rect 8527 16612 9036 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 9214 16600 9220 16652
rect 9272 16640 9278 16652
rect 10042 16640 10048 16652
rect 9272 16612 10048 16640
rect 9272 16600 9278 16612
rect 10042 16600 10048 16612
rect 10100 16600 10106 16652
rect 10410 16600 10416 16652
rect 10468 16640 10474 16652
rect 10873 16643 10931 16649
rect 10873 16640 10885 16643
rect 10468 16612 10885 16640
rect 10468 16600 10474 16612
rect 10873 16609 10885 16612
rect 10919 16640 10931 16643
rect 11238 16640 11244 16652
rect 10919 16612 11244 16640
rect 10919 16609 10931 16612
rect 10873 16603 10931 16609
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 11606 16640 11612 16652
rect 11567 16612 11612 16640
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 12345 16643 12403 16649
rect 12345 16640 12357 16643
rect 11756 16612 12357 16640
rect 11756 16600 11762 16612
rect 12345 16609 12357 16612
rect 12391 16609 12403 16643
rect 13078 16640 13084 16652
rect 13039 16612 13084 16640
rect 12345 16603 12403 16609
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 13817 16643 13875 16649
rect 13817 16609 13829 16643
rect 13863 16609 13875 16643
rect 13817 16603 13875 16609
rect 8570 16572 8576 16584
rect 8404 16544 8576 16572
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 8757 16575 8815 16581
rect 8757 16572 8769 16575
rect 8667 16544 8769 16572
rect 3142 16464 3148 16516
rect 3200 16504 3206 16516
rect 3421 16507 3479 16513
rect 3421 16504 3433 16507
rect 3200 16476 3433 16504
rect 3200 16464 3206 16476
rect 3421 16473 3433 16476
rect 3467 16473 3479 16507
rect 6365 16507 6423 16513
rect 6365 16504 6377 16507
rect 3421 16467 3479 16473
rect 5644 16476 6377 16504
rect 198 16396 204 16448
rect 256 16436 262 16448
rect 4062 16436 4068 16448
rect 256 16408 4068 16436
rect 256 16396 262 16408
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 4246 16396 4252 16448
rect 4304 16436 4310 16448
rect 4706 16436 4712 16448
rect 4304 16408 4712 16436
rect 4304 16396 4310 16408
rect 4706 16396 4712 16408
rect 4764 16396 4770 16448
rect 4982 16396 4988 16448
rect 5040 16436 5046 16448
rect 5644 16436 5672 16476
rect 6365 16473 6377 16476
rect 6411 16473 6423 16507
rect 8687 16504 8715 16544
rect 8757 16541 8769 16544
rect 8803 16572 8815 16575
rect 9306 16572 9312 16584
rect 8803 16544 9312 16572
rect 8803 16541 8815 16544
rect 8757 16535 8815 16541
rect 9306 16532 9312 16544
rect 9364 16532 9370 16584
rect 10134 16572 10140 16584
rect 10095 16544 10140 16572
rect 10134 16532 10140 16544
rect 10192 16532 10198 16584
rect 10321 16575 10379 16581
rect 10321 16541 10333 16575
rect 10367 16572 10379 16575
rect 10962 16572 10968 16584
rect 10367 16544 10968 16572
rect 10367 16541 10379 16544
rect 10321 16535 10379 16541
rect 10336 16504 10364 16535
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 13832 16572 13860 16603
rect 11624 16544 13860 16572
rect 11624 16516 11652 16544
rect 13998 16532 14004 16584
rect 14056 16572 14062 16584
rect 14553 16575 14611 16581
rect 14553 16572 14565 16575
rect 14056 16544 14565 16572
rect 14056 16532 14062 16544
rect 14553 16541 14565 16544
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 6365 16467 6423 16473
rect 6472 16476 8715 16504
rect 8772 16476 10364 16504
rect 5040 16408 5672 16436
rect 5721 16439 5779 16445
rect 5040 16396 5046 16408
rect 5721 16405 5733 16439
rect 5767 16436 5779 16439
rect 5810 16436 5816 16448
rect 5767 16408 5816 16436
rect 5767 16405 5779 16408
rect 5721 16399 5779 16405
rect 5810 16396 5816 16408
rect 5868 16396 5874 16448
rect 5902 16396 5908 16448
rect 5960 16436 5966 16448
rect 6472 16436 6500 16476
rect 5960 16408 6500 16436
rect 5960 16396 5966 16408
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 8113 16439 8171 16445
rect 8113 16436 8125 16439
rect 6972 16408 8125 16436
rect 6972 16396 6978 16408
rect 8113 16405 8125 16408
rect 8159 16405 8171 16439
rect 8113 16399 8171 16405
rect 8202 16396 8208 16448
rect 8260 16436 8266 16448
rect 8772 16436 8800 16476
rect 11606 16464 11612 16516
rect 11664 16464 11670 16516
rect 8260 16408 8800 16436
rect 8260 16396 8266 16408
rect 8846 16396 8852 16448
rect 8904 16436 8910 16448
rect 9677 16439 9735 16445
rect 9677 16436 9689 16439
rect 8904 16408 9689 16436
rect 8904 16396 8910 16408
rect 9677 16405 9689 16408
rect 9723 16405 9735 16439
rect 9677 16399 9735 16405
rect 11146 16396 11152 16448
rect 11204 16436 11210 16448
rect 11882 16436 11888 16448
rect 11204 16408 11888 16436
rect 11204 16396 11210 16408
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 12158 16396 12164 16448
rect 12216 16436 12222 16448
rect 14001 16439 14059 16445
rect 14001 16436 14013 16439
rect 12216 16408 14013 16436
rect 12216 16396 12222 16408
rect 14001 16405 14013 16408
rect 14047 16405 14059 16439
rect 14001 16399 14059 16405
rect 14274 16396 14280 16448
rect 14332 16436 14338 16448
rect 14550 16436 14556 16448
rect 14332 16408 14556 16436
rect 14332 16396 14338 16408
rect 14550 16396 14556 16408
rect 14608 16396 14614 16448
rect 1104 16346 15824 16368
rect 1104 16294 3447 16346
rect 3499 16294 3511 16346
rect 3563 16294 3575 16346
rect 3627 16294 3639 16346
rect 3691 16294 8378 16346
rect 8430 16294 8442 16346
rect 8494 16294 8506 16346
rect 8558 16294 8570 16346
rect 8622 16294 13308 16346
rect 13360 16294 13372 16346
rect 13424 16294 13436 16346
rect 13488 16294 13500 16346
rect 13552 16294 15824 16346
rect 1104 16272 15824 16294
rect 1581 16235 1639 16241
rect 1581 16201 1593 16235
rect 1627 16232 1639 16235
rect 2866 16232 2872 16244
rect 1627 16204 2872 16232
rect 1627 16201 1639 16204
rect 1581 16195 1639 16201
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 3145 16235 3203 16241
rect 3145 16201 3157 16235
rect 3191 16232 3203 16235
rect 5718 16232 5724 16244
rect 3191 16204 5724 16232
rect 3191 16201 3203 16204
rect 3145 16195 3203 16201
rect 5718 16192 5724 16204
rect 5776 16192 5782 16244
rect 6917 16235 6975 16241
rect 6917 16201 6929 16235
rect 6963 16232 6975 16235
rect 7006 16232 7012 16244
rect 6963 16204 7012 16232
rect 6963 16201 6975 16204
rect 6917 16195 6975 16201
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 7098 16192 7104 16244
rect 7156 16232 7162 16244
rect 8846 16232 8852 16244
rect 7156 16204 8852 16232
rect 7156 16192 7162 16204
rect 8846 16192 8852 16204
rect 8904 16192 8910 16244
rect 9766 16232 9772 16244
rect 8956 16204 9772 16232
rect 3970 16164 3976 16176
rect 3620 16136 3976 16164
rect 2501 16099 2559 16105
rect 2501 16065 2513 16099
rect 2547 16096 2559 16099
rect 2774 16096 2780 16108
rect 2547 16068 2780 16096
rect 2547 16065 2559 16068
rect 2501 16059 2559 16065
rect 2774 16056 2780 16068
rect 2832 16056 2838 16108
rect 3620 16105 3648 16136
rect 3970 16124 3976 16136
rect 4028 16124 4034 16176
rect 4341 16167 4399 16173
rect 4341 16133 4353 16167
rect 4387 16164 4399 16167
rect 5166 16164 5172 16176
rect 4387 16136 5172 16164
rect 4387 16133 4399 16136
rect 4341 16127 4399 16133
rect 5166 16124 5172 16136
rect 5224 16124 5230 16176
rect 5258 16124 5264 16176
rect 5316 16164 5322 16176
rect 8297 16167 8355 16173
rect 8297 16164 8309 16167
rect 5316 16136 8309 16164
rect 5316 16124 5322 16136
rect 8297 16133 8309 16136
rect 8343 16133 8355 16167
rect 8297 16127 8355 16133
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16065 3663 16099
rect 3605 16059 3663 16065
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16096 3847 16099
rect 4614 16096 4620 16108
rect 3835 16068 4620 16096
rect 3835 16065 3847 16068
rect 3789 16059 3847 16065
rect 4614 16056 4620 16068
rect 4672 16056 4678 16108
rect 4798 16096 4804 16108
rect 4759 16068 4804 16096
rect 4798 16056 4804 16068
rect 4856 16056 4862 16108
rect 4982 16096 4988 16108
rect 4895 16068 4988 16096
rect 4982 16056 4988 16068
rect 5040 16096 5046 16108
rect 5902 16096 5908 16108
rect 5040 16068 5908 16096
rect 5040 16056 5046 16068
rect 5902 16056 5908 16068
rect 5960 16056 5966 16108
rect 6181 16099 6239 16105
rect 6181 16065 6193 16099
rect 6227 16096 6239 16099
rect 7190 16096 7196 16108
rect 6227 16068 7196 16096
rect 6227 16065 6239 16068
rect 6181 16059 6239 16065
rect 7190 16056 7196 16068
rect 7248 16056 7254 16108
rect 7466 16056 7472 16108
rect 7524 16056 7530 16108
rect 7561 16099 7619 16105
rect 7561 16065 7573 16099
rect 7607 16096 7619 16099
rect 7607 16068 7696 16096
rect 7607 16065 7619 16068
rect 7561 16059 7619 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 1397 15991 1455 15997
rect 2225 16031 2283 16037
rect 2225 15997 2237 16031
rect 2271 16028 2283 16031
rect 5074 16028 5080 16040
rect 2271 16000 5080 16028
rect 2271 15997 2283 16000
rect 2225 15991 2283 15997
rect 1412 15960 1440 15991
rect 5074 15988 5080 16000
rect 5132 15988 5138 16040
rect 5997 16031 6055 16037
rect 5997 15997 6009 16031
rect 6043 16028 6055 16031
rect 7484 16028 7512 16056
rect 6043 16000 7512 16028
rect 6043 15997 6055 16000
rect 5997 15991 6055 15997
rect 1412 15932 2084 15960
rect 2056 15892 2084 15932
rect 2314 15920 2320 15972
rect 2372 15960 2378 15972
rect 5905 15963 5963 15969
rect 2372 15932 5663 15960
rect 2372 15920 2378 15932
rect 2774 15892 2780 15904
rect 2056 15864 2780 15892
rect 2774 15852 2780 15864
rect 2832 15852 2838 15904
rect 3234 15852 3240 15904
rect 3292 15892 3298 15904
rect 3513 15895 3571 15901
rect 3513 15892 3525 15895
rect 3292 15864 3525 15892
rect 3292 15852 3298 15864
rect 3513 15861 3525 15864
rect 3559 15861 3571 15895
rect 3513 15855 3571 15861
rect 4709 15895 4767 15901
rect 4709 15861 4721 15895
rect 4755 15892 4767 15895
rect 4890 15892 4896 15904
rect 4755 15864 4896 15892
rect 4755 15861 4767 15864
rect 4709 15855 4767 15861
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 5074 15852 5080 15904
rect 5132 15892 5138 15904
rect 5537 15895 5595 15901
rect 5537 15892 5549 15895
rect 5132 15864 5549 15892
rect 5132 15852 5138 15864
rect 5537 15861 5549 15864
rect 5583 15861 5595 15895
rect 5635 15892 5663 15932
rect 5905 15929 5917 15963
rect 5951 15960 5963 15963
rect 7466 15960 7472 15972
rect 5951 15932 7472 15960
rect 5951 15929 5963 15932
rect 5905 15923 5963 15929
rect 7466 15920 7472 15932
rect 7524 15920 7530 15972
rect 7558 15920 7564 15972
rect 7616 15960 7622 15972
rect 7668 15960 7696 16068
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 8956 16096 8984 16204
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 10962 16192 10968 16244
rect 11020 16232 11026 16244
rect 11330 16232 11336 16244
rect 11020 16204 11336 16232
rect 11020 16192 11026 16204
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 9674 16124 9680 16176
rect 9732 16164 9738 16176
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 9732 16136 11805 16164
rect 9732 16124 9738 16136
rect 11793 16133 11805 16136
rect 11839 16133 11851 16167
rect 11793 16127 11851 16133
rect 11882 16124 11888 16176
rect 11940 16164 11946 16176
rect 13817 16167 13875 16173
rect 13817 16164 13829 16167
rect 11940 16136 13829 16164
rect 11940 16124 11946 16136
rect 13817 16133 13829 16136
rect 13863 16133 13875 16167
rect 13817 16127 13875 16133
rect 7800 16068 8984 16096
rect 7800 16056 7806 16068
rect 9122 16056 9128 16108
rect 9180 16056 9186 16108
rect 9490 16056 9496 16108
rect 9548 16096 9554 16108
rect 9769 16099 9827 16105
rect 9769 16096 9781 16099
rect 9548 16068 9781 16096
rect 9548 16056 9554 16068
rect 9769 16065 9781 16068
rect 9815 16065 9827 16099
rect 10962 16096 10968 16108
rect 9769 16059 9827 16065
rect 9968 16068 10180 16096
rect 10923 16068 10968 16096
rect 8018 15988 8024 16040
rect 8076 16028 8082 16040
rect 8113 16031 8171 16037
rect 8113 16028 8125 16031
rect 8076 16000 8125 16028
rect 8076 15988 8082 16000
rect 8113 15997 8125 16000
rect 8159 15997 8171 16031
rect 8113 15991 8171 15997
rect 8294 15988 8300 16040
rect 8352 16028 8358 16040
rect 9140 16028 9168 16056
rect 8352 16000 9168 16028
rect 8352 15988 8358 16000
rect 9214 15988 9220 16040
rect 9272 15988 9278 16040
rect 9585 16031 9643 16037
rect 9585 15997 9597 16031
rect 9631 16028 9643 16031
rect 9968 16028 9996 16068
rect 9631 16000 9996 16028
rect 10152 16028 10180 16068
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 12710 16096 12716 16108
rect 11348 16068 12716 16096
rect 11348 16028 11376 16068
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 12986 16096 12992 16108
rect 12820 16068 12992 16096
rect 10152 16000 11376 16028
rect 9631 15997 9643 16000
rect 9585 15991 9643 15997
rect 11422 15988 11428 16040
rect 11480 16028 11486 16040
rect 11609 16031 11667 16037
rect 11609 16028 11621 16031
rect 11480 16000 11621 16028
rect 11480 15988 11486 16000
rect 11609 15997 11621 16000
rect 11655 15997 11667 16031
rect 11609 15991 11667 15997
rect 11698 15988 11704 16040
rect 11756 16028 11762 16040
rect 12820 16037 12848 16068
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 14921 16099 14979 16105
rect 14921 16065 14933 16099
rect 14967 16096 14979 16099
rect 16758 16096 16764 16108
rect 14967 16068 16764 16096
rect 14967 16065 14979 16068
rect 14921 16059 14979 16065
rect 16758 16056 16764 16068
rect 16816 16056 16822 16108
rect 12437 16031 12495 16037
rect 12437 16028 12449 16031
rect 11756 16000 12449 16028
rect 11756 15988 11762 16000
rect 12437 15997 12449 16000
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 12805 16031 12863 16037
rect 12805 15997 12817 16031
rect 12851 15997 12863 16031
rect 12805 15991 12863 15997
rect 9122 15960 9128 15972
rect 7616 15932 7696 15960
rect 8404 15932 9128 15960
rect 7616 15920 7622 15932
rect 7098 15892 7104 15904
rect 5635 15864 7104 15892
rect 5537 15855 5595 15861
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 7282 15892 7288 15904
rect 7243 15864 7288 15892
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 7377 15895 7435 15901
rect 7377 15861 7389 15895
rect 7423 15892 7435 15895
rect 8404 15892 8432 15932
rect 9122 15920 9128 15932
rect 9180 15920 9186 15972
rect 9232 15960 9260 15988
rect 10873 15963 10931 15969
rect 9232 15932 10456 15960
rect 7423 15864 8432 15892
rect 7423 15861 7435 15864
rect 7377 15855 7435 15861
rect 8478 15852 8484 15904
rect 8536 15892 8542 15904
rect 9217 15895 9275 15901
rect 9217 15892 9229 15895
rect 8536 15864 9229 15892
rect 8536 15852 8542 15864
rect 9217 15861 9229 15864
rect 9263 15861 9275 15895
rect 9217 15855 9275 15861
rect 9582 15852 9588 15904
rect 9640 15892 9646 15904
rect 9677 15895 9735 15901
rect 9677 15892 9689 15895
rect 9640 15864 9689 15892
rect 9640 15852 9646 15864
rect 9677 15861 9689 15864
rect 9723 15861 9735 15895
rect 9677 15855 9735 15861
rect 9766 15852 9772 15904
rect 9824 15892 9830 15904
rect 10134 15892 10140 15904
rect 9824 15864 10140 15892
rect 9824 15852 9830 15864
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 10428 15901 10456 15932
rect 10873 15929 10885 15963
rect 10919 15960 10931 15963
rect 12452 15960 12480 15991
rect 12894 15988 12900 16040
rect 12952 16028 12958 16040
rect 13633 16031 13691 16037
rect 13633 16028 13645 16031
rect 12952 16000 13645 16028
rect 12952 15988 12958 16000
rect 13633 15997 13645 16000
rect 13679 15997 13691 16031
rect 14642 16028 14648 16040
rect 14603 16000 14648 16028
rect 13633 15991 13691 15997
rect 14642 15988 14648 16000
rect 14700 15988 14706 16040
rect 13265 15963 13323 15969
rect 13265 15960 13277 15963
rect 10919 15932 11928 15960
rect 12452 15932 13277 15960
rect 10919 15929 10931 15932
rect 10873 15923 10931 15929
rect 10413 15895 10471 15901
rect 10413 15861 10425 15895
rect 10459 15861 10471 15895
rect 10413 15855 10471 15861
rect 10781 15895 10839 15901
rect 10781 15861 10793 15895
rect 10827 15892 10839 15895
rect 11238 15892 11244 15904
rect 10827 15864 11244 15892
rect 10827 15861 10839 15864
rect 10781 15855 10839 15861
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 11900 15892 11928 15932
rect 13265 15929 13277 15932
rect 13311 15929 13323 15963
rect 13265 15923 13323 15929
rect 12802 15892 12808 15904
rect 11900 15864 12808 15892
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 13630 15892 13636 15904
rect 12943 15864 13636 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 13630 15852 13636 15864
rect 13688 15852 13694 15904
rect 1104 15802 15824 15824
rect 1104 15750 5912 15802
rect 5964 15750 5976 15802
rect 6028 15750 6040 15802
rect 6092 15750 6104 15802
rect 6156 15750 10843 15802
rect 10895 15750 10907 15802
rect 10959 15750 10971 15802
rect 11023 15750 11035 15802
rect 11087 15750 15824 15802
rect 1104 15728 15824 15750
rect 3145 15691 3203 15697
rect 3145 15657 3157 15691
rect 3191 15688 3203 15691
rect 5074 15688 5080 15700
rect 3191 15660 5080 15688
rect 3191 15657 3203 15660
rect 3145 15651 3203 15657
rect 5074 15648 5080 15660
rect 5132 15648 5138 15700
rect 5350 15688 5356 15700
rect 5311 15660 5356 15688
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 6914 15688 6920 15700
rect 6875 15660 6920 15688
rect 6914 15648 6920 15660
rect 6972 15648 6978 15700
rect 8113 15691 8171 15697
rect 8113 15657 8125 15691
rect 8159 15688 8171 15691
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 8159 15660 9689 15688
rect 8159 15657 8171 15660
rect 8113 15651 8171 15657
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 9677 15651 9735 15657
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 10137 15691 10195 15697
rect 10137 15688 10149 15691
rect 9824 15660 10149 15688
rect 9824 15648 9830 15660
rect 10137 15657 10149 15660
rect 10183 15657 10195 15691
rect 10137 15651 10195 15657
rect 10410 15648 10416 15700
rect 10468 15688 10474 15700
rect 10686 15688 10692 15700
rect 10468 15660 10692 15688
rect 10468 15648 10474 15660
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 12250 15648 12256 15700
rect 12308 15688 12314 15700
rect 13446 15688 13452 15700
rect 12308 15660 13308 15688
rect 13407 15660 13452 15688
rect 12308 15648 12314 15660
rect 6086 15620 6092 15632
rect 4356 15592 6092 15620
rect 1210 15512 1216 15564
rect 1268 15552 1274 15564
rect 1857 15555 1915 15561
rect 1857 15552 1869 15555
rect 1268 15524 1869 15552
rect 1268 15512 1274 15524
rect 1857 15521 1869 15524
rect 1903 15521 1915 15555
rect 1857 15515 1915 15521
rect 3237 15555 3295 15561
rect 3237 15521 3249 15555
rect 3283 15552 3295 15555
rect 4154 15552 4160 15564
rect 3283 15524 4160 15552
rect 3283 15521 3295 15524
rect 3237 15515 3295 15521
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15484 2191 15487
rect 2958 15484 2964 15496
rect 2179 15456 2964 15484
rect 2179 15453 2191 15456
rect 2133 15447 2191 15453
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 3421 15487 3479 15493
rect 3421 15484 3433 15487
rect 3068 15456 3433 15484
rect 2866 15376 2872 15428
rect 2924 15416 2930 15428
rect 3068 15416 3096 15456
rect 3421 15453 3433 15456
rect 3467 15484 3479 15487
rect 4356 15484 4384 15592
rect 6086 15580 6092 15592
rect 6144 15580 6150 15632
rect 10962 15620 10968 15632
rect 7024 15592 10968 15620
rect 4522 15552 4528 15564
rect 4483 15524 4528 15552
rect 4522 15512 4528 15524
rect 4580 15512 4586 15564
rect 4614 15512 4620 15564
rect 4672 15552 4678 15564
rect 7024 15561 7052 15592
rect 10962 15580 10968 15592
rect 11020 15580 11026 15632
rect 11333 15623 11391 15629
rect 11333 15589 11345 15623
rect 11379 15620 11391 15623
rect 11422 15620 11428 15632
rect 11379 15592 11428 15620
rect 11379 15589 11391 15592
rect 11333 15583 11391 15589
rect 11422 15580 11428 15592
rect 11480 15580 11486 15632
rect 12066 15580 12072 15632
rect 12124 15620 12130 15632
rect 12124 15592 12664 15620
rect 12124 15580 12130 15592
rect 5721 15555 5779 15561
rect 4672 15524 4717 15552
rect 4672 15512 4678 15524
rect 5721 15521 5733 15555
rect 5767 15552 5779 15555
rect 7009 15555 7067 15561
rect 5767 15524 6960 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 3467 15456 4384 15484
rect 4801 15487 4859 15493
rect 3467 15453 3479 15456
rect 3421 15447 3479 15453
rect 4801 15453 4813 15487
rect 4847 15484 4859 15487
rect 5258 15484 5264 15496
rect 4847 15456 5264 15484
rect 4847 15453 4859 15456
rect 4801 15447 4859 15453
rect 5258 15444 5264 15456
rect 5316 15444 5322 15496
rect 5810 15484 5816 15496
rect 5771 15456 5816 15484
rect 5810 15444 5816 15456
rect 5868 15444 5874 15496
rect 5997 15487 6055 15493
rect 5997 15453 6009 15487
rect 6043 15484 6055 15487
rect 6454 15484 6460 15496
rect 6043 15456 6460 15484
rect 6043 15453 6055 15456
rect 5997 15447 6055 15453
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 6932 15484 6960 15524
rect 7009 15521 7021 15555
rect 7055 15521 7067 15555
rect 7009 15515 7067 15521
rect 7466 15512 7472 15564
rect 7524 15512 7530 15564
rect 8205 15555 8263 15561
rect 8205 15521 8217 15555
rect 8251 15552 8263 15555
rect 8251 15524 8616 15552
rect 8251 15521 8263 15524
rect 8205 15515 8263 15521
rect 7098 15484 7104 15496
rect 6932 15456 7104 15484
rect 7098 15444 7104 15456
rect 7156 15444 7162 15496
rect 7193 15487 7251 15493
rect 7193 15453 7205 15487
rect 7239 15453 7251 15487
rect 7484 15484 7512 15512
rect 7484 15456 7788 15484
rect 7193 15447 7251 15453
rect 2924 15388 3096 15416
rect 2924 15376 2930 15388
rect 3234 15376 3240 15428
rect 3292 15416 3298 15428
rect 7006 15416 7012 15428
rect 3292 15388 7012 15416
rect 3292 15376 3298 15388
rect 7006 15376 7012 15388
rect 7064 15376 7070 15428
rect 7208 15416 7236 15447
rect 7466 15416 7472 15428
rect 7208 15388 7472 15416
rect 7466 15376 7472 15388
rect 7524 15376 7530 15428
rect 7760 15425 7788 15456
rect 7834 15444 7840 15496
rect 7892 15484 7898 15496
rect 8110 15484 8116 15496
rect 7892 15456 8116 15484
rect 7892 15444 7898 15456
rect 8110 15444 8116 15456
rect 8168 15484 8174 15496
rect 8297 15487 8355 15493
rect 8297 15484 8309 15487
rect 8168 15456 8309 15484
rect 8168 15444 8174 15456
rect 8297 15453 8309 15456
rect 8343 15453 8355 15487
rect 8297 15447 8355 15453
rect 7745 15419 7803 15425
rect 7745 15385 7757 15419
rect 7791 15385 7803 15419
rect 8588 15416 8616 15524
rect 8662 15512 8668 15564
rect 8720 15512 8726 15564
rect 8846 15512 8852 15564
rect 8904 15552 8910 15564
rect 9306 15552 9312 15564
rect 8904 15524 9312 15552
rect 8904 15512 8910 15524
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 10045 15555 10103 15561
rect 10045 15521 10057 15555
rect 10091 15552 10103 15555
rect 10091 15524 10456 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 8680 15484 8708 15512
rect 10428 15496 10456 15524
rect 11054 15512 11060 15564
rect 11112 15552 11118 15564
rect 11241 15555 11299 15561
rect 11241 15552 11253 15555
rect 11112 15524 11253 15552
rect 11112 15512 11118 15524
rect 11241 15521 11253 15524
rect 11287 15521 11299 15555
rect 11241 15515 11299 15521
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8680 15456 8953 15484
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 8941 15447 8999 15453
rect 9048 15456 10241 15484
rect 8846 15416 8852 15428
rect 8588 15388 8852 15416
rect 7745 15379 7803 15385
rect 8846 15376 8852 15388
rect 8904 15376 8910 15428
rect 2777 15351 2835 15357
rect 2777 15317 2789 15351
rect 2823 15348 2835 15351
rect 3970 15348 3976 15360
rect 2823 15320 3976 15348
rect 2823 15317 2835 15320
rect 2777 15311 2835 15317
rect 3970 15308 3976 15320
rect 4028 15308 4034 15360
rect 4154 15348 4160 15360
rect 4115 15320 4160 15348
rect 4154 15308 4160 15320
rect 4212 15308 4218 15360
rect 6546 15348 6552 15360
rect 6507 15320 6552 15348
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 7558 15308 7564 15360
rect 7616 15348 7622 15360
rect 8110 15348 8116 15360
rect 7616 15320 8116 15348
rect 7616 15308 7622 15320
rect 8110 15308 8116 15320
rect 8168 15348 8174 15360
rect 9048 15348 9076 15456
rect 10060 15428 10088 15456
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 10410 15444 10416 15496
rect 10468 15444 10474 15496
rect 10870 15444 10876 15496
rect 10928 15484 10934 15496
rect 11425 15487 11483 15493
rect 11425 15484 11437 15487
rect 10928 15456 11437 15484
rect 10928 15444 10934 15456
rect 11425 15453 11437 15456
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 11882 15444 11888 15496
rect 11940 15484 11946 15496
rect 12084 15484 12112 15580
rect 12434 15512 12440 15564
rect 12492 15552 12498 15564
rect 12492 15524 12537 15552
rect 12492 15512 12498 15524
rect 12526 15484 12532 15496
rect 11940 15456 12112 15484
rect 12487 15456 12532 15484
rect 11940 15444 11946 15456
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 12636 15493 12664 15592
rect 12802 15512 12808 15564
rect 12860 15512 12866 15564
rect 13280 15561 13308 15660
rect 13446 15648 13452 15660
rect 13504 15648 13510 15700
rect 14182 15688 14188 15700
rect 14143 15660 14188 15688
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 13265 15555 13323 15561
rect 13265 15521 13277 15555
rect 13311 15521 13323 15555
rect 13265 15515 13323 15521
rect 14001 15555 14059 15561
rect 14001 15521 14013 15555
rect 14047 15552 14059 15555
rect 14090 15552 14096 15564
rect 14047 15524 14096 15552
rect 14047 15521 14059 15524
rect 14001 15515 14059 15521
rect 14090 15512 14096 15524
rect 14148 15512 14154 15564
rect 12621 15487 12679 15493
rect 12621 15453 12633 15487
rect 12667 15453 12679 15487
rect 12820 15484 12848 15512
rect 15286 15484 15292 15496
rect 12820 15456 15292 15484
rect 12621 15447 12679 15453
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 9214 15376 9220 15428
rect 9272 15416 9278 15428
rect 9674 15416 9680 15428
rect 9272 15388 9680 15416
rect 9272 15376 9278 15388
rect 9674 15376 9680 15388
rect 9732 15376 9738 15428
rect 10042 15376 10048 15428
rect 10100 15376 10106 15428
rect 10962 15376 10968 15428
rect 11020 15416 11026 15428
rect 12342 15416 12348 15428
rect 11020 15388 12348 15416
rect 11020 15376 11026 15388
rect 12342 15376 12348 15388
rect 12400 15376 12406 15428
rect 8168 15320 9076 15348
rect 8168 15308 8174 15320
rect 9122 15308 9128 15360
rect 9180 15348 9186 15360
rect 10873 15351 10931 15357
rect 10873 15348 10885 15351
rect 9180 15320 10885 15348
rect 9180 15308 9186 15320
rect 10873 15317 10885 15320
rect 10919 15317 10931 15351
rect 12066 15348 12072 15360
rect 12027 15320 12072 15348
rect 10873 15311 10931 15317
rect 12066 15308 12072 15320
rect 12124 15308 12130 15360
rect 1104 15258 15824 15280
rect 1104 15206 3447 15258
rect 3499 15206 3511 15258
rect 3563 15206 3575 15258
rect 3627 15206 3639 15258
rect 3691 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 13308 15258
rect 13360 15206 13372 15258
rect 13424 15206 13436 15258
rect 13488 15206 13500 15258
rect 13552 15206 15824 15258
rect 1104 15184 15824 15206
rect 2498 15104 2504 15156
rect 2556 15144 2562 15156
rect 4338 15144 4344 15156
rect 2556 15116 4344 15144
rect 2556 15104 2562 15116
rect 4338 15104 4344 15116
rect 4396 15104 4402 15156
rect 5350 15144 5356 15156
rect 4448 15116 5356 15144
rect 3145 15079 3203 15085
rect 3145 15045 3157 15079
rect 3191 15076 3203 15079
rect 3878 15076 3884 15088
rect 3191 15048 3884 15076
rect 3191 15045 3203 15048
rect 3145 15039 3203 15045
rect 3878 15036 3884 15048
rect 3936 15036 3942 15088
rect 2593 15011 2651 15017
rect 2593 14977 2605 15011
rect 2639 15008 2651 15011
rect 2866 15008 2872 15020
rect 2639 14980 2872 15008
rect 2639 14977 2651 14980
rect 2593 14971 2651 14977
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 3786 15008 3792 15020
rect 3747 14980 3792 15008
rect 3786 14968 3792 14980
rect 3844 14968 3850 15020
rect 4448 15008 4476 15116
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 5810 15104 5816 15156
rect 5868 15144 5874 15156
rect 6825 15147 6883 15153
rect 6825 15144 6837 15147
rect 5868 15116 6837 15144
rect 5868 15104 5874 15116
rect 6825 15113 6837 15116
rect 6871 15113 6883 15147
rect 6825 15107 6883 15113
rect 7374 15104 7380 15156
rect 7432 15144 7438 15156
rect 9582 15144 9588 15156
rect 7432 15116 9588 15144
rect 7432 15104 7438 15116
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 10686 15104 10692 15156
rect 10744 15144 10750 15156
rect 13357 15147 13415 15153
rect 13357 15144 13369 15147
rect 10744 15116 13369 15144
rect 10744 15104 10750 15116
rect 13357 15113 13369 15116
rect 13403 15113 13415 15147
rect 13357 15107 13415 15113
rect 4706 15036 4712 15088
rect 4764 15076 4770 15088
rect 8938 15076 8944 15088
rect 4764 15048 8944 15076
rect 4764 15036 4770 15048
rect 8938 15036 8944 15048
rect 8996 15036 9002 15088
rect 9858 15076 9864 15088
rect 9048 15048 9343 15076
rect 9819 15048 9864 15076
rect 4982 15008 4988 15020
rect 3988 14980 4476 15008
rect 4943 14980 4988 15008
rect 1670 14832 1676 14884
rect 1728 14872 1734 14884
rect 2409 14875 2467 14881
rect 2409 14872 2421 14875
rect 1728 14844 2421 14872
rect 1728 14832 1734 14844
rect 2409 14841 2421 14844
rect 2455 14872 2467 14875
rect 2682 14872 2688 14884
rect 2455 14844 2688 14872
rect 2455 14841 2467 14844
rect 2409 14835 2467 14841
rect 2682 14832 2688 14844
rect 2740 14832 2746 14884
rect 2774 14832 2780 14884
rect 2832 14872 2838 14884
rect 3605 14875 3663 14881
rect 3605 14872 3617 14875
rect 2832 14844 3617 14872
rect 2832 14832 2838 14844
rect 3605 14841 3617 14844
rect 3651 14841 3663 14875
rect 3605 14835 3663 14841
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 1949 14807 2007 14813
rect 1949 14804 1961 14807
rect 1820 14776 1961 14804
rect 1820 14764 1826 14776
rect 1949 14773 1961 14776
rect 1995 14773 2007 14807
rect 1949 14767 2007 14773
rect 2317 14807 2375 14813
rect 2317 14773 2329 14807
rect 2363 14804 2375 14807
rect 2866 14804 2872 14816
rect 2363 14776 2872 14804
rect 2363 14773 2375 14776
rect 2317 14767 2375 14773
rect 2866 14764 2872 14776
rect 2924 14764 2930 14816
rect 3513 14807 3571 14813
rect 3513 14773 3525 14807
rect 3559 14804 3571 14807
rect 3988 14804 4016 14980
rect 4982 14968 4988 14980
rect 5040 14968 5046 15020
rect 5350 14968 5356 15020
rect 5408 15008 5414 15020
rect 5408 14980 5764 15008
rect 5408 14968 5414 14980
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4614 14940 4620 14952
rect 4120 14912 4620 14940
rect 4120 14900 4126 14912
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 5626 14940 5632 14952
rect 5184 14912 5632 14940
rect 4709 14875 4767 14881
rect 4709 14841 4721 14875
rect 4755 14872 4767 14875
rect 4755 14844 4936 14872
rect 4755 14841 4767 14844
rect 4709 14835 4767 14841
rect 4338 14804 4344 14816
rect 3559 14776 4016 14804
rect 4299 14776 4344 14804
rect 3559 14773 3571 14776
rect 3513 14767 3571 14773
rect 4338 14764 4344 14776
rect 4396 14764 4402 14816
rect 4798 14804 4804 14816
rect 4759 14776 4804 14804
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 4908 14804 4936 14844
rect 5184 14804 5212 14912
rect 5626 14900 5632 14912
rect 5684 14900 5690 14952
rect 5736 14940 5764 14980
rect 5810 14968 5816 15020
rect 5868 15008 5874 15020
rect 5997 15011 6055 15017
rect 5997 15008 6009 15011
rect 5868 14980 6009 15008
rect 5868 14968 5874 14980
rect 5997 14977 6009 14980
rect 6043 14977 6055 15011
rect 5997 14971 6055 14977
rect 6086 14968 6092 15020
rect 6144 15008 6150 15020
rect 7469 15011 7527 15017
rect 6144 14980 6189 15008
rect 6144 14968 6150 14980
rect 7469 14977 7481 15011
rect 7515 15008 7527 15011
rect 7558 15008 7564 15020
rect 7515 14980 7564 15008
rect 7515 14977 7527 14980
rect 7469 14971 7527 14977
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 7926 14968 7932 15020
rect 7984 15008 7990 15020
rect 9048 15008 9076 15048
rect 9214 15008 9220 15020
rect 7984 14980 9076 15008
rect 9175 14980 9220 15008
rect 7984 14968 7990 14980
rect 9214 14968 9220 14980
rect 9272 14968 9278 15020
rect 9315 15008 9343 15048
rect 9858 15036 9864 15048
rect 9916 15036 9922 15088
rect 10042 15036 10048 15088
rect 10100 15076 10106 15088
rect 12621 15079 12679 15085
rect 10100 15048 10456 15076
rect 10100 15036 10106 15048
rect 10428 15017 10456 15048
rect 12621 15045 12633 15079
rect 12667 15076 12679 15079
rect 13078 15076 13084 15088
rect 12667 15048 13084 15076
rect 12667 15045 12679 15048
rect 12621 15039 12679 15045
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 13814 15036 13820 15088
rect 13872 15076 13878 15088
rect 14093 15079 14151 15085
rect 14093 15076 14105 15079
rect 13872 15048 14105 15076
rect 13872 15036 13878 15048
rect 14093 15045 14105 15048
rect 14139 15045 14151 15079
rect 14093 15039 14151 15045
rect 10321 15011 10379 15017
rect 10321 15008 10333 15011
rect 9315 14980 10333 15008
rect 10321 14977 10333 14980
rect 10367 14977 10379 15011
rect 10321 14971 10379 14977
rect 10413 15011 10471 15017
rect 10413 14977 10425 15011
rect 10459 15008 10471 15011
rect 11882 15008 11888 15020
rect 10459 14980 11888 15008
rect 10459 14977 10471 14980
rect 10413 14971 10471 14977
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 5905 14943 5963 14949
rect 5905 14940 5917 14943
rect 5736 14912 5917 14940
rect 5905 14909 5917 14912
rect 5951 14940 5963 14943
rect 6362 14940 6368 14952
rect 5951 14912 6368 14940
rect 5951 14909 5963 14912
rect 5905 14903 5963 14909
rect 6362 14900 6368 14912
rect 6420 14900 6426 14952
rect 7193 14943 7251 14949
rect 7193 14909 7205 14943
rect 7239 14940 7251 14943
rect 7742 14940 7748 14952
rect 7239 14912 7748 14940
rect 7239 14909 7251 14912
rect 7193 14903 7251 14909
rect 7742 14900 7748 14912
rect 7800 14900 7806 14952
rect 8478 14900 8484 14952
rect 8536 14940 8542 14952
rect 9232 14940 9260 14968
rect 10870 14940 10876 14952
rect 8536 14912 9260 14940
rect 9600 14912 10876 14940
rect 8536 14900 8542 14912
rect 6914 14832 6920 14884
rect 6972 14872 6978 14884
rect 9600 14872 9628 14912
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 11057 14943 11115 14949
rect 11057 14909 11069 14943
rect 11103 14940 11115 14943
rect 12066 14940 12072 14952
rect 11103 14912 12072 14940
rect 11103 14909 11115 14912
rect 11057 14903 11115 14909
rect 12066 14900 12072 14912
rect 12124 14900 12130 14952
rect 12434 14940 12440 14952
rect 12395 14912 12440 14940
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 13078 14900 13084 14952
rect 13136 14940 13142 14952
rect 13173 14943 13231 14949
rect 13173 14940 13185 14943
rect 13136 14912 13185 14940
rect 13136 14900 13142 14912
rect 13173 14909 13185 14912
rect 13219 14909 13231 14943
rect 13173 14903 13231 14909
rect 13909 14943 13967 14949
rect 13909 14909 13921 14943
rect 13955 14940 13967 14943
rect 15194 14940 15200 14952
rect 13955 14912 15200 14940
rect 13955 14909 13967 14912
rect 13909 14903 13967 14909
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 14458 14872 14464 14884
rect 6972 14844 9628 14872
rect 9692 14844 14464 14872
rect 6972 14832 6978 14844
rect 5534 14804 5540 14816
rect 4908 14776 5212 14804
rect 5495 14776 5540 14804
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 7282 14804 7288 14816
rect 7243 14776 7288 14804
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 8018 14804 8024 14816
rect 7979 14776 8024 14804
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 8662 14804 8668 14816
rect 8623 14776 8668 14804
rect 8662 14764 8668 14776
rect 8720 14764 8726 14816
rect 8846 14764 8852 14816
rect 8904 14804 8910 14816
rect 9033 14807 9091 14813
rect 9033 14804 9045 14807
rect 8904 14776 9045 14804
rect 8904 14764 8910 14776
rect 9033 14773 9045 14776
rect 9079 14773 9091 14807
rect 9033 14767 9091 14773
rect 9125 14807 9183 14813
rect 9125 14773 9137 14807
rect 9171 14804 9183 14807
rect 9692 14804 9720 14844
rect 14458 14832 14464 14844
rect 14516 14832 14522 14884
rect 9171 14776 9720 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 10134 14764 10140 14816
rect 10192 14804 10198 14816
rect 10229 14807 10287 14813
rect 10229 14804 10241 14807
rect 10192 14776 10241 14804
rect 10192 14764 10198 14776
rect 10229 14773 10241 14776
rect 10275 14773 10287 14807
rect 10229 14767 10287 14773
rect 11241 14807 11299 14813
rect 11241 14773 11253 14807
rect 11287 14804 11299 14807
rect 11514 14804 11520 14816
rect 11287 14776 11520 14804
rect 11287 14773 11299 14776
rect 11241 14767 11299 14773
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 1104 14714 15824 14736
rect 1104 14662 5912 14714
rect 5964 14662 5976 14714
rect 6028 14662 6040 14714
rect 6092 14662 6104 14714
rect 6156 14662 10843 14714
rect 10895 14662 10907 14714
rect 10959 14662 10971 14714
rect 11023 14662 11035 14714
rect 11087 14662 15824 14714
rect 1104 14640 15824 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 2682 14560 2688 14612
rect 2740 14600 2746 14612
rect 3234 14600 3240 14612
rect 2740 14572 3240 14600
rect 2740 14560 2746 14572
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 4157 14603 4215 14609
rect 4157 14569 4169 14603
rect 4203 14600 4215 14603
rect 4246 14600 4252 14612
rect 4203 14572 4252 14600
rect 4203 14569 4215 14572
rect 4157 14563 4215 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 4525 14603 4583 14609
rect 4525 14569 4537 14603
rect 4571 14600 4583 14603
rect 4571 14572 7236 14600
rect 4571 14569 4583 14572
rect 4525 14563 4583 14569
rect 1949 14535 2007 14541
rect 1949 14501 1961 14535
rect 1995 14532 2007 14535
rect 6546 14532 6552 14544
rect 1995 14504 6552 14532
rect 1995 14501 2007 14504
rect 1949 14495 2007 14501
rect 6546 14492 6552 14504
rect 6604 14492 6610 14544
rect 7208 14532 7236 14572
rect 7282 14560 7288 14612
rect 7340 14600 7346 14612
rect 12069 14603 12127 14609
rect 12069 14600 12081 14603
rect 7340 14572 12081 14600
rect 7340 14560 7346 14572
rect 12069 14569 12081 14572
rect 12115 14569 12127 14603
rect 12069 14563 12127 14569
rect 12342 14560 12348 14612
rect 12400 14600 12406 14612
rect 13265 14603 13323 14609
rect 13265 14600 13277 14603
rect 12400 14572 13277 14600
rect 12400 14560 12406 14572
rect 13265 14569 13277 14572
rect 13311 14569 13323 14603
rect 13265 14563 13323 14569
rect 10502 14532 10508 14544
rect 7208 14504 10508 14532
rect 10502 14492 10508 14504
rect 10560 14492 10566 14544
rect 12529 14535 12587 14541
rect 12529 14501 12541 14535
rect 12575 14532 12587 14535
rect 13078 14532 13084 14544
rect 12575 14504 13084 14532
rect 12575 14501 12587 14504
rect 12529 14495 12587 14501
rect 13078 14492 13084 14504
rect 13136 14492 13142 14544
rect 13170 14492 13176 14544
rect 13228 14532 13234 14544
rect 13633 14535 13691 14541
rect 13633 14532 13645 14535
rect 13228 14504 13645 14532
rect 13228 14492 13234 14504
rect 13633 14501 13645 14504
rect 13679 14532 13691 14535
rect 14918 14532 14924 14544
rect 13679 14504 14924 14532
rect 13679 14501 13691 14504
rect 13633 14495 13691 14501
rect 14918 14492 14924 14504
rect 14976 14492 14982 14544
rect 3142 14464 3148 14476
rect 3103 14436 3148 14464
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 4617 14467 4675 14473
rect 4617 14433 4629 14467
rect 4663 14464 4675 14467
rect 4706 14464 4712 14476
rect 4663 14436 4712 14464
rect 4663 14433 4675 14436
rect 4617 14427 4675 14433
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 5620 14467 5678 14473
rect 5620 14464 5632 14467
rect 4816 14436 5632 14464
rect 2038 14396 2044 14408
rect 1999 14368 2044 14396
rect 2038 14356 2044 14368
rect 2096 14356 2102 14408
rect 2130 14356 2136 14408
rect 2188 14396 2194 14408
rect 3234 14396 3240 14408
rect 2188 14368 2233 14396
rect 3195 14368 3240 14396
rect 2188 14356 2194 14368
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 4430 14396 4436 14408
rect 3467 14368 4436 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 4430 14356 4436 14368
rect 4488 14356 4494 14408
rect 4816 14405 4844 14436
rect 5620 14433 5632 14436
rect 5666 14464 5678 14467
rect 5902 14464 5908 14476
rect 5666 14436 5908 14464
rect 5666 14433 5678 14436
rect 5620 14427 5678 14433
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 7460 14467 7518 14473
rect 7460 14433 7472 14467
rect 7506 14464 7518 14467
rect 7834 14464 7840 14476
rect 7506 14436 7840 14464
rect 7506 14433 7518 14436
rect 7460 14427 7518 14433
rect 7834 14424 7840 14436
rect 7892 14424 7898 14476
rect 8202 14424 8208 14476
rect 8260 14464 8266 14476
rect 9217 14467 9275 14473
rect 9217 14464 9229 14467
rect 8260 14436 9229 14464
rect 8260 14424 8266 14436
rect 9217 14433 9229 14436
rect 9263 14433 9275 14467
rect 9217 14427 9275 14433
rect 9306 14424 9312 14476
rect 9364 14464 9370 14476
rect 10045 14467 10103 14473
rect 10045 14464 10057 14467
rect 9364 14436 10057 14464
rect 9364 14424 9370 14436
rect 10045 14433 10057 14436
rect 10091 14464 10103 14467
rect 10091 14436 11008 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 4801 14399 4859 14405
rect 4801 14365 4813 14399
rect 4847 14365 4859 14399
rect 4801 14359 4859 14365
rect 3786 14288 3792 14340
rect 3844 14328 3850 14340
rect 4816 14328 4844 14359
rect 4890 14356 4896 14408
rect 4948 14396 4954 14408
rect 5350 14396 5356 14408
rect 4948 14368 5356 14396
rect 4948 14356 4954 14368
rect 5350 14356 5356 14368
rect 5408 14356 5414 14408
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 7193 14399 7251 14405
rect 7193 14396 7205 14399
rect 6880 14368 7205 14396
rect 6880 14356 6886 14368
rect 7193 14365 7205 14368
rect 7239 14365 7251 14399
rect 9766 14396 9772 14408
rect 7193 14359 7251 14365
rect 8588 14368 9772 14396
rect 8588 14340 8616 14368
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 10134 14396 10140 14408
rect 10095 14368 10140 14396
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 8570 14328 8576 14340
rect 3844 14300 4844 14328
rect 6656 14300 7236 14328
rect 8531 14300 8576 14328
rect 3844 14288 3850 14300
rect 2777 14263 2835 14269
rect 2777 14229 2789 14263
rect 2823 14260 2835 14263
rect 6656 14260 6684 14300
rect 2823 14232 6684 14260
rect 2823 14229 2835 14232
rect 2777 14223 2835 14229
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 7006 14260 7012 14272
rect 6788 14232 7012 14260
rect 6788 14220 6794 14232
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7208 14260 7236 14300
rect 8570 14288 8576 14300
rect 8628 14288 8634 14340
rect 9674 14328 9680 14340
rect 9635 14300 9680 14328
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 10042 14288 10048 14340
rect 10100 14328 10106 14340
rect 10244 14328 10272 14359
rect 10100 14300 10272 14328
rect 10100 14288 10106 14300
rect 8202 14260 8208 14272
rect 7208 14232 8208 14260
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 8938 14220 8944 14272
rect 8996 14260 9002 14272
rect 9033 14263 9091 14269
rect 9033 14260 9045 14263
rect 8996 14232 9045 14260
rect 8996 14220 9002 14232
rect 9033 14229 9045 14232
rect 9079 14229 9091 14263
rect 9033 14223 9091 14229
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 10873 14263 10931 14269
rect 10873 14260 10885 14263
rect 9916 14232 10885 14260
rect 9916 14220 9922 14232
rect 10873 14229 10885 14232
rect 10919 14229 10931 14263
rect 10980 14260 11008 14436
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 11241 14467 11299 14473
rect 11241 14464 11253 14467
rect 11112 14436 11253 14464
rect 11112 14424 11118 14436
rect 11241 14433 11253 14436
rect 11287 14464 11299 14467
rect 11606 14464 11612 14476
rect 11287 14436 11612 14464
rect 11287 14433 11299 14436
rect 11241 14427 11299 14433
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 12710 14464 12716 14476
rect 12483 14436 12716 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 13538 14424 13544 14476
rect 13596 14464 13602 14476
rect 13725 14467 13783 14473
rect 13725 14464 13737 14467
rect 13596 14436 13737 14464
rect 13596 14424 13602 14436
rect 13725 14433 13737 14436
rect 13771 14433 13783 14467
rect 13725 14427 13783 14433
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14365 11391 14399
rect 11333 14359 11391 14365
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14396 11575 14399
rect 11882 14396 11888 14408
rect 11563 14368 11888 14396
rect 11563 14365 11575 14368
rect 11517 14359 11575 14365
rect 11348 14328 11376 14359
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 12342 14356 12348 14408
rect 12400 14396 12406 14408
rect 12621 14399 12679 14405
rect 12621 14396 12633 14399
rect 12400 14368 12633 14396
rect 12400 14356 12406 14368
rect 12621 14365 12633 14368
rect 12667 14365 12679 14399
rect 12621 14359 12679 14365
rect 13556 14328 13584 14424
rect 13814 14396 13820 14408
rect 13775 14368 13820 14396
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 11348 14300 13584 14328
rect 13170 14260 13176 14272
rect 10980 14232 13176 14260
rect 10873 14223 10931 14229
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 1104 14170 15824 14192
rect 1104 14118 3447 14170
rect 3499 14118 3511 14170
rect 3563 14118 3575 14170
rect 3627 14118 3639 14170
rect 3691 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 13308 14170
rect 13360 14118 13372 14170
rect 13424 14118 13436 14170
rect 13488 14118 13500 14170
rect 13552 14118 15824 14170
rect 1104 14096 15824 14118
rect 2498 14056 2504 14068
rect 2459 14028 2504 14056
rect 2498 14016 2504 14028
rect 2556 14016 2562 14068
rect 4062 14016 4068 14068
rect 4120 14056 4126 14068
rect 9306 14056 9312 14068
rect 4120 14028 8616 14056
rect 4120 14016 4126 14028
rect 8588 14000 8616 14028
rect 8680 14028 9312 14056
rect 2590 13948 2596 14000
rect 2648 13988 2654 14000
rect 3697 13991 3755 13997
rect 3697 13988 3709 13991
rect 2648 13960 3709 13988
rect 2648 13948 2654 13960
rect 3697 13957 3709 13960
rect 3743 13957 3755 13991
rect 3697 13951 3755 13957
rect 6273 13991 6331 13997
rect 6273 13957 6285 13991
rect 6319 13988 6331 13991
rect 6638 13988 6644 14000
rect 6319 13960 6644 13988
rect 6319 13957 6331 13960
rect 6273 13951 6331 13957
rect 6638 13948 6644 13960
rect 6696 13948 6702 14000
rect 8110 13948 8116 14000
rect 8168 13988 8174 14000
rect 8205 13991 8263 13997
rect 8205 13988 8217 13991
rect 8168 13960 8217 13988
rect 8168 13948 8174 13960
rect 8205 13957 8217 13960
rect 8251 13957 8263 13991
rect 8205 13951 8263 13957
rect 8570 13948 8576 14000
rect 8628 13948 8634 14000
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 3786 13920 3792 13932
rect 3191 13892 3792 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 3786 13880 3792 13892
rect 3844 13880 3850 13932
rect 4154 13920 4160 13932
rect 4115 13892 4160 13920
rect 4154 13880 4160 13892
rect 4212 13880 4218 13932
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4387 13892 5028 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13852 1915 13855
rect 2866 13852 2872 13864
rect 1903 13824 2872 13852
rect 1903 13821 1915 13824
rect 1857 13815 1915 13821
rect 2866 13812 2872 13824
rect 2924 13812 2930 13864
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13852 3019 13855
rect 4246 13852 4252 13864
rect 3007 13824 4252 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 4890 13852 4896 13864
rect 4851 13824 4896 13852
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 5000 13852 5028 13892
rect 6362 13880 6368 13932
rect 6420 13920 6426 13932
rect 6546 13920 6552 13932
rect 6420 13892 6552 13920
rect 6420 13880 6426 13892
rect 6546 13880 6552 13892
rect 6604 13880 6610 13932
rect 8478 13880 8484 13932
rect 8536 13920 8542 13932
rect 8680 13929 8708 14028
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 9398 14016 9404 14068
rect 9456 14056 9462 14068
rect 10502 14056 10508 14068
rect 9456 14028 9720 14056
rect 10463 14028 10508 14056
rect 9456 14016 9462 14028
rect 8665 13923 8723 13929
rect 8665 13920 8677 13923
rect 8536 13892 8677 13920
rect 8536 13880 8542 13892
rect 8665 13889 8677 13892
rect 8711 13889 8723 13923
rect 9692 13920 9720 14028
rect 10502 14016 10508 14028
rect 10560 14016 10566 14068
rect 11701 14059 11759 14065
rect 11701 14056 11713 14059
rect 10612 14028 11713 14056
rect 9950 13948 9956 14000
rect 10008 13988 10014 14000
rect 10045 13991 10103 13997
rect 10045 13988 10057 13991
rect 10008 13960 10057 13988
rect 10008 13948 10014 13960
rect 10045 13957 10057 13960
rect 10091 13957 10103 13991
rect 10045 13951 10103 13957
rect 10134 13948 10140 14000
rect 10192 13988 10198 14000
rect 10612 13988 10640 14028
rect 11701 14025 11713 14028
rect 11747 14025 11759 14059
rect 13814 14056 13820 14068
rect 11701 14019 11759 14025
rect 11788 14028 13820 14056
rect 11788 13988 11816 14028
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 10192 13960 10640 13988
rect 10704 13960 11816 13988
rect 10192 13948 10198 13960
rect 10704 13920 10732 13960
rect 12710 13948 12716 14000
rect 12768 13988 12774 14000
rect 13354 13988 13360 14000
rect 12768 13960 13360 13988
rect 12768 13948 12774 13960
rect 13354 13948 13360 13960
rect 13412 13948 13418 14000
rect 9692 13892 10732 13920
rect 11149 13923 11207 13929
rect 8665 13883 8723 13889
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 11330 13920 11336 13932
rect 11195 13892 11336 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 11330 13880 11336 13892
rect 11388 13880 11394 13932
rect 11606 13880 11612 13932
rect 11664 13920 11670 13932
rect 11664 13892 12020 13920
rect 11664 13880 11670 13892
rect 6270 13852 6276 13864
rect 5000 13824 6276 13852
rect 6270 13812 6276 13824
rect 6328 13812 6334 13864
rect 6822 13852 6828 13864
rect 6783 13824 6828 13852
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7024 13824 8340 13852
rect 5160 13787 5218 13793
rect 5160 13753 5172 13787
rect 5206 13784 5218 13787
rect 6362 13784 6368 13796
rect 5206 13756 6368 13784
rect 5206 13753 5218 13756
rect 5160 13747 5218 13753
rect 6362 13744 6368 13756
rect 6420 13744 6426 13796
rect 6454 13744 6460 13796
rect 6512 13784 6518 13796
rect 7024 13784 7052 13824
rect 6512 13756 7052 13784
rect 7092 13787 7150 13793
rect 6512 13744 6518 13756
rect 7092 13753 7104 13787
rect 7138 13784 7150 13787
rect 7374 13784 7380 13796
rect 7138 13756 7380 13784
rect 7138 13753 7150 13756
rect 7092 13747 7150 13753
rect 7374 13744 7380 13756
rect 7432 13784 7438 13796
rect 7742 13784 7748 13796
rect 7432 13756 7748 13784
rect 7432 13744 7438 13756
rect 7742 13744 7748 13756
rect 7800 13744 7806 13796
rect 8312 13784 8340 13824
rect 8680 13824 8953 13852
rect 8680 13784 8708 13824
rect 8925 13793 8953 13824
rect 9674 13812 9680 13864
rect 9732 13852 9738 13864
rect 9950 13852 9956 13864
rect 9732 13824 9956 13852
rect 9732 13812 9738 13824
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 10042 13812 10048 13864
rect 10100 13852 10106 13864
rect 10686 13852 10692 13864
rect 10100 13824 10692 13852
rect 10100 13812 10106 13824
rect 10686 13812 10692 13824
rect 10744 13812 10750 13864
rect 11882 13852 11888 13864
rect 11843 13824 11888 13852
rect 11882 13812 11888 13824
rect 11940 13812 11946 13864
rect 11992 13852 12020 13892
rect 12342 13880 12348 13932
rect 12400 13920 12406 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12400 13892 13001 13920
rect 12400 13880 12406 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 15562 13920 15568 13932
rect 12989 13883 13047 13889
rect 13556 13892 15568 13920
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 11992 13824 12817 13852
rect 12805 13821 12817 13824
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13852 12955 13855
rect 13262 13852 13268 13864
rect 12943 13824 13268 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 13262 13812 13268 13824
rect 13320 13852 13326 13864
rect 13556 13852 13584 13892
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 13320 13824 13584 13852
rect 13320 13812 13326 13824
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 13944 13855 14002 13861
rect 13944 13852 13956 13855
rect 13688 13824 13956 13852
rect 13688 13812 13694 13824
rect 13944 13821 13956 13824
rect 13990 13821 14002 13855
rect 13944 13815 14002 13821
rect 8312 13756 8708 13784
rect 8910 13787 8968 13793
rect 8910 13753 8922 13787
rect 8956 13753 8968 13787
rect 8910 13747 8968 13753
rect 9306 13744 9312 13796
rect 9364 13784 9370 13796
rect 9582 13784 9588 13796
rect 9364 13756 9588 13784
rect 9364 13744 9370 13756
rect 9582 13744 9588 13756
rect 9640 13784 9646 13796
rect 12250 13784 12256 13796
rect 9640 13756 12256 13784
rect 9640 13744 9646 13756
rect 12250 13744 12256 13756
rect 12308 13744 12314 13796
rect 16390 13784 16396 13796
rect 12348 13756 16396 13784
rect 2314 13676 2320 13728
rect 2372 13716 2378 13728
rect 2869 13719 2927 13725
rect 2869 13716 2881 13719
rect 2372 13688 2881 13716
rect 2372 13676 2378 13688
rect 2869 13685 2881 13688
rect 2915 13685 2927 13719
rect 2869 13679 2927 13685
rect 4065 13719 4123 13725
rect 4065 13685 4077 13719
rect 4111 13716 4123 13719
rect 9950 13716 9956 13728
rect 4111 13688 9956 13716
rect 4111 13685 4123 13688
rect 4065 13679 4123 13685
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 10686 13676 10692 13728
rect 10744 13716 10750 13728
rect 10873 13719 10931 13725
rect 10873 13716 10885 13719
rect 10744 13688 10885 13716
rect 10744 13676 10750 13688
rect 10873 13685 10885 13688
rect 10919 13685 10931 13719
rect 10873 13679 10931 13685
rect 10965 13719 11023 13725
rect 10965 13685 10977 13719
rect 11011 13716 11023 13719
rect 12348 13716 12376 13756
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 11011 13688 12376 13716
rect 11011 13685 11023 13688
rect 10965 13679 11023 13685
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12492 13688 12537 13716
rect 12492 13676 12498 13688
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 14047 13719 14105 13725
rect 14047 13716 14059 13719
rect 13872 13688 14059 13716
rect 13872 13676 13878 13688
rect 14047 13685 14059 13688
rect 14093 13685 14105 13719
rect 14047 13679 14105 13685
rect 1104 13626 15824 13648
rect 1104 13574 5912 13626
rect 5964 13574 5976 13626
rect 6028 13574 6040 13626
rect 6092 13574 6104 13626
rect 6156 13574 10843 13626
rect 10895 13574 10907 13626
rect 10959 13574 10971 13626
rect 11023 13574 11035 13626
rect 11087 13574 15824 13626
rect 1104 13552 15824 13574
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 3237 13515 3295 13521
rect 1995 13484 3188 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 2041 13447 2099 13453
rect 2041 13413 2053 13447
rect 2087 13444 2099 13447
rect 2222 13444 2228 13456
rect 2087 13416 2228 13444
rect 2087 13413 2099 13416
rect 2041 13407 2099 13413
rect 2222 13404 2228 13416
rect 2280 13404 2286 13456
rect 3160 13444 3188 13484
rect 3237 13481 3249 13515
rect 3283 13512 3295 13515
rect 4614 13512 4620 13524
rect 3283 13484 4620 13512
rect 3283 13481 3295 13484
rect 3237 13475 3295 13481
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 5074 13472 5080 13524
rect 5132 13512 5138 13524
rect 5350 13512 5356 13524
rect 5132 13484 5356 13512
rect 5132 13472 5138 13484
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 6362 13512 6368 13524
rect 6275 13484 6368 13512
rect 6362 13472 6368 13484
rect 6420 13512 6426 13524
rect 6914 13512 6920 13524
rect 6420 13484 6920 13512
rect 6420 13472 6426 13484
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7834 13512 7840 13524
rect 7156 13484 7840 13512
rect 7156 13472 7162 13484
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 8202 13512 8208 13524
rect 8163 13484 8208 13512
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 9490 13472 9496 13524
rect 9548 13512 9554 13524
rect 10502 13512 10508 13524
rect 9548 13484 10508 13512
rect 9548 13472 9554 13484
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 11885 13515 11943 13521
rect 11885 13481 11897 13515
rect 11931 13512 11943 13515
rect 11974 13512 11980 13524
rect 11931 13484 11980 13512
rect 11931 13481 11943 13484
rect 11885 13475 11943 13481
rect 11974 13472 11980 13484
rect 12032 13472 12038 13524
rect 12250 13472 12256 13524
rect 12308 13512 12314 13524
rect 12713 13515 12771 13521
rect 12713 13512 12725 13515
rect 12308 13484 12725 13512
rect 12308 13472 12314 13484
rect 12713 13481 12725 13484
rect 12759 13481 12771 13515
rect 13906 13512 13912 13524
rect 12713 13475 12771 13481
rect 12820 13484 13912 13512
rect 3786 13444 3792 13456
rect 3160 13416 3792 13444
rect 3786 13404 3792 13416
rect 3844 13404 3850 13456
rect 12618 13444 12624 13456
rect 4080 13416 12624 13444
rect 2498 13336 2504 13388
rect 2556 13376 2562 13388
rect 2682 13376 2688 13388
rect 2556 13348 2688 13376
rect 2556 13336 2562 13348
rect 2682 13336 2688 13348
rect 2740 13376 2746 13388
rect 4080 13385 4108 13416
rect 12618 13404 12624 13416
rect 12676 13404 12682 13456
rect 3145 13379 3203 13385
rect 3145 13376 3157 13379
rect 2740 13348 3157 13376
rect 2740 13336 2746 13348
rect 3145 13345 3157 13348
rect 3191 13345 3203 13379
rect 3145 13339 3203 13345
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13345 4123 13379
rect 4065 13339 4123 13345
rect 4614 13336 4620 13388
rect 4672 13376 4678 13388
rect 7098 13385 7104 13388
rect 5241 13379 5299 13385
rect 5241 13376 5253 13379
rect 4672 13348 5253 13376
rect 4672 13336 4678 13348
rect 5241 13345 5253 13348
rect 5287 13345 5299 13379
rect 7092 13376 7104 13385
rect 7059 13348 7104 13376
rect 5241 13339 5299 13345
rect 7092 13339 7104 13348
rect 7098 13336 7104 13339
rect 7156 13336 7162 13388
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 8665 13379 8723 13385
rect 8665 13376 8677 13379
rect 8352 13348 8677 13376
rect 8352 13336 8358 13348
rect 8665 13345 8677 13348
rect 8711 13345 8723 13379
rect 8665 13339 8723 13345
rect 9582 13336 9588 13388
rect 9640 13376 9646 13388
rect 9677 13379 9735 13385
rect 9677 13376 9689 13379
rect 9640 13348 9689 13376
rect 9640 13336 9646 13348
rect 9677 13345 9689 13348
rect 9723 13345 9735 13379
rect 9677 13339 9735 13345
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 9933 13379 9991 13385
rect 9933 13376 9945 13379
rect 9824 13348 9945 13376
rect 9824 13336 9830 13348
rect 9933 13345 9945 13348
rect 9979 13345 9991 13379
rect 9933 13339 9991 13345
rect 10502 13336 10508 13388
rect 10560 13376 10566 13388
rect 10560 13348 10732 13376
rect 10560 13336 10566 13348
rect 1486 13268 1492 13320
rect 1544 13308 1550 13320
rect 2133 13311 2191 13317
rect 2133 13308 2145 13311
rect 1544 13280 2145 13308
rect 1544 13268 1550 13280
rect 2133 13277 2145 13280
rect 2179 13277 2191 13311
rect 2133 13271 2191 13277
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13277 3479 13311
rect 4246 13308 4252 13320
rect 4207 13280 4252 13308
rect 3421 13271 3479 13277
rect 1581 13243 1639 13249
rect 1581 13209 1593 13243
rect 1627 13240 1639 13243
rect 2406 13240 2412 13252
rect 1627 13212 2412 13240
rect 1627 13209 1639 13212
rect 1581 13203 1639 13209
rect 2406 13200 2412 13212
rect 2464 13200 2470 13252
rect 2774 13200 2780 13252
rect 2832 13240 2838 13252
rect 2832 13212 2877 13240
rect 2832 13200 2838 13212
rect 1854 13132 1860 13184
rect 1912 13172 1918 13184
rect 3234 13172 3240 13184
rect 1912 13144 3240 13172
rect 1912 13132 1918 13144
rect 3234 13132 3240 13144
rect 3292 13132 3298 13184
rect 3436 13172 3464 13271
rect 4246 13268 4252 13280
rect 4304 13268 4310 13320
rect 4890 13268 4896 13320
rect 4948 13308 4954 13320
rect 4985 13311 5043 13317
rect 4985 13308 4997 13311
rect 4948 13280 4997 13308
rect 4948 13268 4954 13280
rect 4985 13277 4997 13280
rect 5031 13277 5043 13311
rect 6822 13308 6828 13320
rect 6783 13280 6828 13308
rect 4985 13271 5043 13277
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 8846 13308 8852 13320
rect 8807 13280 8852 13308
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 10704 13308 10732 13348
rect 11514 13336 11520 13388
rect 11572 13376 11578 13388
rect 11977 13379 12035 13385
rect 11977 13376 11989 13379
rect 11572 13348 11989 13376
rect 11572 13336 11578 13348
rect 11977 13345 11989 13348
rect 12023 13376 12035 13379
rect 12820 13376 12848 13484
rect 13906 13472 13912 13484
rect 13964 13512 13970 13524
rect 14826 13512 14832 13524
rect 13964 13484 14832 13512
rect 13964 13472 13970 13484
rect 14826 13472 14832 13484
rect 14884 13472 14890 13524
rect 13814 13444 13820 13456
rect 13775 13416 13820 13444
rect 13814 13404 13820 13416
rect 13872 13404 13878 13456
rect 12023 13348 12848 13376
rect 12897 13379 12955 13385
rect 12023 13345 12035 13348
rect 11977 13339 12035 13345
rect 12897 13345 12909 13379
rect 12943 13376 12955 13379
rect 13262 13376 13268 13388
rect 12943 13348 13268 13376
rect 12943 13345 12955 13348
rect 12897 13339 12955 13345
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 12069 13311 12127 13317
rect 12069 13308 12081 13311
rect 10704 13280 12081 13308
rect 12069 13277 12081 13280
rect 12115 13308 12127 13311
rect 12342 13308 12348 13320
rect 12115 13280 12348 13308
rect 12115 13277 12127 13280
rect 12069 13271 12127 13277
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 13722 13308 13728 13320
rect 13683 13280 13728 13308
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 13998 13308 14004 13320
rect 13959 13280 14004 13308
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 7834 13200 7840 13252
rect 7892 13240 7898 13252
rect 9674 13240 9680 13252
rect 7892 13212 9680 13240
rect 7892 13200 7898 13212
rect 9674 13200 9680 13212
rect 9732 13200 9738 13252
rect 11054 13240 11060 13252
rect 11015 13212 11060 13240
rect 11054 13200 11060 13212
rect 11112 13200 11118 13252
rect 13814 13240 13820 13252
rect 11348 13212 13820 13240
rect 6638 13172 6644 13184
rect 3436 13144 6644 13172
rect 6638 13132 6644 13144
rect 6696 13132 6702 13184
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 11348 13172 11376 13212
rect 13814 13200 13820 13212
rect 13872 13200 13878 13252
rect 11514 13172 11520 13184
rect 7248 13144 11376 13172
rect 11475 13144 11520 13172
rect 7248 13132 7254 13144
rect 11514 13132 11520 13144
rect 11572 13132 11578 13184
rect 1104 13082 15824 13104
rect 1104 13030 3447 13082
rect 3499 13030 3511 13082
rect 3563 13030 3575 13082
rect 3627 13030 3639 13082
rect 3691 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 13308 13082
rect 13360 13030 13372 13082
rect 13424 13030 13436 13082
rect 13488 13030 13500 13082
rect 13552 13030 15824 13082
rect 1104 13008 15824 13030
rect 1854 12968 1860 12980
rect 1815 12940 1860 12968
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 2222 12928 2228 12980
rect 2280 12968 2286 12980
rect 4154 12968 4160 12980
rect 2280 12940 4160 12968
rect 2280 12928 2286 12940
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 4430 12968 4436 12980
rect 4391 12940 4436 12968
rect 4430 12928 4436 12940
rect 4488 12928 4494 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 4580 12940 6837 12968
rect 4580 12928 4586 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 9122 12968 9128 12980
rect 6825 12931 6883 12937
rect 7208 12940 9128 12968
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12801 2559 12835
rect 3050 12832 3056 12844
rect 3011 12804 3056 12832
rect 2501 12795 2559 12801
rect 2516 12764 2544 12795
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 4706 12792 4712 12844
rect 4764 12832 4770 12844
rect 4890 12832 4896 12844
rect 4764 12804 4896 12832
rect 4764 12792 4770 12804
rect 4890 12792 4896 12804
rect 4948 12792 4954 12844
rect 2516 12736 3363 12764
rect 3335 12705 3363 12736
rect 4430 12724 4436 12776
rect 4488 12764 4494 12776
rect 5149 12767 5207 12773
rect 5149 12764 5161 12767
rect 4488 12736 5161 12764
rect 4488 12724 4494 12736
rect 5149 12733 5161 12736
rect 5195 12733 5207 12767
rect 5149 12727 5207 12733
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 7208 12773 7236 12940
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9582 12928 9588 12980
rect 9640 12968 9646 12980
rect 9640 12940 9904 12968
rect 9640 12928 9646 12940
rect 7650 12860 7656 12912
rect 7708 12900 7714 12912
rect 8294 12900 8300 12912
rect 7708 12872 8300 12900
rect 7708 12860 7714 12872
rect 8294 12860 8300 12872
rect 8352 12860 8358 12912
rect 8386 12860 8392 12912
rect 8444 12900 8450 12912
rect 9766 12900 9772 12912
rect 8444 12872 9772 12900
rect 8444 12860 8450 12872
rect 9766 12860 9772 12872
rect 9824 12860 9830 12912
rect 9876 12900 9904 12940
rect 9950 12928 9956 12980
rect 10008 12968 10014 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 10008 12940 10609 12968
rect 10008 12928 10014 12940
rect 10597 12937 10609 12940
rect 10643 12937 10655 12971
rect 10597 12931 10655 12937
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 12986 12968 12992 12980
rect 11112 12940 12992 12968
rect 11112 12928 11118 12940
rect 12986 12928 12992 12940
rect 13044 12928 13050 12980
rect 13078 12928 13084 12980
rect 13136 12968 13142 12980
rect 13633 12971 13691 12977
rect 13633 12968 13645 12971
rect 13136 12940 13645 12968
rect 13136 12928 13142 12940
rect 13633 12937 13645 12940
rect 13679 12937 13691 12971
rect 13633 12931 13691 12937
rect 12437 12903 12495 12909
rect 12437 12900 12449 12903
rect 9876 12872 12449 12900
rect 12437 12869 12449 12872
rect 12483 12869 12495 12903
rect 12437 12863 12495 12869
rect 12618 12860 12624 12912
rect 12676 12900 12682 12912
rect 12676 12872 13032 12900
rect 12676 12860 12682 12872
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12832 7527 12835
rect 7834 12832 7840 12844
rect 7515 12804 7840 12832
rect 7515 12801 7527 12804
rect 7469 12795 7527 12801
rect 7834 12792 7840 12804
rect 7892 12792 7898 12844
rect 7926 12792 7932 12844
rect 7984 12832 7990 12844
rect 9030 12832 9036 12844
rect 7984 12804 8953 12832
rect 8991 12804 9036 12832
rect 7984 12792 7990 12804
rect 7193 12767 7251 12773
rect 7193 12764 7205 12767
rect 5500 12736 7205 12764
rect 5500 12724 5506 12736
rect 7193 12733 7205 12736
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 7374 12724 7380 12776
rect 7432 12764 7438 12776
rect 8297 12767 8355 12773
rect 8297 12764 8309 12767
rect 7432 12736 8309 12764
rect 7432 12724 7438 12736
rect 8297 12733 8309 12736
rect 8343 12733 8355 12767
rect 8297 12727 8355 12733
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 8925 12764 8953 12804
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 11149 12835 11207 12841
rect 11149 12832 11161 12835
rect 10928 12804 11161 12832
rect 10928 12792 10934 12804
rect 11149 12801 11161 12804
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 11514 12792 11520 12844
rect 11572 12832 11578 12844
rect 13004 12841 13032 12872
rect 12897 12835 12955 12841
rect 12897 12832 12909 12835
rect 11572 12804 12909 12832
rect 11572 12792 11578 12804
rect 12897 12801 12909 12804
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13872 12804 14197 12832
rect 13872 12792 13878 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 9582 12764 9588 12776
rect 8444 12736 8489 12764
rect 8925 12736 9588 12764
rect 8444 12724 8450 12736
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 9674 12724 9680 12776
rect 9732 12764 9738 12776
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 9732 12736 10517 12764
rect 9732 12724 9738 12736
rect 10505 12733 10517 12736
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 10594 12724 10600 12776
rect 10652 12764 10658 12776
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 10652 12736 10977 12764
rect 10652 12724 10658 12736
rect 10965 12733 10977 12736
rect 11011 12733 11023 12767
rect 11977 12767 12035 12773
rect 11977 12764 11989 12767
rect 10965 12727 11023 12733
rect 11164 12736 11989 12764
rect 3320 12699 3378 12705
rect 3320 12665 3332 12699
rect 3366 12696 3378 12699
rect 3418 12696 3424 12708
rect 3366 12668 3424 12696
rect 3366 12665 3378 12668
rect 3320 12659 3378 12665
rect 3418 12656 3424 12668
rect 3476 12656 3482 12708
rect 3786 12656 3792 12708
rect 3844 12696 3850 12708
rect 7285 12699 7343 12705
rect 7285 12696 7297 12699
rect 3844 12668 7297 12696
rect 3844 12656 3850 12668
rect 7285 12665 7297 12668
rect 7331 12696 7343 12699
rect 7926 12696 7932 12708
rect 7331 12668 7932 12696
rect 7331 12665 7343 12668
rect 7285 12659 7343 12665
rect 7926 12656 7932 12668
rect 7984 12656 7990 12708
rect 8938 12696 8944 12708
rect 8128 12668 8944 12696
rect 1946 12588 1952 12640
rect 2004 12628 2010 12640
rect 2225 12631 2283 12637
rect 2225 12628 2237 12631
rect 2004 12600 2237 12628
rect 2004 12588 2010 12600
rect 2225 12597 2237 12600
rect 2271 12597 2283 12631
rect 2225 12591 2283 12597
rect 2317 12631 2375 12637
rect 2317 12597 2329 12631
rect 2363 12628 2375 12631
rect 4338 12628 4344 12640
rect 2363 12600 4344 12628
rect 2363 12597 2375 12600
rect 2317 12591 2375 12597
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 5718 12588 5724 12640
rect 5776 12628 5782 12640
rect 6273 12631 6331 12637
rect 6273 12628 6285 12631
rect 5776 12600 6285 12628
rect 5776 12588 5782 12600
rect 6273 12597 6285 12600
rect 6319 12628 6331 12631
rect 6914 12628 6920 12640
rect 6319 12600 6920 12628
rect 6319 12597 6331 12600
rect 6273 12591 6331 12597
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 8128 12637 8156 12668
rect 8938 12656 8944 12668
rect 8996 12696 9002 12708
rect 8996 12668 10640 12696
rect 8996 12656 9002 12668
rect 8113 12631 8171 12637
rect 8113 12597 8125 12631
rect 8159 12597 8171 12631
rect 8113 12591 8171 12597
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 9214 12628 9220 12640
rect 8260 12600 9220 12628
rect 8260 12588 8266 12600
rect 9214 12588 9220 12600
rect 9272 12588 9278 12640
rect 9677 12631 9735 12637
rect 9677 12597 9689 12631
rect 9723 12628 9735 12631
rect 9766 12628 9772 12640
rect 9723 12600 9772 12628
rect 9723 12597 9735 12600
rect 9677 12591 9735 12597
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 10008 12600 10333 12628
rect 10008 12588 10014 12600
rect 10321 12597 10333 12600
rect 10367 12597 10379 12631
rect 10612 12628 10640 12668
rect 10686 12656 10692 12708
rect 10744 12696 10750 12708
rect 11057 12699 11115 12705
rect 11057 12696 11069 12699
rect 10744 12668 11069 12696
rect 10744 12656 10750 12668
rect 11057 12665 11069 12668
rect 11103 12665 11115 12699
rect 11057 12659 11115 12665
rect 11164 12628 11192 12736
rect 11977 12733 11989 12736
rect 12023 12733 12035 12767
rect 11977 12727 12035 12733
rect 12066 12724 12072 12776
rect 12124 12764 12130 12776
rect 12342 12764 12348 12776
rect 12124 12736 12348 12764
rect 12124 12724 12130 12736
rect 12342 12724 12348 12736
rect 12400 12724 12406 12776
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12492 12736 12817 12764
rect 12492 12724 12498 12736
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 13630 12656 13636 12708
rect 13688 12696 13694 12708
rect 14093 12699 14151 12705
rect 14093 12696 14105 12699
rect 13688 12668 14105 12696
rect 13688 12656 13694 12668
rect 14093 12665 14105 12668
rect 14139 12665 14151 12699
rect 14093 12659 14151 12665
rect 10612 12600 11192 12628
rect 10321 12591 10379 12597
rect 11514 12588 11520 12640
rect 11572 12628 11578 12640
rect 11793 12631 11851 12637
rect 11793 12628 11805 12631
rect 11572 12600 11805 12628
rect 11572 12588 11578 12600
rect 11793 12597 11805 12600
rect 11839 12597 11851 12631
rect 11793 12591 11851 12597
rect 13078 12588 13084 12640
rect 13136 12628 13142 12640
rect 14001 12631 14059 12637
rect 14001 12628 14013 12631
rect 13136 12600 14013 12628
rect 13136 12588 13142 12600
rect 14001 12597 14013 12600
rect 14047 12597 14059 12631
rect 14001 12591 14059 12597
rect 1104 12538 15824 12560
rect 1104 12486 5912 12538
rect 5964 12486 5976 12538
rect 6028 12486 6040 12538
rect 6092 12486 6104 12538
rect 6156 12486 10843 12538
rect 10895 12486 10907 12538
rect 10959 12486 10971 12538
rect 11023 12486 11035 12538
rect 11087 12486 15824 12538
rect 1104 12464 15824 12486
rect 1578 12384 1584 12436
rect 1636 12424 1642 12436
rect 1673 12427 1731 12433
rect 1673 12424 1685 12427
rect 1636 12396 1685 12424
rect 1636 12384 1642 12396
rect 1673 12393 1685 12396
rect 1719 12393 1731 12427
rect 1673 12387 1731 12393
rect 2041 12427 2099 12433
rect 2041 12393 2053 12427
rect 2087 12424 2099 12427
rect 5718 12424 5724 12436
rect 2087 12396 5724 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 5718 12384 5724 12396
rect 5776 12384 5782 12436
rect 6089 12427 6147 12433
rect 6089 12393 6101 12427
rect 6135 12424 6147 12427
rect 6454 12424 6460 12436
rect 6135 12396 6460 12424
rect 6135 12393 6147 12396
rect 6089 12387 6147 12393
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 6549 12427 6607 12433
rect 6549 12393 6561 12427
rect 6595 12393 6607 12427
rect 6549 12387 6607 12393
rect 4065 12359 4123 12365
rect 4065 12325 4077 12359
rect 4111 12356 4123 12359
rect 4341 12359 4399 12365
rect 4341 12356 4353 12359
rect 4111 12328 4353 12356
rect 4111 12325 4123 12328
rect 4065 12319 4123 12325
rect 4341 12325 4353 12328
rect 4387 12356 4399 12359
rect 6362 12356 6368 12368
rect 4387 12328 6368 12356
rect 4387 12325 4399 12328
rect 4341 12319 4399 12325
rect 6362 12316 6368 12328
rect 6420 12316 6426 12368
rect 6564 12356 6592 12387
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7190 12424 7196 12436
rect 6972 12396 7196 12424
rect 6972 12384 6978 12396
rect 7190 12384 7196 12396
rect 7248 12424 7254 12436
rect 7374 12424 7380 12436
rect 7248 12396 7380 12424
rect 7248 12384 7254 12396
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 7469 12427 7527 12433
rect 7469 12393 7481 12427
rect 7515 12424 7527 12427
rect 8478 12424 8484 12436
rect 7515 12396 8484 12424
rect 7515 12393 7527 12396
rect 7469 12387 7527 12393
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 8757 12427 8815 12433
rect 8757 12393 8769 12427
rect 8803 12424 8815 12427
rect 8846 12424 8852 12436
rect 8803 12396 8852 12424
rect 8803 12393 8815 12396
rect 8757 12387 8815 12393
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 9306 12424 9312 12436
rect 9140 12396 9312 12424
rect 8202 12356 8208 12368
rect 6564 12328 8208 12356
rect 2682 12288 2688 12300
rect 2643 12260 2688 12288
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 4706 12288 4712 12300
rect 4667 12260 4712 12288
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 4976 12291 5034 12297
rect 4976 12257 4988 12291
rect 5022 12288 5034 12291
rect 5258 12288 5264 12300
rect 5022 12260 5264 12288
rect 5022 12257 5034 12260
rect 4976 12251 5034 12257
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 6564 12232 6592 12328
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 8662 12356 8668 12368
rect 8623 12328 8668 12356
rect 8662 12316 8668 12328
rect 8720 12356 8726 12368
rect 9140 12356 9168 12396
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 10042 12424 10048 12436
rect 9723 12396 10048 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 10873 12427 10931 12433
rect 10873 12424 10885 12427
rect 10744 12396 10885 12424
rect 10744 12384 10750 12396
rect 10873 12393 10885 12396
rect 10919 12393 10931 12427
rect 10873 12387 10931 12393
rect 11241 12427 11299 12433
rect 11241 12393 11253 12427
rect 11287 12424 11299 12427
rect 15194 12424 15200 12436
rect 11287 12396 15200 12424
rect 11287 12393 11299 12396
rect 11241 12387 11299 12393
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 8720 12328 9168 12356
rect 8720 12316 8726 12328
rect 9214 12316 9220 12368
rect 9272 12356 9278 12368
rect 9272 12328 10456 12356
rect 9272 12316 9278 12328
rect 6730 12288 6736 12300
rect 6691 12260 6736 12288
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 8570 12288 8576 12300
rect 7116 12260 8576 12288
rect 2130 12220 2136 12232
rect 2091 12192 2136 12220
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 3329 12223 3387 12229
rect 2363 12192 3280 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 3252 12084 3280 12192
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 3344 12152 3372 12183
rect 6546 12180 6552 12232
rect 6604 12180 6610 12232
rect 7116 12161 7144 12260
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 8754 12248 8760 12300
rect 8812 12288 8818 12300
rect 9766 12288 9772 12300
rect 8812 12260 9772 12288
rect 8812 12248 8818 12260
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 10226 12288 10232 12300
rect 10100 12260 10232 12288
rect 10100 12248 10106 12260
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 10428 12297 10456 12328
rect 10962 12316 10968 12368
rect 11020 12356 11026 12368
rect 11020 12328 12020 12356
rect 11020 12316 11026 12328
rect 10413 12291 10471 12297
rect 10413 12257 10425 12291
rect 10459 12257 10471 12291
rect 10413 12251 10471 12257
rect 10781 12291 10839 12297
rect 10781 12257 10793 12291
rect 10827 12288 10839 12291
rect 11330 12288 11336 12300
rect 10827 12260 11336 12288
rect 10827 12257 10839 12260
rect 10781 12251 10839 12257
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 11882 12288 11888 12300
rect 11532 12260 11888 12288
rect 7561 12223 7619 12229
rect 7561 12189 7573 12223
rect 7607 12189 7619 12223
rect 7561 12183 7619 12189
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 7834 12220 7840 12232
rect 7791 12192 7840 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 7101 12155 7159 12161
rect 3344 12124 4752 12152
rect 4154 12084 4160 12096
rect 3252 12056 4160 12084
rect 4154 12044 4160 12056
rect 4212 12044 4218 12096
rect 4724 12084 4752 12124
rect 7101 12121 7113 12155
rect 7147 12121 7159 12155
rect 7101 12115 7159 12121
rect 7006 12084 7012 12096
rect 4724 12056 7012 12084
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 7576 12084 7604 12183
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 8294 12220 8300 12232
rect 7944 12192 8300 12220
rect 7524 12056 7604 12084
rect 7524 12044 7530 12056
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 7944 12084 7972 12192
rect 8294 12180 8300 12192
rect 8352 12220 8358 12232
rect 8941 12223 8999 12229
rect 8941 12220 8953 12223
rect 8352 12192 8953 12220
rect 8352 12180 8358 12192
rect 8941 12189 8953 12192
rect 8987 12220 8999 12223
rect 9493 12223 9551 12229
rect 8987 12192 9444 12220
rect 8987 12189 8999 12192
rect 8941 12183 8999 12189
rect 8018 12112 8024 12164
rect 8076 12152 8082 12164
rect 9416 12152 9444 12192
rect 9493 12189 9505 12223
rect 9539 12220 9551 12223
rect 11425 12223 11483 12229
rect 11425 12220 11437 12223
rect 9539 12192 11437 12220
rect 9539 12189 9551 12192
rect 9493 12183 9551 12189
rect 11425 12189 11437 12192
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 10229 12155 10287 12161
rect 8076 12124 9076 12152
rect 9416 12124 9628 12152
rect 8076 12112 8082 12124
rect 7800 12056 7972 12084
rect 7800 12044 7806 12056
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8297 12087 8355 12093
rect 8297 12084 8309 12087
rect 8260 12056 8309 12084
rect 8260 12044 8266 12056
rect 8297 12053 8309 12056
rect 8343 12053 8355 12087
rect 9048 12084 9076 12124
rect 9122 12084 9128 12096
rect 9048 12056 9128 12084
rect 8297 12047 8355 12053
rect 9122 12044 9128 12056
rect 9180 12084 9186 12096
rect 9493 12087 9551 12093
rect 9493 12084 9505 12087
rect 9180 12056 9505 12084
rect 9180 12044 9186 12056
rect 9493 12053 9505 12056
rect 9539 12053 9551 12087
rect 9600 12084 9628 12124
rect 10229 12121 10241 12155
rect 10275 12152 10287 12155
rect 11532 12152 11560 12260
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 11992 12288 12020 12328
rect 12158 12316 12164 12368
rect 12216 12356 12222 12368
rect 13262 12356 13268 12368
rect 12216 12328 13268 12356
rect 12216 12316 12222 12328
rect 13262 12316 13268 12328
rect 13320 12356 13326 12368
rect 13633 12359 13691 12365
rect 13633 12356 13645 12359
rect 13320 12328 13645 12356
rect 13320 12316 13326 12328
rect 13633 12325 13645 12328
rect 13679 12325 13691 12359
rect 13633 12319 13691 12325
rect 12437 12291 12495 12297
rect 12437 12288 12449 12291
rect 11992 12260 12449 12288
rect 12437 12257 12449 12260
rect 12483 12257 12495 12291
rect 12437 12251 12495 12257
rect 12529 12291 12587 12297
rect 12529 12257 12541 12291
rect 12575 12288 12587 12291
rect 12802 12288 12808 12300
rect 12575 12260 12808 12288
rect 12575 12257 12587 12260
rect 12529 12251 12587 12257
rect 12802 12248 12808 12260
rect 12860 12288 12866 12300
rect 14274 12288 14280 12300
rect 12860 12260 14280 12288
rect 12860 12248 12866 12260
rect 14274 12248 14280 12260
rect 14332 12248 14338 12300
rect 12618 12220 12624 12232
rect 12579 12192 12624 12220
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 12894 12180 12900 12232
rect 12952 12220 12958 12232
rect 13725 12223 13783 12229
rect 13725 12220 13737 12223
rect 12952 12192 13737 12220
rect 12952 12180 12958 12192
rect 13725 12189 13737 12192
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 13817 12223 13875 12229
rect 13817 12189 13829 12223
rect 13863 12189 13875 12223
rect 13817 12183 13875 12189
rect 10275 12124 11560 12152
rect 11624 12124 12376 12152
rect 10275 12121 10287 12124
rect 10229 12115 10287 12121
rect 11624 12084 11652 12124
rect 9600 12056 11652 12084
rect 12069 12087 12127 12093
rect 9493 12047 9551 12053
rect 12069 12053 12081 12087
rect 12115 12084 12127 12087
rect 12250 12084 12256 12096
rect 12115 12056 12256 12084
rect 12115 12053 12127 12056
rect 12069 12047 12127 12053
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 12348 12084 12376 12124
rect 12802 12112 12808 12164
rect 12860 12152 12866 12164
rect 13265 12155 13323 12161
rect 13265 12152 13277 12155
rect 12860 12124 13277 12152
rect 12860 12112 12866 12124
rect 13265 12121 13277 12124
rect 13311 12121 13323 12155
rect 13265 12115 13323 12121
rect 13832 12084 13860 12183
rect 12348 12056 13860 12084
rect 1104 11994 15824 12016
rect 1104 11942 3447 11994
rect 3499 11942 3511 11994
rect 3563 11942 3575 11994
rect 3627 11942 3639 11994
rect 3691 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 13308 11994
rect 13360 11942 13372 11994
rect 13424 11942 13436 11994
rect 13488 11942 13500 11994
rect 13552 11942 15824 11994
rect 1104 11920 15824 11942
rect 3234 11880 3240 11892
rect 3068 11852 3240 11880
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 2314 11608 2320 11620
rect 2275 11580 2320 11608
rect 2314 11568 2320 11580
rect 2372 11568 2378 11620
rect 2516 11608 2544 11707
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 3068 11753 3096 11852
rect 3234 11840 3240 11852
rect 3292 11840 3298 11892
rect 4433 11883 4491 11889
rect 4433 11849 4445 11883
rect 4479 11880 4491 11883
rect 7834 11880 7840 11892
rect 4479 11852 7840 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 7834 11840 7840 11852
rect 7892 11880 7898 11892
rect 7892 11852 9720 11880
rect 7892 11840 7898 11852
rect 3053 11747 3111 11753
rect 3053 11744 3065 11747
rect 2832 11716 3065 11744
rect 2832 11704 2838 11716
rect 3053 11713 3065 11716
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4764 11716 4905 11744
rect 4764 11704 4770 11716
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 6822 11744 6828 11756
rect 6783 11716 6828 11744
rect 4893 11707 4951 11713
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 9692 11744 9720 11852
rect 10502 11840 10508 11892
rect 10560 11880 10566 11892
rect 10870 11880 10876 11892
rect 10560 11852 10876 11880
rect 10560 11840 10566 11852
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 12437 11883 12495 11889
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 12710 11880 12716 11892
rect 12483 11852 12716 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 9858 11772 9864 11824
rect 9916 11812 9922 11824
rect 9916 11784 14228 11812
rect 9916 11772 9922 11784
rect 11057 11747 11115 11753
rect 11057 11744 11069 11747
rect 7852 11716 8800 11744
rect 9692 11716 11069 11744
rect 3320 11679 3378 11685
rect 3320 11645 3332 11679
rect 3366 11676 3378 11679
rect 3366 11648 5672 11676
rect 3366 11645 3378 11648
rect 3320 11639 3378 11645
rect 5644 11620 5672 11648
rect 6638 11636 6644 11688
rect 6696 11676 6702 11688
rect 7081 11679 7139 11685
rect 7081 11676 7093 11679
rect 6696 11648 7093 11676
rect 6696 11636 6702 11648
rect 7081 11645 7093 11648
rect 7127 11645 7139 11679
rect 7852 11676 7880 11716
rect 7081 11639 7139 11645
rect 7300 11648 7880 11676
rect 3418 11608 3424 11620
rect 2516 11580 3424 11608
rect 3418 11568 3424 11580
rect 3476 11568 3482 11620
rect 5160 11611 5218 11617
rect 5160 11577 5172 11611
rect 5206 11608 5218 11611
rect 5350 11608 5356 11620
rect 5206 11580 5356 11608
rect 5206 11577 5218 11580
rect 5160 11571 5218 11577
rect 5350 11568 5356 11580
rect 5408 11568 5414 11620
rect 5626 11568 5632 11620
rect 5684 11608 5690 11620
rect 7190 11608 7196 11620
rect 5684 11580 7196 11608
rect 5684 11568 5690 11580
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 1857 11543 1915 11549
rect 1857 11509 1869 11543
rect 1903 11540 1915 11543
rect 2038 11540 2044 11552
rect 1903 11512 2044 11540
rect 1903 11509 1915 11512
rect 1857 11503 1915 11509
rect 2038 11500 2044 11512
rect 2096 11500 2102 11552
rect 2225 11543 2283 11549
rect 2225 11509 2237 11543
rect 2271 11540 2283 11543
rect 2682 11540 2688 11552
rect 2271 11512 2688 11540
rect 2271 11509 2283 11512
rect 2225 11503 2283 11509
rect 2682 11500 2688 11512
rect 2740 11500 2746 11552
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 6273 11543 6331 11549
rect 6273 11540 6285 11543
rect 4672 11512 6285 11540
rect 4672 11500 4678 11512
rect 6273 11509 6285 11512
rect 6319 11509 6331 11543
rect 6273 11503 6331 11509
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7300 11540 7328 11648
rect 8294 11636 8300 11688
rect 8352 11676 8358 11688
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 8352 11648 8677 11676
rect 8352 11636 8358 11648
rect 8665 11645 8677 11648
rect 8711 11645 8723 11679
rect 8772 11676 8800 11716
rect 11057 11713 11069 11716
rect 11103 11713 11115 11747
rect 11057 11707 11115 11713
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 14200 11753 14228 11784
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 11664 11716 13001 11744
rect 11664 11704 11670 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 15470 11744 15476 11756
rect 14792 11716 15476 11744
rect 14792 11704 14798 11716
rect 15470 11704 15476 11716
rect 15528 11704 15534 11756
rect 8921 11679 8979 11685
rect 8921 11676 8933 11679
rect 8772 11648 8933 11676
rect 8665 11639 8723 11645
rect 8921 11645 8933 11648
rect 8967 11645 8979 11679
rect 10870 11676 10876 11688
rect 8921 11639 8979 11645
rect 9048 11648 10732 11676
rect 10783 11648 10876 11676
rect 7650 11568 7656 11620
rect 7708 11608 7714 11620
rect 7708 11580 8432 11608
rect 7708 11568 7714 11580
rect 8202 11540 8208 11552
rect 7156 11512 7328 11540
rect 8163 11512 8208 11540
rect 7156 11500 7162 11512
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8404 11540 8432 11580
rect 8478 11568 8484 11620
rect 8536 11608 8542 11620
rect 9048 11608 9076 11648
rect 8536 11580 9076 11608
rect 8536 11568 8542 11580
rect 9858 11568 9864 11620
rect 9916 11608 9922 11620
rect 10704 11608 10732 11648
rect 10870 11636 10876 11648
rect 10928 11676 10934 11688
rect 12434 11676 12440 11688
rect 10928 11648 12440 11676
rect 10928 11636 10934 11648
rect 12434 11636 12440 11648
rect 12492 11636 12498 11688
rect 12805 11679 12863 11685
rect 12805 11645 12817 11679
rect 12851 11676 12863 11679
rect 12851 11648 13032 11676
rect 12851 11645 12863 11648
rect 12805 11639 12863 11645
rect 13004 11620 13032 11648
rect 14458 11636 14464 11688
rect 14516 11676 14522 11688
rect 14829 11679 14887 11685
rect 14829 11676 14841 11679
rect 14516 11648 14841 11676
rect 14516 11636 14522 11648
rect 14829 11645 14841 11648
rect 14875 11676 14887 11679
rect 16390 11676 16396 11688
rect 14875 11648 16396 11676
rect 14875 11645 14887 11648
rect 14829 11639 14887 11645
rect 16390 11636 16396 11648
rect 16448 11636 16454 11688
rect 10778 11608 10784 11620
rect 9916 11580 10548 11608
rect 10704 11580 10784 11608
rect 9916 11568 9922 11580
rect 10520 11549 10548 11580
rect 10778 11568 10784 11580
rect 10836 11568 10842 11620
rect 11422 11568 11428 11620
rect 11480 11568 11486 11620
rect 11701 11611 11759 11617
rect 11701 11577 11713 11611
rect 11747 11608 11759 11611
rect 12618 11608 12624 11620
rect 11747 11580 12624 11608
rect 11747 11577 11759 11580
rect 11701 11571 11759 11577
rect 12618 11568 12624 11580
rect 12676 11568 12682 11620
rect 12710 11568 12716 11620
rect 12768 11608 12774 11620
rect 12897 11611 12955 11617
rect 12897 11608 12909 11611
rect 12768 11580 12909 11608
rect 12768 11568 12774 11580
rect 12897 11577 12909 11580
rect 12943 11577 12955 11611
rect 12897 11571 12955 11577
rect 12986 11568 12992 11620
rect 13044 11568 13050 11620
rect 14001 11611 14059 11617
rect 14001 11577 14013 11611
rect 14047 11608 14059 11611
rect 14734 11608 14740 11620
rect 14047 11580 14740 11608
rect 14047 11577 14059 11580
rect 14001 11571 14059 11577
rect 14734 11568 14740 11580
rect 14792 11568 14798 11620
rect 10045 11543 10103 11549
rect 10045 11540 10057 11543
rect 8404 11512 10057 11540
rect 10045 11509 10057 11512
rect 10091 11509 10103 11543
rect 10045 11503 10103 11509
rect 10505 11543 10563 11549
rect 10505 11509 10517 11543
rect 10551 11509 10563 11543
rect 10505 11503 10563 11509
rect 10965 11543 11023 11549
rect 10965 11509 10977 11543
rect 11011 11540 11023 11543
rect 11440 11540 11468 11568
rect 13446 11540 13452 11552
rect 11011 11512 13452 11540
rect 11011 11509 11023 11512
rect 10965 11503 11023 11509
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 13630 11540 13636 11552
rect 13591 11512 13636 11540
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 14090 11500 14096 11552
rect 14148 11540 14154 11552
rect 15010 11540 15016 11552
rect 14148 11512 14193 11540
rect 14971 11512 15016 11540
rect 14148 11500 14154 11512
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 1104 11450 15824 11472
rect 1104 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 6104 11450
rect 6156 11398 10843 11450
rect 10895 11398 10907 11450
rect 10959 11398 10971 11450
rect 11023 11398 11035 11450
rect 11087 11398 15824 11450
rect 1104 11376 15824 11398
rect 11330 11336 11336 11348
rect 1596 11308 11336 11336
rect 1596 11209 1624 11308
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 11514 11336 11520 11348
rect 11475 11308 11520 11336
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 11977 11339 12035 11345
rect 11977 11336 11989 11339
rect 11756 11308 11989 11336
rect 11756 11296 11762 11308
rect 11977 11305 11989 11308
rect 12023 11305 12035 11339
rect 11977 11299 12035 11305
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 12713 11339 12771 11345
rect 12713 11336 12725 11339
rect 12584 11308 12725 11336
rect 12584 11296 12590 11308
rect 12713 11305 12725 11308
rect 12759 11305 12771 11339
rect 12713 11299 12771 11305
rect 12802 11296 12808 11348
rect 12860 11336 12866 11348
rect 12986 11336 12992 11348
rect 12860 11308 12992 11336
rect 12860 11296 12866 11308
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 13909 11339 13967 11345
rect 13909 11305 13921 11339
rect 13955 11336 13967 11339
rect 14090 11336 14096 11348
rect 13955 11308 14096 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 1854 11268 1860 11280
rect 1815 11240 1860 11268
rect 1854 11228 1860 11240
rect 1912 11228 1918 11280
rect 2774 11268 2780 11280
rect 2148 11240 2780 11268
rect 2148 11209 2176 11240
rect 2774 11228 2780 11240
rect 2832 11268 2838 11280
rect 4890 11268 4896 11280
rect 2832 11240 4108 11268
rect 2832 11228 2838 11240
rect 4080 11209 4108 11240
rect 4172 11240 4896 11268
rect 1581 11203 1639 11209
rect 1581 11169 1593 11203
rect 1627 11169 1639 11203
rect 1581 11163 1639 11169
rect 2133 11203 2191 11209
rect 2133 11169 2145 11203
rect 2179 11169 2191 11203
rect 2133 11163 2191 11169
rect 2400 11203 2458 11209
rect 2400 11169 2412 11203
rect 2446 11200 2458 11203
rect 4065 11203 4123 11209
rect 2446 11172 4016 11200
rect 2446 11169 2458 11172
rect 2400 11163 2458 11169
rect 3988 11132 4016 11172
rect 4065 11169 4077 11203
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 4172 11132 4200 11240
rect 4890 11228 4896 11240
rect 4948 11228 4954 11280
rect 6273 11271 6331 11277
rect 6273 11237 6285 11271
rect 6319 11268 6331 11271
rect 7184 11271 7242 11277
rect 6319 11240 7144 11268
rect 6319 11237 6331 11240
rect 6273 11231 6331 11237
rect 4332 11203 4390 11209
rect 4332 11169 4344 11203
rect 4378 11200 4390 11203
rect 4706 11200 4712 11212
rect 4378 11172 4712 11200
rect 4378 11169 4390 11172
rect 4332 11163 4390 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11200 6147 11203
rect 6546 11200 6552 11212
rect 6135 11172 6552 11200
rect 6135 11169 6147 11172
rect 6089 11163 6147 11169
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 7116 11200 7144 11240
rect 7184 11237 7196 11271
rect 7230 11268 7242 11271
rect 7374 11268 7380 11280
rect 7230 11240 7380 11268
rect 7230 11237 7242 11240
rect 7184 11231 7242 11237
rect 7374 11228 7380 11240
rect 7432 11228 7438 11280
rect 8202 11228 8208 11280
rect 8260 11268 8266 11280
rect 9398 11268 9404 11280
rect 8260 11240 9404 11268
rect 8260 11228 8266 11240
rect 9398 11228 9404 11240
rect 9456 11268 9462 11280
rect 9922 11271 9980 11277
rect 9922 11268 9934 11271
rect 9456 11240 9934 11268
rect 9456 11228 9462 11240
rect 9922 11237 9934 11240
rect 9968 11237 9980 11271
rect 9922 11231 9980 11237
rect 10502 11228 10508 11280
rect 10560 11268 10566 11280
rect 10778 11268 10784 11280
rect 10560 11240 10784 11268
rect 10560 11228 10566 11240
rect 10778 11228 10784 11240
rect 10836 11228 10842 11280
rect 13170 11228 13176 11280
rect 13228 11268 13234 11280
rect 14369 11271 14427 11277
rect 14369 11268 14381 11271
rect 13228 11240 14381 11268
rect 13228 11228 13234 11240
rect 14369 11237 14381 11240
rect 14415 11237 14427 11271
rect 14369 11231 14427 11237
rect 11514 11200 11520 11212
rect 7116 11172 11520 11200
rect 11514 11160 11520 11172
rect 11572 11160 11578 11212
rect 11885 11203 11943 11209
rect 11885 11169 11897 11203
rect 11931 11169 11943 11203
rect 11885 11163 11943 11169
rect 3988 11104 4200 11132
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6880 11104 6929 11132
rect 6880 11092 6886 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 8754 11132 8760 11144
rect 8715 11104 8760 11132
rect 6917 11095 6975 11101
rect 8754 11092 8760 11104
rect 8812 11092 8818 11144
rect 9674 11132 9680 11144
rect 9635 11104 9680 11132
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 10686 11092 10692 11144
rect 10744 11132 10750 11144
rect 11790 11132 11796 11144
rect 10744 11104 11796 11132
rect 10744 11092 10750 11104
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 3234 11024 3240 11076
rect 3292 11064 3298 11076
rect 3418 11064 3424 11076
rect 3292 11036 3424 11064
rect 3292 11024 3298 11036
rect 3418 11024 3424 11036
rect 3476 11064 3482 11076
rect 3513 11067 3571 11073
rect 3513 11064 3525 11067
rect 3476 11036 3525 11064
rect 3476 11024 3482 11036
rect 3513 11033 3525 11036
rect 3559 11033 3571 11067
rect 3513 11027 3571 11033
rect 3786 11024 3792 11076
rect 3844 11064 3850 11076
rect 4062 11064 4068 11076
rect 3844 11036 4068 11064
rect 3844 11024 3850 11036
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 5074 11024 5080 11076
rect 5132 11064 5138 11076
rect 5445 11067 5503 11073
rect 5445 11064 5457 11067
rect 5132 11036 5457 11064
rect 5132 11024 5138 11036
rect 5445 11033 5457 11036
rect 5491 11033 5503 11067
rect 5445 11027 5503 11033
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 5905 11067 5963 11073
rect 5905 11064 5917 11067
rect 5592 11036 5917 11064
rect 5592 11024 5598 11036
rect 5905 11033 5917 11036
rect 5951 11033 5963 11067
rect 5905 11027 5963 11033
rect 8018 11024 8024 11076
rect 8076 11064 8082 11076
rect 8297 11067 8355 11073
rect 8297 11064 8309 11067
rect 8076 11036 8309 11064
rect 8076 11024 8082 11036
rect 8297 11033 8309 11036
rect 8343 11064 8355 11067
rect 9490 11064 9496 11076
rect 8343 11036 9496 11064
rect 8343 11033 8355 11036
rect 8297 11027 8355 11033
rect 9490 11024 9496 11036
rect 9548 11024 9554 11076
rect 10778 11024 10784 11076
rect 10836 11064 10842 11076
rect 11057 11067 11115 11073
rect 11057 11064 11069 11067
rect 10836 11036 11069 11064
rect 10836 11024 10842 11036
rect 11057 11033 11069 11036
rect 11103 11033 11115 11067
rect 11900 11064 11928 11163
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 13078 11200 13084 11212
rect 12492 11172 13084 11200
rect 12492 11160 12498 11172
rect 13078 11160 13084 11172
rect 13136 11160 13142 11212
rect 13538 11200 13544 11212
rect 13188 11172 13544 11200
rect 12066 11132 12072 11144
rect 12027 11104 12072 11132
rect 12066 11092 12072 11104
rect 12124 11092 12130 11144
rect 13188 11141 13216 11172
rect 13538 11160 13544 11172
rect 13596 11200 13602 11212
rect 14090 11200 14096 11212
rect 13596 11172 14096 11200
rect 13596 11160 13602 11172
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 14274 11200 14280 11212
rect 14235 11172 14280 11200
rect 14274 11160 14280 11172
rect 14332 11160 14338 11212
rect 13173 11135 13231 11141
rect 13173 11101 13185 11135
rect 13219 11101 13231 11135
rect 13173 11095 13231 11101
rect 13262 11092 13268 11144
rect 13320 11132 13326 11144
rect 14553 11135 14611 11141
rect 13320 11104 13365 11132
rect 13320 11092 13326 11104
rect 14553 11101 14565 11135
rect 14599 11132 14611 11135
rect 14642 11132 14648 11144
rect 14599 11104 14648 11132
rect 14599 11101 14611 11104
rect 14553 11095 14611 11101
rect 13998 11064 14004 11076
rect 11900 11036 14004 11064
rect 11057 11027 11115 11033
rect 13998 11024 14004 11036
rect 14056 11024 14062 11076
rect 2498 10956 2504 11008
rect 2556 10996 2562 11008
rect 4246 10996 4252 11008
rect 2556 10968 4252 10996
rect 2556 10956 2562 10968
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 5350 10956 5356 11008
rect 5408 10996 5414 11008
rect 14568 10996 14596 11095
rect 14642 11092 14648 11104
rect 14700 11092 14706 11144
rect 5408 10968 14596 10996
rect 5408 10956 5414 10968
rect 1104 10906 15824 10928
rect 1104 10854 3447 10906
rect 3499 10854 3511 10906
rect 3563 10854 3575 10906
rect 3627 10854 3639 10906
rect 3691 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 13308 10906
rect 13360 10854 13372 10906
rect 13424 10854 13436 10906
rect 13488 10854 13500 10906
rect 13552 10854 15824 10906
rect 1104 10832 15824 10854
rect 1302 10752 1308 10804
rect 1360 10792 1366 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1360 10764 1593 10792
rect 1360 10752 1366 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 1581 10755 1639 10761
rect 1857 10795 1915 10801
rect 1857 10761 1869 10795
rect 1903 10792 1915 10795
rect 2130 10792 2136 10804
rect 1903 10764 2136 10792
rect 1903 10761 1915 10764
rect 1857 10755 1915 10761
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 6270 10792 6276 10804
rect 2280 10764 4200 10792
rect 6231 10764 6276 10792
rect 2280 10752 2286 10764
rect 4172 10736 4200 10764
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 6546 10752 6552 10804
rect 6604 10792 6610 10804
rect 11238 10792 11244 10804
rect 6604 10764 11244 10792
rect 6604 10752 6610 10764
rect 11238 10752 11244 10764
rect 11296 10752 11302 10804
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 12894 10792 12900 10804
rect 11756 10764 12900 10792
rect 11756 10752 11762 10764
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 13630 10792 13636 10804
rect 13591 10764 13636 10792
rect 13630 10752 13636 10764
rect 13688 10752 13694 10804
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14090 10792 14096 10804
rect 13964 10764 14096 10792
rect 13964 10752 13970 10764
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 4154 10684 4160 10736
rect 4212 10684 4218 10736
rect 7926 10684 7932 10736
rect 7984 10724 7990 10736
rect 8205 10727 8263 10733
rect 8205 10724 8217 10727
rect 7984 10696 8217 10724
rect 7984 10684 7990 10696
rect 8205 10693 8217 10696
rect 8251 10693 8263 10727
rect 8205 10687 8263 10693
rect 11790 10684 11796 10736
rect 11848 10724 11854 10736
rect 11885 10727 11943 10733
rect 11885 10724 11897 10727
rect 11848 10696 11897 10724
rect 11848 10684 11854 10696
rect 11885 10693 11897 10696
rect 11931 10693 11943 10727
rect 13446 10724 13452 10736
rect 11885 10687 11943 10693
rect 12820 10696 13452 10724
rect 2498 10656 2504 10668
rect 2459 10628 2504 10656
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 4062 10616 4068 10668
rect 4120 10656 4126 10668
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4120 10628 4905 10656
rect 4120 10616 4126 10628
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 6822 10656 6828 10668
rect 6783 10628 6828 10656
rect 4893 10619 4951 10625
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 10134 10656 10140 10668
rect 9732 10628 10140 10656
rect 9732 10616 9738 10628
rect 10134 10616 10140 10628
rect 10192 10656 10198 10668
rect 10505 10659 10563 10665
rect 10505 10656 10517 10659
rect 10192 10628 10517 10656
rect 10192 10616 10198 10628
rect 10505 10625 10517 10628
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 11572 10628 11836 10656
rect 11572 10616 11578 10628
rect 1394 10588 1400 10600
rect 1355 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10548 1458 10600
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 3053 10591 3111 10597
rect 3053 10588 3065 10591
rect 2832 10560 3065 10588
rect 2832 10548 2838 10560
rect 3053 10557 3065 10560
rect 3099 10557 3111 10591
rect 3053 10551 3111 10557
rect 7092 10591 7150 10597
rect 7092 10557 7104 10591
rect 7138 10588 7150 10591
rect 8018 10588 8024 10600
rect 7138 10560 8024 10588
rect 7138 10557 7150 10560
rect 7092 10551 7150 10557
rect 8018 10548 8024 10560
rect 8076 10548 8082 10600
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 8294 10588 8300 10600
rect 8260 10560 8300 10588
rect 8260 10548 8266 10560
rect 8294 10548 8300 10560
rect 8352 10588 8358 10600
rect 8665 10591 8723 10597
rect 8665 10588 8677 10591
rect 8352 10560 8677 10588
rect 8352 10548 8358 10560
rect 8665 10557 8677 10560
rect 8711 10588 8723 10591
rect 9692 10588 9720 10616
rect 11808 10600 11836 10628
rect 11606 10588 11612 10600
rect 8711 10560 9720 10588
rect 10612 10560 11612 10588
rect 8711 10557 8723 10560
rect 8665 10551 8723 10557
rect 1854 10480 1860 10532
rect 1912 10520 1918 10532
rect 2317 10523 2375 10529
rect 2317 10520 2329 10523
rect 1912 10492 2329 10520
rect 1912 10480 1918 10492
rect 2317 10489 2329 10492
rect 2363 10489 2375 10523
rect 2317 10483 2375 10489
rect 3320 10523 3378 10529
rect 3320 10489 3332 10523
rect 3366 10520 3378 10523
rect 3366 10492 3556 10520
rect 3366 10489 3378 10492
rect 3320 10483 3378 10489
rect 2222 10452 2228 10464
rect 2183 10424 2228 10452
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 3528 10452 3556 10492
rect 5074 10480 5080 10532
rect 5132 10529 5138 10532
rect 5132 10523 5196 10529
rect 5132 10489 5150 10523
rect 5184 10489 5196 10523
rect 8910 10523 8968 10529
rect 8910 10520 8922 10523
rect 5132 10483 5196 10489
rect 5368 10492 8922 10520
rect 5132 10480 5138 10483
rect 4338 10452 4344 10464
rect 3528 10424 4344 10452
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 4982 10452 4988 10464
rect 4479 10424 4988 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 4982 10412 4988 10424
rect 5040 10452 5046 10464
rect 5368 10452 5396 10492
rect 8910 10489 8922 10492
rect 8956 10489 8968 10523
rect 10612 10520 10640 10560
rect 11606 10548 11612 10560
rect 11664 10548 11670 10600
rect 11790 10548 11796 10600
rect 11848 10548 11854 10600
rect 12820 10597 12848 10696
rect 13446 10684 13452 10696
rect 13504 10724 13510 10736
rect 14918 10724 14924 10736
rect 13504 10696 14924 10724
rect 13504 10684 13510 10696
rect 14918 10684 14924 10696
rect 14976 10684 14982 10736
rect 12986 10656 12992 10668
rect 12947 10628 12992 10656
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13170 10616 13176 10668
rect 13228 10656 13234 10668
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 13228 10628 14197 10656
rect 13228 10616 13234 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 12805 10591 12863 10597
rect 12805 10557 12817 10591
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10588 12955 10591
rect 14090 10588 14096 10600
rect 12943 10560 14096 10588
rect 12943 10557 12955 10560
rect 12897 10551 12955 10557
rect 14090 10548 14096 10560
rect 14148 10588 14154 10600
rect 14366 10588 14372 10600
rect 14148 10560 14372 10588
rect 14148 10548 14154 10560
rect 14366 10548 14372 10560
rect 14424 10548 14430 10600
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 14829 10591 14887 10597
rect 14829 10588 14841 10591
rect 14608 10560 14841 10588
rect 14608 10548 14614 10560
rect 14829 10557 14841 10560
rect 14875 10557 14887 10591
rect 14829 10551 14887 10557
rect 8910 10483 8968 10489
rect 9048 10492 10640 10520
rect 10772 10523 10830 10529
rect 5040 10424 5396 10452
rect 5040 10412 5046 10424
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 9048 10452 9076 10492
rect 10772 10489 10784 10523
rect 10818 10520 10830 10523
rect 11146 10520 11152 10532
rect 10818 10492 11152 10520
rect 10818 10489 10830 10492
rect 10772 10483 10830 10489
rect 11146 10480 11152 10492
rect 11204 10520 11210 10532
rect 13262 10520 13268 10532
rect 11204 10492 13268 10520
rect 11204 10480 11210 10492
rect 13262 10480 13268 10492
rect 13320 10480 13326 10532
rect 13906 10480 13912 10532
rect 13964 10520 13970 10532
rect 13964 10492 14136 10520
rect 13964 10480 13970 10492
rect 10042 10452 10048 10464
rect 5500 10424 9076 10452
rect 9955 10424 10048 10452
rect 5500 10412 5506 10424
rect 10042 10412 10048 10424
rect 10100 10452 10106 10464
rect 11514 10452 11520 10464
rect 10100 10424 11520 10452
rect 10100 10412 10106 10424
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12492 10424 12537 10452
rect 12492 10412 12498 10424
rect 12894 10412 12900 10464
rect 12952 10452 12958 10464
rect 13078 10452 13084 10464
rect 12952 10424 13084 10452
rect 12952 10412 12958 10424
rect 13078 10412 13084 10424
rect 13136 10452 13142 10464
rect 14108 10461 14136 10492
rect 14001 10455 14059 10461
rect 14001 10452 14013 10455
rect 13136 10424 14013 10452
rect 13136 10412 13142 10424
rect 14001 10421 14013 10424
rect 14047 10421 14059 10455
rect 14001 10415 14059 10421
rect 14093 10455 14151 10461
rect 14093 10421 14105 10455
rect 14139 10421 14151 10455
rect 15010 10452 15016 10464
rect 14971 10424 15016 10452
rect 14093 10415 14151 10421
rect 15010 10412 15016 10424
rect 15068 10412 15074 10464
rect 1104 10362 15824 10384
rect 1104 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 6104 10362
rect 6156 10310 10843 10362
rect 10895 10310 10907 10362
rect 10959 10310 10971 10362
rect 11023 10310 11035 10362
rect 11087 10310 15824 10362
rect 1104 10288 15824 10310
rect 4614 10248 4620 10260
rect 1412 10220 2544 10248
rect 1412 10121 1440 10220
rect 2406 10189 2412 10192
rect 2400 10180 2412 10189
rect 2367 10152 2412 10180
rect 2400 10143 2412 10152
rect 2406 10140 2412 10143
rect 2464 10140 2470 10192
rect 2516 10180 2544 10220
rect 4356 10220 4620 10248
rect 4356 10180 4384 10220
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 5810 10248 5816 10260
rect 5543 10220 5816 10248
rect 2516 10152 4384 10180
rect 4430 10140 4436 10192
rect 4488 10180 4494 10192
rect 5442 10180 5448 10192
rect 4488 10152 5448 10180
rect 4488 10140 4494 10152
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10081 1455 10115
rect 1397 10075 1455 10081
rect 2133 10115 2191 10121
rect 2133 10081 2145 10115
rect 2179 10112 2191 10115
rect 2774 10112 2780 10124
rect 2179 10084 2780 10112
rect 2179 10081 2191 10084
rect 2133 10075 2191 10081
rect 2774 10072 2780 10084
rect 2832 10112 2838 10124
rect 4062 10112 4068 10124
rect 2832 10084 4068 10112
rect 2832 10072 2838 10084
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 4332 10115 4390 10121
rect 4332 10081 4344 10115
rect 4378 10112 4390 10115
rect 5543 10112 5571 10220
rect 5810 10208 5816 10220
rect 5868 10248 5874 10260
rect 6546 10248 6552 10260
rect 5868 10220 6552 10248
rect 5868 10208 5874 10220
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 7285 10251 7343 10257
rect 7285 10217 7297 10251
rect 7331 10248 7343 10251
rect 7374 10248 7380 10260
rect 7331 10220 7380 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 7374 10208 7380 10220
rect 7432 10248 7438 10260
rect 7742 10248 7748 10260
rect 7432 10220 7748 10248
rect 7432 10208 7438 10220
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 8846 10248 8852 10260
rect 8260 10220 8852 10248
rect 8260 10208 8266 10220
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 9122 10248 9128 10260
rect 9083 10220 9128 10248
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9306 10208 9312 10260
rect 9364 10248 9370 10260
rect 9490 10248 9496 10260
rect 9364 10220 9496 10248
rect 9364 10208 9370 10220
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 10502 10208 10508 10260
rect 10560 10248 10566 10260
rect 11606 10248 11612 10260
rect 10560 10220 11612 10248
rect 10560 10208 10566 10220
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 11885 10251 11943 10257
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 12158 10248 12164 10260
rect 11931 10220 12164 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 13173 10251 13231 10257
rect 13173 10248 13185 10251
rect 12492 10220 13185 10248
rect 12492 10208 12498 10220
rect 13173 10217 13185 10220
rect 13219 10217 13231 10251
rect 13173 10211 13231 10217
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 13872 10220 13921 10248
rect 13872 10208 13878 10220
rect 13909 10217 13921 10220
rect 13955 10217 13967 10251
rect 13909 10211 13967 10217
rect 6172 10183 6230 10189
rect 6172 10149 6184 10183
rect 6218 10180 6230 10183
rect 6270 10180 6276 10192
rect 6218 10152 6276 10180
rect 6218 10149 6230 10152
rect 6172 10143 6230 10149
rect 6270 10140 6276 10152
rect 6328 10140 6334 10192
rect 7834 10140 7840 10192
rect 7892 10180 7898 10192
rect 7990 10183 8048 10189
rect 7990 10180 8002 10183
rect 7892 10152 8002 10180
rect 7892 10140 7898 10152
rect 7990 10149 8002 10152
rect 8036 10149 8048 10183
rect 7990 10143 8048 10149
rect 8110 10140 8116 10192
rect 8168 10180 8174 10192
rect 14277 10183 14335 10189
rect 14277 10180 14289 10183
rect 8168 10152 12480 10180
rect 8168 10140 8174 10152
rect 12452 10124 12480 10152
rect 12544 10152 14289 10180
rect 7745 10115 7803 10121
rect 7745 10112 7757 10115
rect 4378 10084 5571 10112
rect 5920 10084 7757 10112
rect 4378 10081 4390 10084
rect 4332 10075 4390 10081
rect 5258 10004 5264 10056
rect 5316 10044 5322 10056
rect 5920 10053 5948 10084
rect 7745 10081 7757 10084
rect 7791 10112 7803 10115
rect 8294 10112 8300 10124
rect 7791 10084 8300 10112
rect 7791 10081 7803 10084
rect 7745 10075 7803 10081
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 9933 10115 9991 10121
rect 9933 10112 9945 10115
rect 8772 10084 9945 10112
rect 5905 10047 5963 10053
rect 5905 10044 5917 10047
rect 5316 10016 5917 10044
rect 5316 10004 5322 10016
rect 5905 10013 5917 10016
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 3418 9936 3424 9988
rect 3476 9936 3482 9988
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 5445 9979 5503 9985
rect 5445 9976 5457 9979
rect 5408 9948 5457 9976
rect 5408 9936 5414 9948
rect 5445 9945 5457 9948
rect 5491 9945 5503 9979
rect 5445 9939 5503 9945
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 3436 9908 3464 9936
rect 1627 9880 3464 9908
rect 3513 9911 3571 9917
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 3513 9877 3525 9911
rect 3559 9908 3571 9911
rect 4246 9908 4252 9920
rect 3559 9880 4252 9908
rect 3559 9877 3571 9880
rect 3513 9871 3571 9877
rect 4246 9868 4252 9880
rect 4304 9908 4310 9920
rect 8772 9908 8800 10084
rect 9933 10081 9945 10084
rect 9979 10081 9991 10115
rect 9933 10075 9991 10081
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 10560 10084 11284 10112
rect 10560 10072 10566 10084
rect 8846 10004 8852 10056
rect 8904 10044 8910 10056
rect 9306 10044 9312 10056
rect 8904 10016 9312 10044
rect 8904 10004 8910 10016
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 10778 9936 10784 9988
rect 10836 9976 10842 9988
rect 11057 9979 11115 9985
rect 11057 9976 11069 9979
rect 10836 9948 11069 9976
rect 10836 9936 10842 9948
rect 11057 9945 11069 9948
rect 11103 9976 11115 9979
rect 11146 9976 11152 9988
rect 11103 9948 11152 9976
rect 11103 9945 11115 9948
rect 11057 9939 11115 9945
rect 11146 9936 11152 9948
rect 11204 9936 11210 9988
rect 11256 9976 11284 10084
rect 11514 10072 11520 10124
rect 11572 10112 11578 10124
rect 11572 10084 12112 10112
rect 11572 10072 11578 10084
rect 11698 10004 11704 10056
rect 11756 10044 11762 10056
rect 12084 10053 12112 10084
rect 12434 10072 12440 10124
rect 12492 10072 12498 10124
rect 11977 10047 12035 10053
rect 11977 10044 11989 10047
rect 11756 10016 11989 10044
rect 11756 10004 11762 10016
rect 11977 10013 11989 10016
rect 12023 10013 12035 10047
rect 11977 10007 12035 10013
rect 12069 10047 12127 10053
rect 12069 10013 12081 10047
rect 12115 10013 12127 10047
rect 12544 10044 12572 10152
rect 14277 10149 14289 10152
rect 14323 10149 14335 10183
rect 14277 10143 14335 10149
rect 13078 10112 13084 10124
rect 13039 10084 13084 10112
rect 13078 10072 13084 10084
rect 13136 10072 13142 10124
rect 13630 10072 13636 10124
rect 13688 10072 13694 10124
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 13872 10084 14504 10112
rect 13872 10072 13878 10084
rect 12069 10007 12127 10013
rect 12176 10016 12572 10044
rect 13265 10047 13323 10053
rect 12176 9976 12204 10016
rect 13265 10013 13277 10047
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 11256 9948 12204 9976
rect 12434 9936 12440 9988
rect 12492 9976 12498 9988
rect 12713 9979 12771 9985
rect 12713 9976 12725 9979
rect 12492 9948 12725 9976
rect 12492 9936 12498 9948
rect 12713 9945 12725 9948
rect 12759 9945 12771 9979
rect 12713 9939 12771 9945
rect 4304 9880 8800 9908
rect 4304 9868 4310 9880
rect 8846 9868 8852 9920
rect 8904 9908 8910 9920
rect 9030 9908 9036 9920
rect 8904 9880 9036 9908
rect 8904 9868 8910 9880
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 9214 9868 9220 9920
rect 9272 9908 9278 9920
rect 11517 9911 11575 9917
rect 11517 9908 11529 9911
rect 9272 9880 11529 9908
rect 9272 9868 9278 9880
rect 11517 9877 11529 9880
rect 11563 9877 11575 9911
rect 11517 9871 11575 9877
rect 12158 9868 12164 9920
rect 12216 9908 12222 9920
rect 13280 9908 13308 10007
rect 12216 9880 13308 9908
rect 13648 9908 13676 10072
rect 14476 10056 14504 10084
rect 14366 10044 14372 10056
rect 14327 10016 14372 10044
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 14458 10004 14464 10056
rect 14516 10044 14522 10056
rect 14516 10016 14609 10044
rect 14516 10004 14522 10016
rect 13906 9908 13912 9920
rect 13648 9880 13912 9908
rect 12216 9868 12222 9880
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 1104 9818 15824 9840
rect 1104 9766 3447 9818
rect 3499 9766 3511 9818
rect 3563 9766 3575 9818
rect 3627 9766 3639 9818
rect 3691 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 13308 9818
rect 13360 9766 13372 9818
rect 13424 9766 13436 9818
rect 13488 9766 13500 9818
rect 13552 9766 15824 9818
rect 1104 9744 15824 9766
rect 1854 9704 1860 9716
rect 1815 9676 1860 9704
rect 1854 9664 1860 9676
rect 1912 9664 1918 9716
rect 4430 9704 4436 9716
rect 2976 9676 4016 9704
rect 4391 9676 4436 9704
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2976 9568 3004 9676
rect 3988 9636 4016 9676
rect 4430 9664 4436 9676
rect 4488 9664 4494 9716
rect 5276 9676 6224 9704
rect 3988 9608 4108 9636
rect 2547 9540 3004 9568
rect 4080 9568 4108 9608
rect 4154 9596 4160 9648
rect 4212 9636 4218 9648
rect 4985 9639 5043 9645
rect 4985 9636 4997 9639
rect 4212 9608 4997 9636
rect 4212 9596 4218 9608
rect 4985 9605 4997 9608
rect 5031 9636 5043 9639
rect 5276 9636 5304 9676
rect 5031 9608 5304 9636
rect 6196 9636 6224 9676
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 10042 9704 10048 9716
rect 6604 9676 10048 9704
rect 6604 9664 6610 9676
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 11146 9664 11152 9716
rect 11204 9704 11210 9716
rect 11606 9704 11612 9716
rect 11204 9676 11612 9704
rect 11204 9664 11210 9676
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 11882 9664 11888 9716
rect 11940 9704 11946 9716
rect 12158 9704 12164 9716
rect 11940 9676 12164 9704
rect 11940 9664 11946 9676
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12437 9707 12495 9713
rect 12437 9673 12449 9707
rect 12483 9704 12495 9707
rect 13078 9704 13084 9716
rect 12483 9676 13084 9704
rect 12483 9673 12495 9676
rect 12437 9667 12495 9673
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 15013 9707 15071 9713
rect 15013 9704 15025 9707
rect 13188 9676 15025 9704
rect 7282 9636 7288 9648
rect 6196 9608 7288 9636
rect 5031 9605 5043 9608
rect 4985 9599 5043 9605
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 8018 9596 8024 9648
rect 8076 9636 8082 9648
rect 9030 9636 9036 9648
rect 8076 9608 9036 9636
rect 8076 9596 8082 9608
rect 9030 9596 9036 9608
rect 9088 9596 9094 9648
rect 10413 9639 10471 9645
rect 10413 9605 10425 9639
rect 10459 9605 10471 9639
rect 13188 9636 13216 9676
rect 15013 9673 15025 9676
rect 15059 9673 15071 9707
rect 15013 9667 15071 9673
rect 10413 9599 10471 9605
rect 11716 9608 13216 9636
rect 5074 9568 5080 9580
rect 4080 9540 5080 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 5258 9568 5264 9580
rect 5219 9540 5264 9568
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 7098 9568 7104 9580
rect 6328 9540 7104 9568
rect 6328 9528 6334 9540
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7742 9528 7748 9580
rect 7800 9568 7806 9580
rect 7800 9540 9168 9568
rect 7800 9528 7806 9540
rect 2130 9460 2136 9512
rect 2188 9500 2194 9512
rect 2866 9500 2872 9512
rect 2188 9472 2872 9500
rect 2188 9460 2194 9472
rect 2866 9460 2872 9472
rect 2924 9500 2930 9512
rect 3053 9503 3111 9509
rect 3053 9500 3065 9503
rect 2924 9472 3065 9500
rect 2924 9460 2930 9472
rect 3053 9469 3065 9472
rect 3099 9469 3111 9503
rect 3053 9463 3111 9469
rect 5169 9503 5227 9509
rect 5169 9469 5181 9503
rect 5215 9500 5227 9503
rect 6730 9500 6736 9512
rect 5215 9472 6736 9500
rect 5215 9469 5227 9472
rect 5169 9463 5227 9469
rect 6730 9460 6736 9472
rect 6788 9500 6794 9512
rect 8757 9503 8815 9509
rect 8757 9500 8769 9503
rect 6788 9472 8769 9500
rect 6788 9460 6794 9472
rect 8757 9469 8769 9472
rect 8803 9469 8815 9503
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 8757 9463 8815 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9140 9500 9168 9540
rect 10042 9528 10048 9580
rect 10100 9568 10106 9580
rect 10428 9568 10456 9599
rect 10100 9540 10640 9568
rect 10100 9528 10106 9540
rect 9582 9500 9588 9512
rect 9140 9472 9588 9500
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 9732 9472 10517 9500
rect 9732 9460 9738 9472
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 10612 9500 10640 9540
rect 11606 9500 11612 9512
rect 10612 9472 11612 9500
rect 10505 9463 10563 9469
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 2225 9435 2283 9441
rect 2225 9401 2237 9435
rect 2271 9432 2283 9435
rect 2682 9432 2688 9444
rect 2271 9404 2688 9432
rect 2271 9401 2283 9404
rect 2225 9395 2283 9401
rect 2682 9392 2688 9404
rect 2740 9392 2746 9444
rect 3320 9435 3378 9441
rect 3320 9401 3332 9435
rect 3366 9432 3378 9435
rect 4982 9432 4988 9444
rect 3366 9404 4988 9432
rect 3366 9401 3378 9404
rect 3320 9395 3378 9401
rect 4982 9392 4988 9404
rect 5040 9392 5046 9444
rect 5528 9435 5586 9441
rect 5528 9401 5540 9435
rect 5574 9432 5586 9435
rect 6822 9432 6828 9444
rect 5574 9404 6828 9432
rect 5574 9401 5586 9404
rect 5528 9395 5586 9401
rect 6822 9392 6828 9404
rect 6880 9392 6886 9444
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 7193 9435 7251 9441
rect 7193 9432 7205 9435
rect 7064 9404 7205 9432
rect 7064 9392 7070 9404
rect 7193 9401 7205 9404
rect 7239 9401 7251 9435
rect 7193 9395 7251 9401
rect 7282 9392 7288 9444
rect 7340 9432 7346 9444
rect 8386 9432 8392 9444
rect 7340 9404 8392 9432
rect 7340 9392 7346 9404
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 9300 9435 9358 9441
rect 9300 9401 9312 9435
rect 9346 9432 9358 9435
rect 9398 9432 9404 9444
rect 9346 9404 9404 9432
rect 9346 9401 9358 9404
rect 9300 9395 9358 9401
rect 9398 9392 9404 9404
rect 9456 9392 9462 9444
rect 10594 9392 10600 9444
rect 10652 9432 10658 9444
rect 10772 9435 10830 9441
rect 10772 9432 10784 9435
rect 10652 9404 10784 9432
rect 10652 9392 10658 9404
rect 10772 9401 10784 9404
rect 10818 9432 10830 9435
rect 11514 9432 11520 9444
rect 10818 9404 11520 9432
rect 10818 9401 10830 9404
rect 10772 9395 10830 9401
rect 11514 9392 11520 9404
rect 11572 9392 11578 9444
rect 2314 9324 2320 9376
rect 2372 9364 2378 9376
rect 2372 9336 2417 9364
rect 2372 9324 2378 9336
rect 2590 9324 2596 9376
rect 2648 9364 2654 9376
rect 6638 9364 6644 9376
rect 2648 9336 6644 9364
rect 2648 9324 2654 9336
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 9674 9364 9680 9376
rect 6972 9336 9680 9364
rect 6972 9324 6978 9336
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 11716 9364 11744 9608
rect 13630 9596 13636 9648
rect 13688 9636 13694 9648
rect 15378 9636 15384 9648
rect 13688 9608 15384 9636
rect 13688 9596 13694 9608
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 12986 9568 12992 9580
rect 11900 9540 12992 9568
rect 11900 9376 11928 9540
rect 12986 9528 12992 9540
rect 13044 9568 13050 9580
rect 13081 9571 13139 9577
rect 13081 9568 13093 9571
rect 13044 9540 13093 9568
rect 13044 9528 13050 9540
rect 13081 9537 13093 9540
rect 13127 9568 13139 9571
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 13127 9540 14197 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 12618 9460 12624 9512
rect 12676 9500 12682 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12676 9472 12817 9500
rect 12676 9460 12682 9472
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 12805 9463 12863 9469
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 13262 9500 13268 9512
rect 12943 9472 13268 9500
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 13998 9460 14004 9512
rect 14056 9500 14062 9512
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 14056 9472 14841 9500
rect 14056 9460 14062 9472
rect 14829 9469 14841 9472
rect 14875 9500 14887 9503
rect 14918 9500 14924 9512
rect 14875 9472 14924 9500
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 12434 9392 12440 9444
rect 12492 9432 12498 9444
rect 14093 9435 14151 9441
rect 14093 9432 14105 9435
rect 12492 9404 14105 9432
rect 12492 9392 12498 9404
rect 14093 9401 14105 9404
rect 14139 9401 14151 9435
rect 14093 9395 14151 9401
rect 11882 9364 11888 9376
rect 10008 9336 11744 9364
rect 11843 9336 11888 9364
rect 10008 9324 10014 9336
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 11974 9324 11980 9376
rect 12032 9364 12038 9376
rect 12986 9364 12992 9376
rect 12032 9336 12992 9364
rect 12032 9324 12038 9336
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 13630 9364 13636 9376
rect 13591 9336 13636 9364
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 13998 9364 14004 9376
rect 13959 9336 14004 9364
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 1104 9274 15824 9296
rect 1104 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 6104 9274
rect 6156 9222 10843 9274
rect 10895 9222 10907 9274
rect 10959 9222 10971 9274
rect 11023 9222 11035 9274
rect 11087 9222 15824 9274
rect 1104 9200 15824 9222
rect 2314 9120 2320 9172
rect 2372 9160 2378 9172
rect 9214 9160 9220 9172
rect 2372 9132 9220 9160
rect 2372 9120 2378 9132
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 13817 9163 13875 9169
rect 13817 9160 13829 9163
rect 9640 9132 13829 9160
rect 9640 9120 9646 9132
rect 13817 9129 13829 9132
rect 13863 9129 13875 9163
rect 13817 9123 13875 9129
rect 13998 9120 14004 9172
rect 14056 9160 14062 9172
rect 15102 9160 15108 9172
rect 14056 9132 15108 9160
rect 14056 9120 14062 9132
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 5074 9052 5080 9104
rect 5132 9092 5138 9104
rect 9922 9095 9980 9101
rect 9922 9092 9934 9095
rect 5132 9064 9934 9092
rect 5132 9052 5138 9064
rect 9922 9061 9934 9064
rect 9968 9092 9980 9095
rect 11882 9092 11888 9104
rect 9968 9064 11888 9092
rect 9968 9061 9980 9064
rect 9922 9055 9980 9061
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 13170 9092 13176 9104
rect 11992 9064 13176 9092
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1443 8996 2084 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 1302 8916 1308 8968
rect 1360 8956 1366 8968
rect 1578 8956 1584 8968
rect 1360 8928 1584 8956
rect 1360 8916 1366 8928
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 1210 8780 1216 8832
rect 1268 8820 1274 8832
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 1268 8792 1593 8820
rect 1268 8780 1274 8792
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 2056 8820 2084 8996
rect 2130 8984 2136 9036
rect 2188 9024 2194 9036
rect 2400 9027 2458 9033
rect 2188 8996 2233 9024
rect 2188 8984 2194 8996
rect 2400 8993 2412 9027
rect 2446 9024 2458 9027
rect 4338 9024 4344 9036
rect 2446 8996 4344 9024
rect 2446 8993 2458 8996
rect 2400 8987 2458 8993
rect 4338 8984 4344 8996
rect 4396 8984 4402 9036
rect 4516 9027 4574 9033
rect 4516 8993 4528 9027
rect 4562 9024 4574 9027
rect 5350 9024 5356 9036
rect 4562 8996 5356 9024
rect 4562 8993 4574 8996
rect 4516 8987 4574 8993
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 5721 9027 5779 9033
rect 5721 8993 5733 9027
rect 5767 9024 5779 9027
rect 5810 9024 5816 9036
rect 5767 8996 5816 9024
rect 5767 8993 5779 8996
rect 5721 8987 5779 8993
rect 5810 8984 5816 8996
rect 5868 8984 5874 9036
rect 5988 9027 6046 9033
rect 5988 8993 6000 9027
rect 6034 9024 6046 9027
rect 7006 9024 7012 9036
rect 6034 8996 7012 9024
rect 6034 8993 6046 8996
rect 5988 8987 6046 8993
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 7561 9027 7619 9033
rect 7561 9024 7573 9027
rect 7156 8996 7573 9024
rect 7156 8984 7162 8996
rect 7561 8993 7573 8996
rect 7607 8993 7619 9027
rect 7561 8987 7619 8993
rect 7828 9027 7886 9033
rect 7828 8993 7840 9027
rect 7874 9024 7886 9027
rect 8754 9024 8760 9036
rect 7874 8996 8760 9024
rect 7874 8993 7886 8996
rect 7828 8987 7886 8993
rect 4246 8956 4252 8968
rect 4207 8928 4252 8956
rect 4246 8916 4252 8928
rect 4304 8916 4310 8968
rect 3510 8888 3516 8900
rect 3471 8860 3516 8888
rect 3510 8848 3516 8860
rect 3568 8848 3574 8900
rect 5626 8888 5632 8900
rect 5587 8860 5632 8888
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 6822 8848 6828 8900
rect 6880 8888 6886 8900
rect 7190 8888 7196 8900
rect 6880 8860 7196 8888
rect 6880 8848 6886 8860
rect 7190 8848 7196 8860
rect 7248 8848 7254 8900
rect 4246 8820 4252 8832
rect 2056 8792 4252 8820
rect 1581 8783 1639 8789
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 6914 8820 6920 8832
rect 4488 8792 6920 8820
rect 4488 8780 4494 8792
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 7098 8820 7104 8832
rect 7059 8792 7104 8820
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 7576 8820 7604 8987
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 9398 8984 9404 9036
rect 9456 9024 9462 9036
rect 11773 9027 11831 9033
rect 11773 9024 11785 9027
rect 9456 8996 11785 9024
rect 9456 8984 9462 8996
rect 11773 8993 11785 8996
rect 11819 9024 11831 9027
rect 11992 9024 12020 9064
rect 13170 9052 13176 9064
rect 13228 9052 13234 9104
rect 11819 8996 12020 9024
rect 13725 9027 13783 9033
rect 11819 8993 11831 8996
rect 11773 8987 11831 8993
rect 13725 8993 13737 9027
rect 13771 8993 13783 9027
rect 13725 8987 13783 8993
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 9674 8956 9680 8968
rect 9088 8928 9680 8956
rect 9088 8916 9094 8928
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 11422 8916 11428 8968
rect 11480 8956 11486 8968
rect 11517 8959 11575 8965
rect 11517 8956 11529 8959
rect 11480 8928 11529 8956
rect 11480 8916 11486 8928
rect 11517 8925 11529 8928
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 12710 8956 12716 8968
rect 12584 8928 12716 8956
rect 12584 8916 12590 8928
rect 12710 8916 12716 8928
rect 12768 8916 12774 8968
rect 13170 8916 13176 8968
rect 13228 8956 13234 8968
rect 13740 8956 13768 8987
rect 13228 8928 13768 8956
rect 13228 8916 13234 8928
rect 13814 8916 13820 8968
rect 13872 8956 13878 8968
rect 13909 8959 13967 8965
rect 13909 8956 13921 8959
rect 13872 8928 13921 8956
rect 13872 8916 13878 8928
rect 13909 8925 13921 8928
rect 13955 8925 13967 8959
rect 14550 8956 14556 8968
rect 14511 8928 14556 8956
rect 13909 8919 13967 8925
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 8570 8848 8576 8900
rect 8628 8888 8634 8900
rect 8941 8891 8999 8897
rect 8941 8888 8953 8891
rect 8628 8860 8953 8888
rect 8628 8848 8634 8860
rect 8941 8857 8953 8860
rect 8987 8857 8999 8891
rect 8941 8851 8999 8857
rect 9214 8848 9220 8900
rect 9272 8888 9278 8900
rect 9490 8888 9496 8900
rect 9272 8860 9496 8888
rect 9272 8848 9278 8860
rect 9490 8848 9496 8860
rect 9548 8848 9554 8900
rect 13078 8888 13084 8900
rect 12636 8860 13084 8888
rect 7926 8820 7932 8832
rect 7576 8792 7932 8820
rect 7926 8780 7932 8792
rect 7984 8820 7990 8832
rect 8662 8820 8668 8832
rect 7984 8792 8668 8820
rect 7984 8780 7990 8792
rect 8662 8780 8668 8792
rect 8720 8820 8726 8832
rect 9030 8820 9036 8832
rect 8720 8792 9036 8820
rect 8720 8780 8726 8792
rect 9030 8780 9036 8792
rect 9088 8780 9094 8832
rect 9122 8780 9128 8832
rect 9180 8820 9186 8832
rect 9950 8820 9956 8832
rect 9180 8792 9956 8820
rect 9180 8780 9186 8792
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 11057 8823 11115 8829
rect 11057 8789 11069 8823
rect 11103 8820 11115 8823
rect 11238 8820 11244 8832
rect 11103 8792 11244 8820
rect 11103 8789 11115 8792
rect 11057 8783 11115 8789
rect 11238 8780 11244 8792
rect 11296 8780 11302 8832
rect 11330 8780 11336 8832
rect 11388 8820 11394 8832
rect 12636 8820 12664 8860
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 13354 8888 13360 8900
rect 13315 8860 13360 8888
rect 13354 8848 13360 8860
rect 13412 8848 13418 8900
rect 11388 8792 12664 8820
rect 12897 8823 12955 8829
rect 11388 8780 11394 8792
rect 12897 8789 12909 8823
rect 12943 8820 12955 8823
rect 14182 8820 14188 8832
rect 12943 8792 14188 8820
rect 12943 8789 12955 8792
rect 12897 8783 12955 8789
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 1104 8730 15824 8752
rect 1104 8678 3447 8730
rect 3499 8678 3511 8730
rect 3563 8678 3575 8730
rect 3627 8678 3639 8730
rect 3691 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 13308 8730
rect 13360 8678 13372 8730
rect 13424 8678 13436 8730
rect 13488 8678 13500 8730
rect 13552 8678 15824 8730
rect 1104 8656 15824 8678
rect 2056 8588 4292 8616
rect 2056 8489 2084 8588
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8480 2283 8483
rect 2590 8480 2596 8492
rect 2271 8452 2596 8480
rect 2271 8449 2283 8452
rect 2225 8443 2283 8449
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 2866 8440 2872 8492
rect 2924 8480 2930 8492
rect 3053 8483 3111 8489
rect 3053 8480 3065 8483
rect 2924 8452 3065 8480
rect 2924 8440 2930 8452
rect 3053 8449 3065 8452
rect 3099 8449 3111 8483
rect 4264 8480 4292 8588
rect 4338 8576 4344 8628
rect 4396 8616 4402 8628
rect 4396 8588 7788 8616
rect 4396 8576 4402 8588
rect 4430 8548 4436 8560
rect 4391 8520 4436 8548
rect 4430 8508 4436 8520
rect 4488 8508 4494 8560
rect 6273 8551 6331 8557
rect 6273 8517 6285 8551
rect 6319 8548 6331 8551
rect 7760 8548 7788 8588
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 8205 8619 8263 8625
rect 8205 8616 8217 8619
rect 7892 8588 8217 8616
rect 7892 8576 7898 8588
rect 8205 8585 8217 8588
rect 8251 8585 8263 8619
rect 11882 8616 11888 8628
rect 8205 8579 8263 8585
rect 8687 8588 11888 8616
rect 8687 8548 8715 8588
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 13630 8616 13636 8628
rect 12492 8588 12537 8616
rect 13591 8588 13636 8616
rect 12492 8576 12498 8588
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 10042 8548 10048 8560
rect 6319 8520 6500 8548
rect 7760 8520 8715 8548
rect 10003 8520 10048 8548
rect 6319 8517 6331 8520
rect 6273 8511 6331 8517
rect 4264 8452 5028 8480
rect 3053 8443 3111 8449
rect 1946 8412 1952 8424
rect 1907 8384 1952 8412
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8412 3019 8415
rect 4154 8412 4160 8424
rect 3007 8384 4160 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 4154 8372 4160 8384
rect 4212 8372 4218 8424
rect 4522 8372 4528 8424
rect 4580 8412 4586 8424
rect 4890 8412 4896 8424
rect 4580 8384 4896 8412
rect 4580 8372 4586 8384
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 5000 8412 5028 8452
rect 5994 8440 6000 8492
rect 6052 8480 6058 8492
rect 6362 8480 6368 8492
rect 6052 8452 6368 8480
rect 6052 8440 6058 8452
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 6472 8480 6500 8520
rect 10042 8508 10048 8520
rect 10100 8508 10106 8560
rect 11606 8508 11612 8560
rect 11664 8548 11670 8560
rect 12710 8548 12716 8560
rect 11664 8520 12716 8548
rect 11664 8508 11670 8520
rect 12710 8508 12716 8520
rect 12768 8508 12774 8560
rect 15010 8548 15016 8560
rect 14971 8520 15016 8548
rect 15010 8508 15016 8520
rect 15068 8508 15074 8560
rect 6472 8452 6960 8480
rect 5000 8384 5856 8412
rect 3234 8304 3240 8356
rect 3292 8353 3298 8356
rect 3292 8347 3356 8353
rect 3292 8313 3310 8347
rect 3344 8313 3356 8347
rect 4982 8344 4988 8356
rect 3292 8307 3356 8313
rect 3436 8316 4988 8344
rect 3292 8304 3298 8307
rect 1581 8279 1639 8285
rect 1581 8245 1593 8279
rect 1627 8276 1639 8279
rect 2314 8276 2320 8288
rect 1627 8248 2320 8276
rect 1627 8245 1639 8248
rect 1581 8239 1639 8245
rect 2314 8236 2320 8248
rect 2372 8236 2378 8288
rect 2777 8279 2835 8285
rect 2777 8245 2789 8279
rect 2823 8276 2835 8279
rect 3436 8276 3464 8316
rect 4982 8304 4988 8316
rect 5040 8304 5046 8356
rect 5160 8347 5218 8353
rect 5160 8313 5172 8347
rect 5206 8344 5218 8347
rect 5534 8344 5540 8356
rect 5206 8316 5540 8344
rect 5206 8313 5218 8316
rect 5160 8307 5218 8313
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 5828 8344 5856 8384
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 6822 8412 6828 8424
rect 5960 8384 6500 8412
rect 6783 8384 6828 8412
rect 5960 8372 5966 8384
rect 6178 8344 6184 8356
rect 5828 8316 6184 8344
rect 6178 8304 6184 8316
rect 6236 8304 6242 8356
rect 2823 8248 3464 8276
rect 2823 8245 2835 8248
rect 2777 8239 2835 8245
rect 4246 8236 4252 8288
rect 4304 8276 4310 8288
rect 6362 8276 6368 8288
rect 4304 8248 6368 8276
rect 4304 8236 4310 8248
rect 6362 8236 6368 8248
rect 6420 8236 6426 8288
rect 6472 8276 6500 8384
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 6932 8412 6960 8452
rect 8018 8440 8024 8492
rect 8076 8480 8082 8492
rect 8386 8480 8392 8492
rect 8076 8452 8392 8480
rect 8076 8440 8082 8452
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8662 8480 8668 8492
rect 8623 8452 8668 8480
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 9766 8440 9772 8492
rect 9824 8480 9830 8492
rect 9950 8480 9956 8492
rect 9824 8452 9956 8480
rect 9824 8440 9830 8452
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 11514 8440 11520 8492
rect 11572 8480 11578 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 11572 8452 13001 8480
rect 11572 8440 11578 8452
rect 12989 8449 13001 8452
rect 13035 8480 13047 8483
rect 13814 8480 13820 8492
rect 13035 8452 13820 8480
rect 13035 8449 13047 8452
rect 12989 8443 13047 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 14277 8483 14335 8489
rect 14277 8449 14289 8483
rect 14323 8480 14335 8483
rect 14458 8480 14464 8492
rect 14323 8452 14464 8480
rect 14323 8449 14335 8452
rect 14277 8443 14335 8449
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 8921 8415 8979 8421
rect 8921 8412 8933 8415
rect 6932 8384 8933 8412
rect 8921 8381 8933 8384
rect 8967 8412 8979 8415
rect 9214 8412 9220 8424
rect 8967 8384 9220 8412
rect 8967 8381 8979 8384
rect 8921 8375 8979 8381
rect 9214 8372 9220 8384
rect 9272 8372 9278 8424
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 10505 8415 10563 8421
rect 10505 8412 10517 8415
rect 9732 8384 10517 8412
rect 9732 8372 9738 8384
rect 10505 8381 10517 8384
rect 10551 8412 10563 8415
rect 10551 8384 11468 8412
rect 10551 8381 10563 8384
rect 10505 8375 10563 8381
rect 11440 8356 11468 8384
rect 12342 8372 12348 8424
rect 12400 8412 12406 8424
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12400 8384 12909 8412
rect 12400 8372 12406 8384
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 13078 8372 13084 8424
rect 13136 8412 13142 8424
rect 14829 8415 14887 8421
rect 13136 8384 14228 8412
rect 13136 8372 13142 8384
rect 7070 8347 7128 8353
rect 7070 8344 7082 8347
rect 6739 8316 7082 8344
rect 6739 8276 6767 8316
rect 7070 8313 7082 8316
rect 7116 8313 7128 8347
rect 7070 8307 7128 8313
rect 7190 8304 7196 8356
rect 7248 8344 7254 8356
rect 7248 8316 8156 8344
rect 7248 8304 7254 8316
rect 6472 8248 6767 8276
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 7926 8276 7932 8288
rect 6972 8248 7932 8276
rect 6972 8236 6978 8248
rect 7926 8236 7932 8248
rect 7984 8236 7990 8288
rect 8128 8276 8156 8316
rect 8202 8304 8208 8356
rect 8260 8344 8266 8356
rect 10594 8344 10600 8356
rect 8260 8316 10600 8344
rect 8260 8304 8266 8316
rect 10594 8304 10600 8316
rect 10652 8304 10658 8356
rect 10686 8304 10692 8356
rect 10744 8353 10750 8356
rect 10744 8347 10808 8353
rect 10744 8313 10762 8347
rect 10796 8313 10808 8347
rect 10744 8307 10808 8313
rect 10744 8304 10750 8307
rect 11422 8304 11428 8356
rect 11480 8304 11486 8356
rect 12805 8347 12863 8353
rect 12805 8313 12817 8347
rect 12851 8344 12863 8347
rect 13188 8344 13216 8384
rect 12851 8316 13216 8344
rect 12851 8313 12863 8316
rect 12805 8307 12863 8313
rect 13814 8304 13820 8356
rect 13872 8344 13878 8356
rect 14093 8347 14151 8353
rect 14093 8344 14105 8347
rect 13872 8316 14105 8344
rect 13872 8304 13878 8316
rect 14093 8313 14105 8316
rect 14139 8313 14151 8347
rect 14093 8307 14151 8313
rect 8754 8276 8760 8288
rect 8128 8248 8760 8276
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 11606 8276 11612 8288
rect 9088 8248 11612 8276
rect 9088 8236 9094 8248
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 12158 8236 12164 8288
rect 12216 8276 12222 8288
rect 12342 8276 12348 8288
rect 12216 8248 12348 8276
rect 12216 8236 12222 8248
rect 12342 8236 12348 8248
rect 12400 8236 12406 8288
rect 13998 8276 14004 8288
rect 13959 8248 14004 8276
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 14200 8276 14228 8384
rect 14829 8381 14841 8415
rect 14875 8412 14887 8415
rect 15470 8412 15476 8424
rect 14875 8384 15476 8412
rect 14875 8381 14887 8384
rect 14829 8375 14887 8381
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 14458 8276 14464 8288
rect 14200 8248 14464 8276
rect 14458 8236 14464 8248
rect 14516 8236 14522 8288
rect 1104 8186 15824 8208
rect 1104 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 6104 8186
rect 6156 8134 10843 8186
rect 10895 8134 10907 8186
rect 10959 8134 10971 8186
rect 11023 8134 11035 8186
rect 11087 8134 15824 8186
rect 1104 8112 15824 8134
rect 4893 8075 4951 8081
rect 4893 8041 4905 8075
rect 4939 8072 4951 8075
rect 4939 8044 5856 8072
rect 4939 8041 4951 8044
rect 4893 8035 4951 8041
rect 5074 8004 5080 8016
rect 1412 7976 5080 8004
rect 1412 7945 1440 7976
rect 5074 7964 5080 7976
rect 5132 7964 5138 8016
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7905 1455 7939
rect 1397 7899 1455 7905
rect 2400 7939 2458 7945
rect 2400 7905 2412 7939
rect 2446 7936 2458 7939
rect 2682 7936 2688 7948
rect 2446 7908 2688 7936
rect 2446 7905 2458 7908
rect 2400 7899 2458 7905
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 4985 7939 5043 7945
rect 4985 7905 4997 7939
rect 5031 7936 5043 7939
rect 5626 7936 5632 7948
rect 5031 7908 5632 7936
rect 5031 7905 5043 7908
rect 4985 7899 5043 7905
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 5828 7936 5856 8044
rect 6362 8032 6368 8084
rect 6420 8072 6426 8084
rect 6914 8072 6920 8084
rect 6420 8044 6920 8072
rect 6420 8032 6426 8044
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 7101 8075 7159 8081
rect 7101 8072 7113 8075
rect 7024 8044 7113 8072
rect 5994 8013 6000 8016
rect 5988 7967 6000 8013
rect 6052 8004 6058 8016
rect 6052 7976 6088 8004
rect 5994 7964 6000 7967
rect 6052 7964 6058 7976
rect 6730 7964 6736 8016
rect 6788 8004 6794 8016
rect 7024 8004 7052 8044
rect 7101 8041 7113 8044
rect 7147 8041 7159 8075
rect 7742 8072 7748 8084
rect 7101 8035 7159 8041
rect 7484 8044 7748 8072
rect 7484 8004 7512 8044
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 7929 8075 7987 8081
rect 7929 8041 7941 8075
rect 7975 8072 7987 8075
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 7975 8044 8033 8072
rect 7975 8041 7987 8044
rect 7929 8035 7987 8041
rect 8021 8041 8033 8044
rect 8067 8072 8079 8075
rect 8202 8072 8208 8084
rect 8067 8044 8208 8072
rect 8067 8041 8079 8044
rect 8021 8035 8079 8041
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 8386 8032 8392 8084
rect 8444 8072 8450 8084
rect 8757 8075 8815 8081
rect 8757 8072 8769 8075
rect 8444 8044 8769 8072
rect 8444 8032 8450 8044
rect 8757 8041 8769 8044
rect 8803 8041 8815 8075
rect 8757 8035 8815 8041
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 11517 8075 11575 8081
rect 11517 8072 11529 8075
rect 9539 8044 11529 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 11517 8041 11529 8044
rect 11563 8041 11575 8075
rect 11517 8035 11575 8041
rect 11790 8032 11796 8084
rect 11848 8072 11854 8084
rect 11885 8075 11943 8081
rect 11885 8072 11897 8075
rect 11848 8044 11897 8072
rect 11848 8032 11854 8044
rect 11885 8041 11897 8044
rect 11931 8041 11943 8075
rect 11885 8035 11943 8041
rect 13909 8075 13967 8081
rect 13909 8041 13921 8075
rect 13955 8072 13967 8075
rect 13998 8072 14004 8084
rect 13955 8044 14004 8072
rect 13955 8041 13967 8044
rect 13909 8035 13967 8041
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 8662 8004 8668 8016
rect 6788 7976 7052 8004
rect 7116 7976 7512 8004
rect 7760 7976 8668 8004
rect 6788 7964 6794 7976
rect 5828 7908 6875 7936
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5258 7868 5264 7880
rect 5215 7840 5264 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 1486 7692 1492 7744
rect 1544 7732 1550 7744
rect 1581 7735 1639 7741
rect 1581 7732 1593 7735
rect 1544 7704 1593 7732
rect 1544 7692 1550 7704
rect 1581 7701 1593 7704
rect 1627 7701 1639 7735
rect 2148 7732 2176 7831
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5718 7868 5724 7880
rect 5679 7840 5724 7868
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 6847 7868 6875 7908
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7116 7936 7144 7976
rect 7760 7948 7788 7976
rect 8662 7964 8668 7976
rect 8720 7964 8726 8016
rect 9125 8007 9183 8013
rect 8772 7976 8975 8004
rect 6972 7908 7144 7936
rect 6972 7896 6978 7908
rect 7742 7896 7748 7948
rect 7800 7896 7806 7948
rect 8018 7896 8024 7948
rect 8076 7936 8082 7948
rect 8772 7936 8800 7976
rect 8076 7908 8800 7936
rect 8947 7936 8975 7976
rect 9125 7973 9137 8007
rect 9171 8004 9183 8007
rect 14277 8007 14335 8013
rect 14277 8004 14289 8007
rect 9171 7976 14289 8004
rect 9171 7973 9183 7976
rect 9125 7967 9183 7973
rect 14277 7973 14289 7976
rect 14323 7973 14335 8007
rect 14277 7967 14335 7973
rect 8947 7908 9536 7936
rect 8076 7896 8082 7908
rect 8846 7868 8852 7880
rect 6847 7840 8616 7868
rect 8807 7840 8852 7868
rect 3513 7803 3571 7809
rect 3513 7769 3525 7803
rect 3559 7800 3571 7803
rect 4246 7800 4252 7812
rect 3559 7772 4252 7800
rect 3559 7769 3571 7772
rect 3513 7763 3571 7769
rect 4246 7760 4252 7772
rect 4304 7800 4310 7812
rect 8018 7800 8024 7812
rect 4304 7772 5764 7800
rect 4304 7760 4310 7772
rect 2866 7732 2872 7744
rect 2148 7704 2872 7732
rect 1581 7695 1639 7701
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 4522 7732 4528 7744
rect 4483 7704 4528 7732
rect 4522 7692 4528 7704
rect 4580 7692 4586 7744
rect 5736 7732 5764 7772
rect 6656 7772 8024 7800
rect 6656 7732 6684 7772
rect 8018 7760 8024 7772
rect 8076 7760 8082 7812
rect 8588 7800 8616 7840
rect 8846 7828 8852 7840
rect 8904 7868 8910 7880
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 8904 7840 9413 7868
rect 8904 7828 8910 7840
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 9508 7868 9536 7908
rect 9582 7896 9588 7948
rect 9640 7936 9646 7948
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 9640 7908 9689 7936
rect 9640 7896 9646 7908
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9933 7939 9991 7945
rect 9933 7936 9945 7939
rect 9677 7899 9735 7905
rect 9784 7908 9945 7936
rect 9784 7868 9812 7908
rect 9933 7905 9945 7908
rect 9979 7905 9991 7939
rect 9933 7899 9991 7905
rect 10318 7896 10324 7948
rect 10376 7936 10382 7948
rect 10870 7936 10876 7948
rect 10376 7908 10876 7936
rect 10376 7896 10382 7908
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 11974 7936 11980 7948
rect 11935 7908 11980 7936
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 12894 7896 12900 7948
rect 12952 7936 12958 7948
rect 13081 7939 13139 7945
rect 13081 7936 13093 7939
rect 12952 7908 13093 7936
rect 12952 7896 12958 7908
rect 13081 7905 13093 7908
rect 13127 7905 13139 7939
rect 13722 7936 13728 7948
rect 13081 7899 13139 7905
rect 13188 7908 13728 7936
rect 9508 7840 9812 7868
rect 9401 7831 9459 7837
rect 10962 7828 10968 7880
rect 11020 7868 11026 7880
rect 11514 7868 11520 7880
rect 11020 7840 11520 7868
rect 11020 7828 11026 7840
rect 11514 7828 11520 7840
rect 11572 7868 11578 7880
rect 12066 7868 12072 7880
rect 11572 7840 12072 7868
rect 11572 7828 11578 7840
rect 12066 7828 12072 7840
rect 12124 7828 12130 7880
rect 12158 7828 12164 7880
rect 12216 7868 12222 7880
rect 13188 7877 13216 7908
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 13173 7871 13231 7877
rect 13173 7868 13185 7871
rect 12216 7840 13185 7868
rect 12216 7828 12222 7840
rect 13173 7837 13185 7840
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7837 13323 7871
rect 13265 7831 13323 7837
rect 9493 7803 9551 7809
rect 9493 7800 9505 7803
rect 8588 7772 9505 7800
rect 9493 7769 9505 7772
rect 9539 7769 9551 7803
rect 13280 7800 13308 7831
rect 14274 7828 14280 7880
rect 14332 7868 14338 7880
rect 14369 7871 14427 7877
rect 14369 7868 14381 7871
rect 14332 7840 14381 7868
rect 14332 7828 14338 7840
rect 14369 7837 14381 7840
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 9493 7763 9551 7769
rect 10704 7772 13308 7800
rect 5736 7704 6684 7732
rect 8297 7735 8355 7741
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 8662 7732 8668 7744
rect 8343 7704 8668 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 9030 7732 9036 7744
rect 8812 7704 9036 7732
rect 8812 7692 8818 7704
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 10042 7732 10048 7744
rect 9447 7704 10048 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 10042 7692 10048 7704
rect 10100 7732 10106 7744
rect 10704 7732 10732 7772
rect 14182 7760 14188 7812
rect 14240 7800 14246 7812
rect 14476 7800 14504 7831
rect 14240 7772 14504 7800
rect 14240 7760 14246 7772
rect 10100 7704 10732 7732
rect 10100 7692 10106 7704
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 10836 7704 11069 7732
rect 10836 7692 10842 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 12526 7692 12532 7744
rect 12584 7732 12590 7744
rect 12713 7735 12771 7741
rect 12713 7732 12725 7735
rect 12584 7704 12725 7732
rect 12584 7692 12590 7704
rect 12713 7701 12725 7704
rect 12759 7701 12771 7735
rect 12713 7695 12771 7701
rect 1104 7642 15824 7664
rect 1104 7590 3447 7642
rect 3499 7590 3511 7642
rect 3563 7590 3575 7642
rect 3627 7590 3639 7642
rect 3691 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 13308 7642
rect 13360 7590 13372 7642
rect 13424 7590 13436 7642
rect 13488 7590 13500 7642
rect 13552 7590 15824 7642
rect 1104 7568 15824 7590
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 2924 7500 3096 7528
rect 2924 7488 2930 7500
rect 1857 7463 1915 7469
rect 1857 7429 1869 7463
rect 1903 7460 1915 7463
rect 1903 7432 2912 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 2884 7404 2912 7432
rect 3068 7404 3096 7500
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 4433 7531 4491 7537
rect 4433 7528 4445 7531
rect 3292 7500 4445 7528
rect 3292 7488 3298 7500
rect 4433 7497 4445 7500
rect 4479 7528 4491 7531
rect 5258 7528 5264 7540
rect 4479 7500 5264 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5626 7488 5632 7540
rect 5684 7528 5690 7540
rect 7558 7528 7564 7540
rect 5684 7500 7564 7528
rect 5684 7488 5690 7500
rect 7558 7488 7564 7500
rect 7616 7488 7622 7540
rect 7834 7488 7840 7540
rect 7892 7528 7898 7540
rect 7892 7500 8708 7528
rect 7892 7488 7898 7500
rect 5902 7420 5908 7472
rect 5960 7460 5966 7472
rect 8205 7463 8263 7469
rect 5960 7432 6868 7460
rect 5960 7420 5966 7432
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 2590 7392 2596 7404
rect 2547 7364 2596 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2590 7352 2596 7364
rect 2648 7352 2654 7404
rect 2866 7352 2872 7404
rect 2924 7352 2930 7404
rect 3050 7392 3056 7404
rect 3011 7364 3056 7392
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 4890 7392 4896 7404
rect 4851 7364 4896 7392
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 6840 7392 6868 7432
rect 8205 7429 8217 7463
rect 8251 7460 8263 7463
rect 8294 7460 8300 7472
rect 8251 7432 8300 7460
rect 8251 7429 8263 7432
rect 8205 7423 8263 7429
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 8680 7401 8708 7500
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 9950 7528 9956 7540
rect 9640 7500 9956 7528
rect 9640 7488 9646 7500
rect 9950 7488 9956 7500
rect 10008 7528 10014 7540
rect 10008 7500 11928 7528
rect 10008 7488 10014 7500
rect 10962 7460 10968 7472
rect 9876 7432 10968 7460
rect 8665 7395 8723 7401
rect 6840 7364 6960 7392
rect 1118 7284 1124 7336
rect 1176 7324 1182 7336
rect 3786 7324 3792 7336
rect 1176 7296 3792 7324
rect 1176 7284 1182 7296
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 4540 7296 5580 7324
rect 3320 7259 3378 7265
rect 3320 7225 3332 7259
rect 3366 7256 3378 7259
rect 4540 7256 4568 7296
rect 3366 7228 4568 7256
rect 3366 7225 3378 7228
rect 3320 7219 3378 7225
rect 4614 7216 4620 7268
rect 4672 7256 4678 7268
rect 5160 7259 5218 7265
rect 5160 7256 5172 7259
rect 4672 7228 5172 7256
rect 4672 7216 4678 7228
rect 5160 7225 5172 7228
rect 5206 7256 5218 7259
rect 5350 7256 5356 7268
rect 5206 7228 5356 7256
rect 5206 7225 5218 7228
rect 5160 7219 5218 7225
rect 5350 7216 5356 7228
rect 5408 7216 5414 7268
rect 5552 7256 5580 7296
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 6638 7324 6644 7336
rect 5684 7296 6644 7324
rect 5684 7284 5690 7296
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 6829 7324 6835 7336
rect 6790 7296 6835 7324
rect 6829 7284 6835 7296
rect 6887 7284 6893 7336
rect 6932 7324 6960 7364
rect 7843 7364 8524 7392
rect 7843 7324 7871 7364
rect 6932 7296 7871 7324
rect 8297 7327 8355 7333
rect 8297 7293 8309 7327
rect 8343 7324 8355 7327
rect 8386 7324 8392 7336
rect 8343 7296 8392 7324
rect 8343 7293 8355 7296
rect 8297 7287 8355 7293
rect 8386 7284 8392 7296
rect 8444 7284 8450 7336
rect 8496 7324 8524 7364
rect 8665 7361 8677 7395
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 9398 7324 9404 7336
rect 8496 7296 9404 7324
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 7092 7259 7150 7265
rect 5552 7228 7052 7256
rect 2222 7188 2228 7200
rect 2183 7160 2228 7188
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 5626 7188 5632 7200
rect 2363 7160 5632 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 6270 7188 6276 7200
rect 6231 7160 6276 7188
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 7024 7188 7052 7228
rect 7092 7225 7104 7259
rect 7138 7256 7150 7259
rect 7374 7256 7380 7268
rect 7138 7228 7380 7256
rect 7138 7225 7150 7228
rect 7092 7219 7150 7225
rect 7374 7216 7380 7228
rect 7432 7216 7438 7268
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 8662 7256 8668 7268
rect 7616 7228 8668 7256
rect 7616 7216 7622 7228
rect 8662 7216 8668 7228
rect 8720 7216 8726 7268
rect 8932 7259 8990 7265
rect 8932 7225 8944 7259
rect 8978 7256 8990 7259
rect 9030 7256 9036 7268
rect 8978 7228 9036 7256
rect 8978 7225 8990 7228
rect 8932 7219 8990 7225
rect 9030 7216 9036 7228
rect 9088 7216 9094 7268
rect 9122 7216 9128 7268
rect 9180 7256 9186 7268
rect 9582 7256 9588 7268
rect 9180 7228 9588 7256
rect 9180 7216 9186 7228
rect 9582 7216 9588 7228
rect 9640 7216 9646 7268
rect 7926 7188 7932 7200
rect 7024 7160 7932 7188
rect 7926 7148 7932 7160
rect 7984 7188 7990 7200
rect 9876 7188 9904 7432
rect 10962 7420 10968 7432
rect 11020 7460 11026 7472
rect 11900 7460 11928 7500
rect 11974 7488 11980 7540
rect 12032 7528 12038 7540
rect 12437 7531 12495 7537
rect 12437 7528 12449 7531
rect 12032 7500 12449 7528
rect 12032 7488 12038 7500
rect 12437 7497 12449 7500
rect 12483 7497 12495 7531
rect 12437 7491 12495 7497
rect 13633 7531 13691 7537
rect 13633 7497 13645 7531
rect 13679 7528 13691 7531
rect 14366 7528 14372 7540
rect 13679 7500 14372 7528
rect 13679 7497 13691 7500
rect 13633 7491 13691 7497
rect 14366 7488 14372 7500
rect 14424 7488 14430 7540
rect 13078 7460 13084 7472
rect 11020 7432 11100 7460
rect 11900 7432 13084 7460
rect 11020 7420 11026 7432
rect 9950 7352 9956 7404
rect 10008 7392 10014 7404
rect 10778 7392 10784 7404
rect 10008 7364 10784 7392
rect 10008 7352 10014 7364
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 11072 7401 11100 7432
rect 13078 7420 13084 7432
rect 13136 7420 13142 7472
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7361 11115 7395
rect 11974 7392 11980 7404
rect 11057 7355 11115 7361
rect 11440 7364 11980 7392
rect 10965 7327 11023 7333
rect 10965 7293 10977 7327
rect 11011 7324 11023 7327
rect 11330 7324 11336 7336
rect 11011 7296 11336 7324
rect 11011 7293 11023 7296
rect 10965 7287 11023 7293
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 10778 7216 10784 7268
rect 10836 7256 10842 7268
rect 10873 7259 10931 7265
rect 10873 7256 10885 7259
rect 10836 7228 10885 7256
rect 10836 7216 10842 7228
rect 10873 7225 10885 7228
rect 10919 7225 10931 7259
rect 10873 7219 10931 7225
rect 11054 7216 11060 7268
rect 11112 7256 11118 7268
rect 11440 7256 11468 7364
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12124 7364 13001 7392
rect 12124 7352 12130 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 14182 7392 14188 7404
rect 12989 7355 13047 7361
rect 13096 7364 14188 7392
rect 11606 7284 11612 7336
rect 11664 7324 11670 7336
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 11664 7296 12817 7324
rect 11664 7284 11670 7296
rect 12805 7293 12817 7296
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 11112 7228 11468 7256
rect 11112 7216 11118 7228
rect 12066 7216 12072 7268
rect 12124 7256 12130 7268
rect 13096 7256 13124 7364
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 14826 7324 14832 7336
rect 14787 7296 14832 7324
rect 14826 7284 14832 7296
rect 14884 7284 14890 7336
rect 12124 7228 13124 7256
rect 12124 7216 12130 7228
rect 13906 7216 13912 7268
rect 13964 7256 13970 7268
rect 14093 7259 14151 7265
rect 14093 7256 14105 7259
rect 13964 7228 14105 7256
rect 13964 7216 13970 7228
rect 14093 7225 14105 7228
rect 14139 7225 14151 7259
rect 14093 7219 14151 7225
rect 7984 7160 9904 7188
rect 10045 7191 10103 7197
rect 7984 7148 7990 7160
rect 10045 7157 10057 7191
rect 10091 7188 10103 7191
rect 10134 7188 10140 7200
rect 10091 7160 10140 7188
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 10226 7148 10232 7200
rect 10284 7188 10290 7200
rect 10505 7191 10563 7197
rect 10505 7188 10517 7191
rect 10284 7160 10517 7188
rect 10284 7148 10290 7160
rect 10505 7157 10517 7160
rect 10551 7157 10563 7191
rect 10505 7151 10563 7157
rect 10594 7148 10600 7200
rect 10652 7188 10658 7200
rect 11330 7188 11336 7200
rect 10652 7160 11336 7188
rect 10652 7148 10658 7160
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11422 7148 11428 7200
rect 11480 7188 11486 7200
rect 11701 7191 11759 7197
rect 11701 7188 11713 7191
rect 11480 7160 11713 7188
rect 11480 7148 11486 7160
rect 11701 7157 11713 7160
rect 11747 7157 11759 7191
rect 11701 7151 11759 7157
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12897 7191 12955 7197
rect 12897 7188 12909 7191
rect 12032 7160 12909 7188
rect 12032 7148 12038 7160
rect 12897 7157 12909 7160
rect 12943 7157 12955 7191
rect 13998 7188 14004 7200
rect 13959 7160 14004 7188
rect 12897 7151 12955 7157
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 15013 7191 15071 7197
rect 15013 7188 15025 7191
rect 14424 7160 15025 7188
rect 14424 7148 14430 7160
rect 15013 7157 15025 7160
rect 15059 7157 15071 7191
rect 15013 7151 15071 7157
rect 1104 7098 15824 7120
rect 1104 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 6104 7098
rect 6156 7046 10843 7098
rect 10895 7046 10907 7098
rect 10959 7046 10971 7098
rect 11023 7046 11035 7098
rect 11087 7046 15824 7098
rect 1104 7024 15824 7046
rect 2222 6944 2228 6996
rect 2280 6984 2286 6996
rect 6730 6984 6736 6996
rect 2280 6956 6736 6984
rect 2280 6944 2286 6956
rect 6730 6944 6736 6956
rect 6788 6944 6794 6996
rect 7190 6984 7196 6996
rect 7151 6956 7196 6984
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 8110 6984 8116 6996
rect 7616 6956 8116 6984
rect 7616 6944 7622 6956
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 9493 6987 9551 6993
rect 9493 6984 9505 6987
rect 8444 6956 9505 6984
rect 8444 6944 8450 6956
rect 9493 6953 9505 6956
rect 9539 6953 9551 6987
rect 9493 6947 9551 6953
rect 10045 6987 10103 6993
rect 10045 6953 10057 6987
rect 10091 6984 10103 6987
rect 10410 6984 10416 6996
rect 10091 6956 10416 6984
rect 10091 6953 10103 6956
rect 10045 6947 10103 6953
rect 10410 6944 10416 6956
rect 10468 6944 10474 6996
rect 10594 6944 10600 6996
rect 10652 6984 10658 6996
rect 12158 6984 12164 6996
rect 10652 6956 12164 6984
rect 10652 6944 10658 6956
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 12437 6987 12495 6993
rect 12437 6953 12449 6987
rect 12483 6984 12495 6987
rect 12618 6984 12624 6996
rect 12483 6956 12624 6984
rect 12483 6953 12495 6956
rect 12437 6947 12495 6953
rect 12618 6944 12624 6956
rect 12676 6984 12682 6996
rect 14182 6984 14188 6996
rect 12676 6956 14188 6984
rect 12676 6944 12682 6956
rect 14182 6944 14188 6956
rect 14240 6944 14246 6996
rect 14645 6987 14703 6993
rect 14645 6953 14657 6987
rect 14691 6953 14703 6987
rect 14645 6947 14703 6953
rect 2590 6916 2596 6928
rect 2148 6888 2596 6916
rect 1302 6808 1308 6860
rect 1360 6848 1366 6860
rect 2148 6857 2176 6888
rect 2590 6876 2596 6888
rect 2648 6876 2654 6928
rect 4893 6919 4951 6925
rect 4893 6885 4905 6919
rect 4939 6916 4951 6919
rect 10226 6916 10232 6928
rect 4939 6888 10232 6916
rect 4939 6885 4951 6888
rect 4893 6879 4951 6885
rect 10226 6876 10232 6888
rect 10284 6876 10290 6928
rect 1397 6851 1455 6857
rect 1397 6848 1409 6851
rect 1360 6820 1409 6848
rect 1360 6808 1366 6820
rect 1397 6817 1409 6820
rect 1443 6817 1455 6851
rect 1397 6811 1455 6817
rect 2133 6851 2191 6857
rect 2133 6817 2145 6851
rect 2179 6817 2191 6851
rect 2133 6811 2191 6817
rect 2400 6851 2458 6857
rect 2400 6817 2412 6851
rect 2446 6848 2458 6851
rect 3786 6848 3792 6860
rect 2446 6820 3792 6848
rect 2446 6817 2458 6820
rect 2400 6811 2458 6817
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 6069 6851 6127 6857
rect 6069 6848 6081 6851
rect 4120 6820 6081 6848
rect 4120 6808 4126 6820
rect 6069 6817 6081 6820
rect 6115 6848 6127 6851
rect 6914 6848 6920 6860
rect 6115 6820 6920 6848
rect 6115 6817 6127 6820
rect 6069 6811 6127 6817
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 7920 6851 7978 6857
rect 7920 6817 7932 6851
rect 7966 6848 7978 6851
rect 9122 6848 9128 6860
rect 7966 6820 9128 6848
rect 7966 6817 7978 6820
rect 7920 6811 7978 6817
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 10137 6851 10195 6857
rect 10137 6848 10149 6851
rect 9456 6820 10149 6848
rect 9456 6808 9462 6820
rect 10137 6817 10149 6820
rect 10183 6817 10195 6851
rect 10428 6848 10456 6944
rect 11054 6876 11060 6928
rect 11112 6916 11118 6928
rect 11241 6919 11299 6925
rect 11241 6916 11253 6919
rect 11112 6888 11253 6916
rect 11112 6876 11118 6888
rect 11241 6885 11253 6888
rect 11287 6916 11299 6919
rect 11287 6888 12664 6916
rect 11287 6885 11299 6888
rect 11241 6879 11299 6885
rect 11606 6848 11612 6860
rect 10428 6820 11612 6848
rect 10137 6811 10195 6817
rect 11606 6808 11612 6820
rect 11664 6808 11670 6860
rect 12158 6808 12164 6860
rect 12216 6848 12222 6860
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12216 6820 12541 6848
rect 12216 6808 12222 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12636 6848 12664 6888
rect 12710 6876 12716 6928
rect 12768 6916 12774 6928
rect 14660 6916 14688 6947
rect 12768 6888 14688 6916
rect 12768 6876 12774 6888
rect 12894 6848 12900 6860
rect 12636 6820 12900 6848
rect 12529 6811 12587 6817
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13630 6848 13636 6860
rect 13591 6820 13636 6848
rect 13630 6808 13636 6820
rect 13688 6808 13694 6860
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 14461 6851 14519 6857
rect 14461 6848 14473 6851
rect 14148 6820 14473 6848
rect 14148 6808 14154 6820
rect 14461 6817 14473 6820
rect 14507 6817 14519 6851
rect 14461 6811 14519 6817
rect 4982 6780 4988 6792
rect 4943 6752 4988 6780
rect 4982 6740 4988 6752
rect 5040 6740 5046 6792
rect 5166 6780 5172 6792
rect 5079 6752 5172 6780
rect 5166 6740 5172 6752
rect 5224 6780 5230 6792
rect 5224 6752 5764 6780
rect 5224 6740 5230 6752
rect 3513 6715 3571 6721
rect 3513 6681 3525 6715
rect 3559 6712 3571 6715
rect 5626 6712 5632 6724
rect 3559 6684 5632 6712
rect 3559 6681 3571 6684
rect 3513 6675 3571 6681
rect 5626 6672 5632 6684
rect 5684 6672 5690 6724
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 4525 6647 4583 6653
rect 4525 6613 4537 6647
rect 4571 6644 4583 6647
rect 4890 6644 4896 6656
rect 4571 6616 4896 6644
rect 4571 6613 4583 6616
rect 4525 6607 4583 6613
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 5736 6644 5764 6752
rect 5810 6740 5816 6792
rect 5868 6780 5874 6792
rect 7650 6780 7656 6792
rect 5868 6752 5913 6780
rect 7611 6752 7656 6780
rect 5868 6740 5874 6752
rect 7650 6740 7656 6752
rect 7708 6740 7714 6792
rect 8662 6740 8668 6792
rect 8720 6740 8726 6792
rect 9766 6780 9772 6792
rect 9048 6752 9772 6780
rect 6914 6672 6920 6724
rect 6972 6712 6978 6724
rect 8680 6712 8708 6740
rect 8846 6712 8852 6724
rect 6972 6684 7236 6712
rect 8680 6684 8852 6712
rect 6972 6672 6978 6684
rect 7098 6644 7104 6656
rect 5736 6616 7104 6644
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7208 6644 7236 6684
rect 8846 6672 8852 6684
rect 8904 6672 8910 6724
rect 9048 6721 9076 6752
rect 9766 6740 9772 6752
rect 9824 6780 9830 6792
rect 9824 6752 9904 6780
rect 9824 6740 9830 6752
rect 9033 6715 9091 6721
rect 9033 6681 9045 6715
rect 9079 6681 9091 6715
rect 9033 6675 9091 6681
rect 9306 6672 9312 6724
rect 9364 6712 9370 6724
rect 9493 6715 9551 6721
rect 9493 6712 9505 6715
rect 9364 6684 9505 6712
rect 9364 6672 9370 6684
rect 9493 6681 9505 6684
rect 9539 6681 9551 6715
rect 9493 6675 9551 6681
rect 9674 6672 9680 6724
rect 9732 6712 9738 6724
rect 9876 6712 9904 6752
rect 10042 6740 10048 6792
rect 10100 6780 10106 6792
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 10100 6752 10241 6780
rect 10100 6740 10106 6752
rect 10229 6749 10241 6752
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 10594 6740 10600 6792
rect 10652 6780 10658 6792
rect 11333 6783 11391 6789
rect 11333 6780 11345 6783
rect 10652 6752 11345 6780
rect 10652 6740 10658 6752
rect 11333 6749 11345 6752
rect 11379 6749 11391 6783
rect 11333 6743 11391 6749
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 11698 6780 11704 6792
rect 11563 6752 11704 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 12618 6780 12624 6792
rect 12579 6752 12624 6780
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 13722 6780 13728 6792
rect 13683 6752 13728 6780
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 13906 6780 13912 6792
rect 13867 6752 13912 6780
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 12250 6712 12256 6724
rect 9732 6684 9777 6712
rect 9876 6684 12256 6712
rect 9732 6672 9738 6684
rect 12250 6672 12256 6684
rect 12308 6672 12314 6724
rect 12986 6672 12992 6724
rect 13044 6712 13050 6724
rect 13998 6712 14004 6724
rect 13044 6684 14004 6712
rect 13044 6672 13050 6684
rect 13998 6672 14004 6684
rect 14056 6672 14062 6724
rect 10873 6647 10931 6653
rect 10873 6644 10885 6647
rect 7208 6616 10885 6644
rect 10873 6613 10885 6616
rect 10919 6613 10931 6647
rect 10873 6607 10931 6613
rect 11974 6604 11980 6656
rect 12032 6644 12038 6656
rect 12069 6647 12127 6653
rect 12069 6644 12081 6647
rect 12032 6616 12081 6644
rect 12032 6604 12038 6616
rect 12069 6613 12081 6616
rect 12115 6613 12127 6647
rect 12069 6607 12127 6613
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 13265 6647 13323 6653
rect 13265 6644 13277 6647
rect 12860 6616 13277 6644
rect 12860 6604 12866 6616
rect 13265 6613 13277 6616
rect 13311 6613 13323 6647
rect 13265 6607 13323 6613
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 1854 6440 1860 6452
rect 1815 6412 1860 6440
rect 1854 6400 1860 6412
rect 1912 6400 1918 6452
rect 3786 6400 3792 6452
rect 3844 6440 3850 6452
rect 4433 6443 4491 6449
rect 4433 6440 4445 6443
rect 3844 6412 4445 6440
rect 3844 6400 3850 6412
rect 4433 6409 4445 6412
rect 4479 6440 4491 6443
rect 4479 6412 7788 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 3050 6332 3056 6384
rect 3108 6332 3114 6384
rect 5902 6332 5908 6384
rect 5960 6372 5966 6384
rect 6270 6372 6276 6384
rect 5960 6344 6276 6372
rect 5960 6332 5966 6344
rect 6270 6332 6276 6344
rect 6328 6332 6334 6384
rect 7760 6372 7788 6412
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 8205 6443 8263 6449
rect 8205 6440 8217 6443
rect 7984 6412 8217 6440
rect 7984 6400 7990 6412
rect 8205 6409 8217 6412
rect 8251 6409 8263 6443
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 8205 6403 8263 6409
rect 8680 6412 10057 6440
rect 8386 6372 8392 6384
rect 7760 6344 8392 6372
rect 8386 6332 8392 6344
rect 8444 6332 8450 6384
rect 8570 6332 8576 6384
rect 8628 6372 8634 6384
rect 8680 6372 8708 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10045 6403 10103 6409
rect 8628 6344 8708 6372
rect 10060 6372 10088 6403
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 10284 6412 10517 6440
rect 10284 6400 10290 6412
rect 10505 6409 10517 6412
rect 10551 6409 10563 6443
rect 10505 6403 10563 6409
rect 12437 6443 12495 6449
rect 12437 6409 12449 6443
rect 12483 6440 12495 6443
rect 13630 6440 13636 6452
rect 12483 6412 13636 6440
rect 12483 6409 12495 6412
rect 12437 6403 12495 6409
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 10318 6372 10324 6384
rect 10060 6344 10324 6372
rect 8628 6332 8634 6344
rect 10318 6332 10324 6344
rect 10376 6372 10382 6384
rect 10376 6344 11192 6372
rect 10376 6332 10382 6344
rect 2406 6304 2412 6316
rect 2367 6276 2412 6304
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 3068 6304 3096 6332
rect 10965 6307 11023 6313
rect 3068 6276 3188 6304
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 2225 6239 2283 6245
rect 2225 6236 2237 6239
rect 1820 6208 2237 6236
rect 1820 6196 1826 6208
rect 2225 6205 2237 6208
rect 2271 6205 2283 6239
rect 2225 6199 2283 6205
rect 3053 6239 3111 6245
rect 3053 6205 3065 6239
rect 3099 6205 3111 6239
rect 3160 6236 3188 6276
rect 6656 6276 6960 6304
rect 3309 6239 3367 6245
rect 3309 6236 3321 6239
rect 3160 6208 3321 6236
rect 3053 6199 3111 6205
rect 3309 6205 3321 6208
rect 3355 6236 3367 6239
rect 4430 6236 4436 6248
rect 3355 6208 4436 6236
rect 3355 6205 3367 6208
rect 3309 6199 3367 6205
rect 2590 6128 2596 6180
rect 2648 6168 2654 6180
rect 3068 6168 3096 6199
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 4893 6239 4951 6245
rect 4893 6236 4905 6239
rect 4856 6208 4905 6236
rect 4856 6196 4862 6208
rect 4893 6205 4905 6208
rect 4939 6205 4951 6239
rect 4893 6199 4951 6205
rect 5718 6196 5724 6248
rect 5776 6236 5782 6248
rect 6656 6236 6684 6276
rect 6822 6236 6828 6248
rect 5776 6208 6684 6236
rect 6735 6208 6828 6236
rect 5776 6196 5782 6208
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 6932 6236 6960 6276
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 11054 6304 11060 6316
rect 11011 6276 11060 6304
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 11054 6264 11060 6276
rect 11112 6264 11118 6316
rect 11164 6313 11192 6344
rect 12158 6332 12164 6384
rect 12216 6372 12222 6384
rect 13262 6372 13268 6384
rect 12216 6344 13268 6372
rect 12216 6332 12222 6344
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 13449 6375 13507 6381
rect 13449 6341 13461 6375
rect 13495 6372 13507 6375
rect 14274 6372 14280 6384
rect 13495 6344 14280 6372
rect 13495 6341 13507 6344
rect 13449 6335 13507 6341
rect 14274 6332 14280 6344
rect 14332 6332 14338 6384
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6273 11207 6307
rect 11698 6304 11704 6316
rect 11659 6276 11704 6304
rect 11149 6267 11207 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 12342 6264 12348 6316
rect 12400 6304 12406 6316
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12400 6276 13001 6304
rect 12400 6264 12406 6276
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 13078 6264 13084 6316
rect 13136 6304 13142 6316
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 13136 6276 14197 6304
rect 13136 6264 13142 6276
rect 14185 6273 14197 6276
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 7081 6239 7139 6245
rect 7081 6236 7093 6239
rect 6932 6208 7093 6236
rect 7081 6205 7093 6208
rect 7127 6236 7139 6239
rect 7374 6236 7380 6248
rect 7127 6208 7380 6236
rect 7127 6205 7139 6208
rect 7081 6199 7139 6205
rect 7374 6196 7380 6208
rect 7432 6236 7438 6248
rect 7558 6236 7564 6248
rect 7432 6208 7564 6236
rect 7432 6196 7438 6208
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 7834 6236 7840 6248
rect 7708 6208 7840 6236
rect 7708 6196 7714 6208
rect 7834 6196 7840 6208
rect 7892 6236 7898 6248
rect 8665 6239 8723 6245
rect 8665 6236 8677 6239
rect 7892 6208 8677 6236
rect 7892 6196 7898 6208
rect 8665 6205 8677 6208
rect 8711 6205 8723 6239
rect 9398 6236 9404 6248
rect 8665 6199 8723 6205
rect 9232 6208 9404 6236
rect 4816 6168 4844 6196
rect 2648 6140 4844 6168
rect 5160 6171 5218 6177
rect 2648 6128 2654 6140
rect 5160 6137 5172 6171
rect 5206 6168 5218 6171
rect 6454 6168 6460 6180
rect 5206 6140 6460 6168
rect 5206 6137 5218 6140
rect 5160 6131 5218 6137
rect 6454 6128 6460 6140
rect 6512 6128 6518 6180
rect 6840 6168 6868 6196
rect 7668 6168 7696 6196
rect 6840 6140 7696 6168
rect 7742 6128 7748 6180
rect 7800 6168 7806 6180
rect 8910 6171 8968 6177
rect 8910 6168 8922 6171
rect 7800 6140 8922 6168
rect 7800 6128 7806 6140
rect 8910 6137 8922 6140
rect 8956 6137 8968 6171
rect 9232 6168 9260 6208
rect 9398 6196 9404 6208
rect 9456 6236 9462 6248
rect 9950 6236 9956 6248
rect 9456 6208 9956 6236
rect 9456 6196 9462 6208
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 10226 6196 10232 6248
rect 10284 6236 10290 6248
rect 12618 6236 12624 6248
rect 10284 6208 12624 6236
rect 10284 6196 10290 6208
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 12802 6236 12808 6248
rect 12763 6208 12808 6236
rect 12802 6196 12808 6208
rect 12860 6236 12866 6248
rect 13265 6239 13323 6245
rect 13265 6236 13277 6239
rect 12860 6208 13277 6236
rect 12860 6196 12866 6208
rect 13265 6205 13277 6208
rect 13311 6205 13323 6239
rect 13265 6199 13323 6205
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6236 14887 6239
rect 15286 6236 15292 6248
rect 14875 6208 15292 6236
rect 14875 6205 14887 6208
rect 14829 6199 14887 6205
rect 15286 6196 15292 6208
rect 15344 6196 15350 6248
rect 13078 6168 13084 6180
rect 8910 6131 8968 6137
rect 9140 6140 9260 6168
rect 9692 6140 13084 6168
rect 2317 6103 2375 6109
rect 2317 6069 2329 6103
rect 2363 6100 2375 6103
rect 4338 6100 4344 6112
rect 2363 6072 4344 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 4430 6060 4436 6112
rect 4488 6100 4494 6112
rect 5810 6100 5816 6112
rect 4488 6072 5816 6100
rect 4488 6060 4494 6072
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 6273 6103 6331 6109
rect 6273 6069 6285 6103
rect 6319 6100 6331 6103
rect 6362 6100 6368 6112
rect 6319 6072 6368 6100
rect 6319 6069 6331 6072
rect 6273 6063 6331 6069
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 7006 6060 7012 6112
rect 7064 6100 7070 6112
rect 8478 6100 8484 6112
rect 7064 6072 8484 6100
rect 7064 6060 7070 6072
rect 8478 6060 8484 6072
rect 8536 6060 8542 6112
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 9140 6100 9168 6140
rect 9692 6112 9720 6140
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 13906 6128 13912 6180
rect 13964 6168 13970 6180
rect 14093 6171 14151 6177
rect 14093 6168 14105 6171
rect 13964 6140 14105 6168
rect 13964 6128 13970 6140
rect 14093 6137 14105 6140
rect 14139 6137 14151 6171
rect 14093 6131 14151 6137
rect 8628 6072 9168 6100
rect 8628 6060 8634 6072
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 9674 6100 9680 6112
rect 9272 6072 9680 6100
rect 9272 6060 9278 6072
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 10873 6103 10931 6109
rect 10873 6069 10885 6103
rect 10919 6100 10931 6103
rect 12618 6100 12624 6112
rect 10919 6072 12624 6100
rect 10919 6069 10931 6072
rect 10873 6063 10931 6069
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 12897 6103 12955 6109
rect 12897 6069 12909 6103
rect 12943 6100 12955 6103
rect 13449 6103 13507 6109
rect 13449 6100 13461 6103
rect 12943 6072 13461 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 13449 6069 13461 6072
rect 13495 6069 13507 6103
rect 13449 6063 13507 6069
rect 13538 6060 13544 6112
rect 13596 6100 13602 6112
rect 13633 6103 13691 6109
rect 13633 6100 13645 6103
rect 13596 6072 13645 6100
rect 13596 6060 13602 6072
rect 13633 6069 13645 6072
rect 13679 6069 13691 6103
rect 13633 6063 13691 6069
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 14001 6103 14059 6109
rect 14001 6100 14013 6103
rect 13780 6072 14013 6100
rect 13780 6060 13786 6072
rect 14001 6069 14013 6072
rect 14047 6069 14059 6103
rect 14001 6063 14059 6069
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 14826 6100 14832 6112
rect 14700 6072 14832 6100
rect 14700 6060 14706 6072
rect 14826 6060 14832 6072
rect 14884 6060 14890 6112
rect 15010 6100 15016 6112
rect 14971 6072 15016 6100
rect 15010 6060 15016 6072
rect 15068 6060 15074 6112
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 1394 5896 1400 5908
rect 1355 5868 1400 5896
rect 1394 5856 1400 5868
rect 1452 5856 1458 5908
rect 3145 5899 3203 5905
rect 3145 5865 3157 5899
rect 3191 5896 3203 5899
rect 4430 5896 4436 5908
rect 3191 5868 4436 5896
rect 3191 5865 3203 5868
rect 3145 5859 3203 5865
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 4890 5896 4896 5908
rect 4851 5868 4896 5896
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 4982 5856 4988 5908
rect 5040 5896 5046 5908
rect 9677 5899 9735 5905
rect 9677 5896 9689 5899
rect 5040 5868 9689 5896
rect 5040 5856 5046 5868
rect 9677 5865 9689 5868
rect 9723 5865 9735 5899
rect 9677 5859 9735 5865
rect 11241 5899 11299 5905
rect 11241 5865 11253 5899
rect 11287 5896 11299 5899
rect 11330 5896 11336 5908
rect 11287 5868 11336 5896
rect 11287 5865 11299 5868
rect 11241 5859 11299 5865
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 14550 5896 14556 5908
rect 12676 5868 14556 5896
rect 12676 5856 12682 5868
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 14642 5856 14648 5908
rect 14700 5896 14706 5908
rect 14700 5868 14745 5896
rect 14700 5856 14706 5868
rect 1302 5788 1308 5840
rect 1360 5828 1366 5840
rect 1765 5831 1823 5837
rect 1765 5828 1777 5831
rect 1360 5800 1777 5828
rect 1360 5788 1366 5800
rect 1765 5797 1777 5800
rect 1811 5797 1823 5831
rect 1765 5791 1823 5797
rect 2038 5788 2044 5840
rect 2096 5828 2102 5840
rect 2501 5831 2559 5837
rect 2096 5800 2268 5828
rect 2096 5788 2102 5800
rect 2240 5769 2268 5800
rect 2501 5797 2513 5831
rect 2547 5828 2559 5831
rect 2774 5828 2780 5840
rect 2547 5800 2780 5828
rect 2547 5797 2559 5800
rect 2501 5791 2559 5797
rect 2774 5788 2780 5800
rect 2832 5788 2838 5840
rect 5442 5828 5448 5840
rect 2884 5800 5448 5828
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5729 2283 5763
rect 2225 5723 2283 5729
rect 2406 5720 2412 5772
rect 2464 5760 2470 5772
rect 2884 5760 2912 5800
rect 5442 5788 5448 5800
rect 5500 5788 5506 5840
rect 5552 5800 6224 5828
rect 2464 5732 2912 5760
rect 3237 5763 3295 5769
rect 2464 5720 2470 5732
rect 3237 5729 3249 5763
rect 3283 5760 3295 5763
rect 5552 5760 5580 5800
rect 5977 5763 6035 5769
rect 5977 5760 5989 5763
rect 3283 5732 5580 5760
rect 5644 5732 5989 5760
rect 3283 5729 3295 5732
rect 3237 5723 3295 5729
rect 5644 5704 5672 5732
rect 5977 5729 5989 5732
rect 6023 5729 6035 5763
rect 6196 5760 6224 5800
rect 6270 5788 6276 5840
rect 6328 5828 6334 5840
rect 7920 5831 7978 5837
rect 6328 5800 7880 5828
rect 6328 5788 6334 5800
rect 7742 5760 7748 5772
rect 6196 5732 7748 5760
rect 5977 5723 6035 5729
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 7852 5760 7880 5800
rect 7920 5797 7932 5831
rect 7966 5828 7978 5831
rect 9766 5828 9772 5840
rect 7966 5800 9772 5828
rect 7966 5797 7978 5800
rect 7920 5791 7978 5797
rect 9766 5788 9772 5800
rect 9824 5788 9830 5840
rect 10045 5831 10103 5837
rect 10045 5797 10057 5831
rect 10091 5828 10103 5831
rect 10686 5828 10692 5840
rect 10091 5800 10692 5828
rect 10091 5797 10103 5800
rect 10045 5791 10103 5797
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 11974 5828 11980 5840
rect 11348 5800 11980 5828
rect 9214 5760 9220 5772
rect 7852 5732 9220 5760
rect 9214 5720 9220 5732
rect 9272 5720 9278 5772
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 11348 5769 11376 5800
rect 11974 5788 11980 5800
rect 12032 5788 12038 5840
rect 12437 5831 12495 5837
rect 12437 5797 12449 5831
rect 12483 5828 12495 5831
rect 13725 5831 13783 5837
rect 12483 5800 12756 5828
rect 12483 5797 12495 5800
rect 12437 5791 12495 5797
rect 10137 5763 10195 5769
rect 10137 5760 10149 5763
rect 9640 5732 10149 5760
rect 9640 5720 9646 5732
rect 10137 5729 10149 5732
rect 10183 5760 10195 5763
rect 11333 5763 11391 5769
rect 10183 5732 11284 5760
rect 10183 5729 10195 5732
rect 10137 5723 10195 5729
rect 1762 5652 1768 5704
rect 1820 5692 1826 5704
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1820 5664 1869 5692
rect 1820 5652 1826 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 4614 5692 4620 5704
rect 3467 5664 4620 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 2056 5624 2084 5655
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4982 5692 4988 5704
rect 4943 5664 4988 5692
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5692 5227 5695
rect 5442 5692 5448 5704
rect 5215 5664 5448 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 5626 5652 5632 5704
rect 5684 5652 5690 5704
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 2222 5624 2228 5636
rect 2056 5596 2228 5624
rect 2222 5584 2228 5596
rect 2280 5584 2286 5636
rect 4525 5627 4583 5633
rect 4525 5593 4537 5627
rect 4571 5624 4583 5627
rect 5350 5624 5356 5636
rect 4571 5596 5356 5624
rect 4571 5593 4583 5596
rect 4525 5587 4583 5593
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5556 2835 5559
rect 4430 5556 4436 5568
rect 2823 5528 4436 5556
rect 2823 5525 2835 5528
rect 2777 5519 2835 5525
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 5736 5556 5764 5655
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 7650 5692 7656 5704
rect 7432 5664 7656 5692
rect 7432 5652 7438 5664
rect 7650 5652 7656 5664
rect 7708 5652 7714 5704
rect 10318 5692 10324 5704
rect 8687 5664 8964 5692
rect 10279 5664 10324 5692
rect 6730 5584 6736 5636
rect 6788 5624 6794 5636
rect 8687 5624 8715 5664
rect 6788 5596 7227 5624
rect 6788 5584 6794 5596
rect 5994 5556 6000 5568
rect 4948 5528 6000 5556
rect 4948 5516 4954 5528
rect 5994 5516 6000 5528
rect 6052 5516 6058 5568
rect 6454 5516 6460 5568
rect 6512 5556 6518 5568
rect 7006 5556 7012 5568
rect 6512 5528 7012 5556
rect 6512 5516 6518 5528
rect 7006 5516 7012 5528
rect 7064 5556 7070 5568
rect 7101 5559 7159 5565
rect 7101 5556 7113 5559
rect 7064 5528 7113 5556
rect 7064 5516 7070 5528
rect 7101 5525 7113 5528
rect 7147 5525 7159 5559
rect 7199 5556 7227 5596
rect 8588 5596 8715 5624
rect 8936 5624 8964 5664
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 10873 5627 10931 5633
rect 10873 5624 10885 5627
rect 8936 5596 10885 5624
rect 8588 5556 8616 5596
rect 10873 5593 10885 5596
rect 10919 5593 10931 5627
rect 11256 5624 11284 5732
rect 11333 5729 11345 5763
rect 11379 5729 11391 5763
rect 11333 5723 11391 5729
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 11756 5732 12296 5760
rect 11756 5720 11762 5732
rect 11514 5652 11520 5704
rect 11572 5692 11578 5704
rect 11572 5664 11617 5692
rect 11572 5652 11578 5664
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 12158 5692 12164 5704
rect 12032 5664 12164 5692
rect 12032 5652 12038 5664
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 12268 5692 12296 5732
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 12728 5760 12756 5800
rect 13725 5797 13737 5831
rect 13771 5828 13783 5831
rect 14918 5828 14924 5840
rect 13771 5800 14924 5828
rect 13771 5797 13783 5800
rect 13725 5791 13783 5797
rect 14918 5788 14924 5800
rect 14976 5788 14982 5840
rect 12986 5760 12992 5772
rect 12400 5732 12664 5760
rect 12728 5732 12992 5760
rect 12400 5720 12406 5732
rect 12636 5701 12664 5732
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 13633 5763 13691 5769
rect 13633 5760 13645 5763
rect 13096 5732 13645 5760
rect 12529 5695 12587 5701
rect 12268 5664 12480 5692
rect 12342 5624 12348 5636
rect 11256 5596 12348 5624
rect 10873 5587 10931 5593
rect 12342 5584 12348 5596
rect 12400 5584 12406 5636
rect 9030 5556 9036 5568
rect 7199 5528 8616 5556
rect 8943 5528 9036 5556
rect 7101 5519 7159 5525
rect 9030 5516 9036 5528
rect 9088 5556 9094 5568
rect 9582 5556 9588 5568
rect 9088 5528 9588 5556
rect 9088 5516 9094 5528
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 11238 5516 11244 5568
rect 11296 5556 11302 5568
rect 11514 5556 11520 5568
rect 11296 5528 11520 5556
rect 11296 5516 11302 5528
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 11698 5516 11704 5568
rect 11756 5556 11762 5568
rect 12069 5559 12127 5565
rect 12069 5556 12081 5559
rect 11756 5528 12081 5556
rect 11756 5516 11762 5528
rect 12069 5525 12081 5528
rect 12115 5525 12127 5559
rect 12452 5556 12480 5664
rect 12529 5661 12541 5695
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5661 12679 5695
rect 13096 5692 13124 5732
rect 13633 5729 13645 5732
rect 13679 5729 13691 5763
rect 13633 5723 13691 5729
rect 14182 5720 14188 5772
rect 14240 5760 14246 5772
rect 14461 5763 14519 5769
rect 14461 5760 14473 5763
rect 14240 5732 14473 5760
rect 14240 5720 14246 5732
rect 14461 5729 14473 5732
rect 14507 5729 14519 5763
rect 14461 5723 14519 5729
rect 12621 5655 12679 5661
rect 12912 5664 13124 5692
rect 12544 5624 12572 5655
rect 12710 5624 12716 5636
rect 12544 5596 12716 5624
rect 12710 5584 12716 5596
rect 12768 5584 12774 5636
rect 12912 5556 12940 5664
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 13817 5695 13875 5701
rect 13817 5692 13829 5695
rect 13320 5664 13829 5692
rect 13320 5652 13326 5664
rect 13817 5661 13829 5664
rect 13863 5661 13875 5695
rect 13817 5655 13875 5661
rect 13078 5584 13084 5636
rect 13136 5624 13142 5636
rect 13538 5624 13544 5636
rect 13136 5596 13544 5624
rect 13136 5584 13142 5596
rect 13538 5584 13544 5596
rect 13596 5584 13602 5636
rect 12452 5528 12940 5556
rect 12069 5519 12127 5525
rect 12986 5516 12992 5568
rect 13044 5556 13050 5568
rect 13265 5559 13323 5565
rect 13265 5556 13277 5559
rect 13044 5528 13277 5556
rect 13044 5516 13050 5528
rect 13265 5525 13277 5528
rect 13311 5525 13323 5559
rect 13265 5519 13323 5525
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 4798 5352 4804 5364
rect 1872 5324 4804 5352
rect 1872 5225 1900 5324
rect 4798 5312 4804 5324
rect 4856 5352 4862 5364
rect 4856 5324 6040 5352
rect 4856 5312 4862 5324
rect 3326 5244 3332 5296
rect 3384 5284 3390 5296
rect 3513 5287 3571 5293
rect 3513 5284 3525 5287
rect 3384 5256 3525 5284
rect 3384 5244 3390 5256
rect 3513 5253 3525 5256
rect 3559 5253 3571 5287
rect 3513 5247 3571 5253
rect 3602 5244 3608 5296
rect 3660 5284 3666 5296
rect 6012 5284 6040 5324
rect 6086 5312 6092 5364
rect 6144 5352 6150 5364
rect 6273 5355 6331 5361
rect 6273 5352 6285 5355
rect 6144 5324 6285 5352
rect 6144 5312 6150 5324
rect 6273 5321 6285 5324
rect 6319 5321 6331 5355
rect 7558 5352 7564 5364
rect 6273 5315 6331 5321
rect 7392 5324 7564 5352
rect 7392 5284 7420 5324
rect 7558 5312 7564 5324
rect 7616 5312 7622 5364
rect 7650 5312 7656 5364
rect 7708 5352 7714 5364
rect 9214 5352 9220 5364
rect 7708 5324 8524 5352
rect 9175 5324 9220 5352
rect 7708 5312 7714 5324
rect 3660 5256 4936 5284
rect 6012 5256 7420 5284
rect 3660 5244 3666 5256
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 1670 5108 1676 5160
rect 1728 5148 1734 5160
rect 1964 5148 1992 5179
rect 2866 5176 2872 5228
rect 2924 5216 2930 5228
rect 2961 5219 3019 5225
rect 2961 5216 2973 5219
rect 2924 5188 2973 5216
rect 2924 5176 2930 5188
rect 2961 5185 2973 5188
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5216 3203 5219
rect 4062 5216 4068 5228
rect 3191 5188 4068 5216
rect 3191 5185 3203 5188
rect 3145 5179 3203 5185
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4614 5216 4620 5228
rect 4387 5188 4620 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 4908 5216 4936 5256
rect 7374 5216 7380 5228
rect 4908 5188 5019 5216
rect 7335 5188 7380 5216
rect 1728 5120 1992 5148
rect 3329 5151 3387 5157
rect 1728 5108 1734 5120
rect 3329 5117 3341 5151
rect 3375 5148 3387 5151
rect 3510 5148 3516 5160
rect 3375 5120 3516 5148
rect 3375 5117 3387 5120
rect 3329 5111 3387 5117
rect 3510 5108 3516 5120
rect 3568 5108 3574 5160
rect 4522 5148 4528 5160
rect 3712 5120 4528 5148
rect 1765 5083 1823 5089
rect 1765 5049 1777 5083
rect 1811 5080 1823 5083
rect 2774 5080 2780 5092
rect 1811 5052 2780 5080
rect 1811 5049 1823 5052
rect 1765 5043 1823 5049
rect 2774 5040 2780 5052
rect 2832 5040 2838 5092
rect 2869 5083 2927 5089
rect 2869 5049 2881 5083
rect 2915 5080 2927 5083
rect 3712 5080 3740 5120
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 4890 5148 4896 5160
rect 4851 5120 4896 5148
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 4991 5148 5019 5188
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 8496 5216 8524 5324
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 9674 5352 9680 5364
rect 9324 5324 9680 5352
rect 8757 5287 8815 5293
rect 8757 5253 8769 5287
rect 8803 5284 8815 5287
rect 9324 5284 9352 5324
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 10413 5355 10471 5361
rect 10413 5321 10425 5355
rect 10459 5352 10471 5355
rect 10502 5352 10508 5364
rect 10459 5324 10508 5352
rect 10459 5321 10471 5324
rect 10413 5315 10471 5321
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 11241 5355 11299 5361
rect 11241 5321 11253 5355
rect 11287 5352 11299 5355
rect 12434 5352 12440 5364
rect 11287 5324 12440 5352
rect 11287 5321 11299 5324
rect 11241 5315 11299 5321
rect 12434 5312 12440 5324
rect 12492 5312 12498 5364
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 13814 5352 13820 5364
rect 12584 5324 13820 5352
rect 12584 5312 12590 5324
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 14090 5312 14096 5364
rect 14148 5352 14154 5364
rect 14550 5352 14556 5364
rect 14148 5324 14556 5352
rect 14148 5312 14154 5324
rect 14550 5312 14556 5324
rect 14608 5312 14614 5364
rect 12158 5284 12164 5296
rect 8803 5256 9352 5284
rect 9416 5256 12164 5284
rect 8803 5253 8815 5256
rect 8757 5247 8815 5253
rect 9416 5216 9444 5256
rect 8496 5188 9444 5216
rect 9490 5176 9496 5228
rect 9548 5216 9554 5228
rect 9769 5219 9827 5225
rect 9769 5216 9781 5219
rect 9548 5188 9781 5216
rect 9548 5176 9554 5188
rect 9769 5185 9781 5188
rect 9815 5185 9827 5219
rect 9769 5179 9827 5185
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10980 5225 11008 5256
rect 12158 5244 12164 5256
rect 12216 5244 12222 5296
rect 12250 5244 12256 5296
rect 12308 5284 12314 5296
rect 12308 5256 13032 5284
rect 12308 5244 12314 5256
rect 10965 5219 11023 5225
rect 10192 5188 10916 5216
rect 10192 5176 10198 5188
rect 7926 5148 7932 5160
rect 4991 5120 7932 5148
rect 7926 5108 7932 5120
rect 7984 5148 7990 5160
rect 8570 5148 8576 5160
rect 7984 5120 8576 5148
rect 7984 5108 7990 5120
rect 8570 5108 8576 5120
rect 8628 5148 8634 5160
rect 8628 5120 9720 5148
rect 8628 5108 8634 5120
rect 2915 5052 3740 5080
rect 4065 5083 4123 5089
rect 2915 5049 2927 5052
rect 2869 5043 2927 5049
rect 4065 5049 4077 5083
rect 4111 5080 4123 5083
rect 4798 5080 4804 5092
rect 4111 5052 4804 5080
rect 4111 5049 4123 5052
rect 4065 5043 4123 5049
rect 4798 5040 4804 5052
rect 4856 5040 4862 5092
rect 5166 5089 5172 5092
rect 5160 5080 5172 5089
rect 5127 5052 5172 5080
rect 5160 5043 5172 5052
rect 5224 5080 5230 5092
rect 5810 5080 5816 5092
rect 5224 5052 5816 5080
rect 5166 5040 5172 5043
rect 5224 5040 5230 5052
rect 5810 5040 5816 5052
rect 5868 5040 5874 5092
rect 6454 5040 6460 5092
rect 6512 5080 6518 5092
rect 7006 5080 7012 5092
rect 6512 5052 7012 5080
rect 6512 5040 6518 5052
rect 7006 5040 7012 5052
rect 7064 5040 7070 5092
rect 7190 5040 7196 5092
rect 7248 5080 7254 5092
rect 7374 5080 7380 5092
rect 7248 5052 7380 5080
rect 7248 5040 7254 5052
rect 7374 5040 7380 5052
rect 7432 5040 7438 5092
rect 7644 5083 7702 5089
rect 7644 5049 7656 5083
rect 7690 5080 7702 5083
rect 8294 5080 8300 5092
rect 7690 5052 8300 5080
rect 7690 5049 7702 5052
rect 7644 5043 7702 5049
rect 8294 5040 8300 5052
rect 8352 5040 8358 5092
rect 9030 5080 9036 5092
rect 8687 5052 9036 5080
rect 1394 5012 1400 5024
rect 1355 4984 1400 5012
rect 1394 4972 1400 4984
rect 1452 4972 1458 5024
rect 2501 5015 2559 5021
rect 2501 4981 2513 5015
rect 2547 5012 2559 5015
rect 3234 5012 3240 5024
rect 2547 4984 3240 5012
rect 2547 4981 2559 4984
rect 2501 4975 2559 4981
rect 3234 4972 3240 4984
rect 3292 4972 3298 5024
rect 3694 5012 3700 5024
rect 3655 4984 3700 5012
rect 3694 4972 3700 4984
rect 3752 4972 3758 5024
rect 4157 5015 4215 5021
rect 4157 4981 4169 5015
rect 4203 5012 4215 5015
rect 5534 5012 5540 5024
rect 4203 4984 5540 5012
rect 4203 4981 4215 4984
rect 4157 4975 4215 4981
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 5626 4972 5632 5024
rect 5684 5012 5690 5024
rect 8687 5012 8715 5052
rect 9030 5040 9036 5052
rect 9088 5040 9094 5092
rect 9585 5083 9643 5089
rect 9585 5080 9597 5083
rect 9416 5052 9597 5080
rect 5684 4984 8715 5012
rect 5684 4972 5690 4984
rect 8754 4972 8760 5024
rect 8812 5012 8818 5024
rect 9416 5012 9444 5052
rect 9585 5049 9597 5052
rect 9631 5049 9643 5083
rect 9692 5080 9720 5120
rect 10410 5108 10416 5160
rect 10468 5148 10474 5160
rect 10781 5151 10839 5157
rect 10781 5148 10793 5151
rect 10468 5120 10793 5148
rect 10468 5108 10474 5120
rect 10781 5117 10793 5120
rect 10827 5117 10839 5151
rect 10888 5148 10916 5188
rect 10965 5185 10977 5219
rect 11011 5216 11023 5219
rect 11885 5219 11943 5225
rect 11011 5188 11045 5216
rect 11440 5188 11816 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 11440 5148 11468 5188
rect 10888 5120 11468 5148
rect 10781 5111 10839 5117
rect 11514 5108 11520 5160
rect 11572 5148 11578 5160
rect 11701 5151 11759 5157
rect 11701 5148 11713 5151
rect 11572 5120 11713 5148
rect 11572 5108 11578 5120
rect 11701 5117 11713 5120
rect 11747 5117 11759 5151
rect 11788 5148 11816 5188
rect 11885 5185 11897 5219
rect 11931 5216 11943 5219
rect 12618 5216 12624 5228
rect 11931 5188 12624 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 13004 5225 13032 5256
rect 13998 5244 14004 5296
rect 14056 5284 14062 5296
rect 14056 5256 14872 5284
rect 14056 5244 14062 5256
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 13354 5176 13360 5228
rect 13412 5216 13418 5228
rect 13906 5216 13912 5228
rect 13412 5188 13912 5216
rect 13412 5176 13418 5188
rect 13906 5176 13912 5188
rect 13964 5176 13970 5228
rect 14090 5176 14096 5228
rect 14148 5216 14154 5228
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 14148 5188 14197 5216
rect 14148 5176 14154 5188
rect 14185 5185 14197 5188
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 12250 5148 12256 5160
rect 11788 5120 12256 5148
rect 11701 5111 11759 5117
rect 12250 5108 12256 5120
rect 12308 5108 12314 5160
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 13078 5148 13084 5160
rect 12943 5120 13084 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 14844 5157 14872 5256
rect 14001 5151 14059 5157
rect 14001 5148 14013 5151
rect 13872 5120 14013 5148
rect 13872 5108 13878 5120
rect 14001 5117 14013 5120
rect 14047 5117 14059 5151
rect 14001 5111 14059 5117
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5117 14887 5151
rect 14829 5111 14887 5117
rect 10873 5083 10931 5089
rect 10873 5080 10885 5083
rect 9692 5052 10885 5080
rect 9585 5043 9643 5049
rect 10873 5049 10885 5052
rect 10919 5049 10931 5083
rect 10873 5043 10931 5049
rect 9674 5012 9680 5024
rect 8812 4984 9444 5012
rect 9635 4984 9680 5012
rect 8812 4972 8818 4984
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 10888 5012 10916 5043
rect 10962 5040 10968 5092
rect 11020 5080 11026 5092
rect 12805 5083 12863 5089
rect 12805 5080 12817 5083
rect 11020 5052 12817 5080
rect 11020 5040 11026 5052
rect 12805 5049 12817 5052
rect 12851 5049 12863 5083
rect 13906 5080 13912 5092
rect 12805 5043 12863 5049
rect 13280 5052 13912 5080
rect 11514 5012 11520 5024
rect 10888 4984 11520 5012
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 11609 5015 11667 5021
rect 11609 4981 11621 5015
rect 11655 5012 11667 5015
rect 11698 5012 11704 5024
rect 11655 4984 11704 5012
rect 11655 4981 11667 4984
rect 11609 4975 11667 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 12437 5015 12495 5021
rect 12437 4981 12449 5015
rect 12483 5012 12495 5015
rect 13280 5012 13308 5052
rect 13906 5040 13912 5052
rect 13964 5040 13970 5092
rect 13630 5012 13636 5024
rect 12483 4984 13308 5012
rect 13591 4984 13636 5012
rect 12483 4981 12495 4984
rect 12437 4975 12495 4981
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 13814 4972 13820 5024
rect 13872 5012 13878 5024
rect 14093 5015 14151 5021
rect 14093 5012 14105 5015
rect 13872 4984 14105 5012
rect 13872 4972 13878 4984
rect 14093 4981 14105 4984
rect 14139 4981 14151 5015
rect 14093 4975 14151 4981
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 15013 5015 15071 5021
rect 15013 5012 15025 5015
rect 14240 4984 15025 5012
rect 14240 4972 14246 4984
rect 15013 4981 15025 4984
rect 15059 4981 15071 5015
rect 15013 4975 15071 4981
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 2958 4808 2964 4820
rect 2823 4780 2964 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 3237 4811 3295 4817
rect 3237 4777 3249 4811
rect 3283 4808 3295 4811
rect 3602 4808 3608 4820
rect 3283 4780 3608 4808
rect 3283 4777 3295 4780
rect 3237 4771 3295 4777
rect 3602 4768 3608 4780
rect 3660 4768 3666 4820
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 4525 4811 4583 4817
rect 4525 4808 4537 4811
rect 3752 4780 4537 4808
rect 3752 4768 3758 4780
rect 4525 4777 4537 4780
rect 4571 4777 4583 4811
rect 4525 4771 4583 4777
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 5040 4780 5273 4808
rect 5040 4768 5046 4780
rect 5261 4777 5273 4780
rect 5307 4777 5319 4811
rect 5261 4771 5319 4777
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 5626 4808 5632 4820
rect 5408 4780 5632 4808
rect 5408 4768 5414 4780
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 8297 4811 8355 4817
rect 8297 4808 8309 4811
rect 5736 4780 8309 4808
rect 1670 4749 1676 4752
rect 1664 4740 1676 4749
rect 1631 4712 1676 4740
rect 1664 4703 1676 4712
rect 1670 4700 1676 4703
rect 1728 4700 1734 4752
rect 4430 4740 4436 4752
rect 4391 4712 4436 4740
rect 4430 4700 4436 4712
rect 4488 4700 4494 4752
rect 4798 4700 4804 4752
rect 4856 4740 4862 4752
rect 5736 4740 5764 4780
rect 8297 4777 8309 4780
rect 8343 4777 8355 4811
rect 8297 4771 8355 4777
rect 8386 4768 8392 4820
rect 8444 4808 8450 4820
rect 8444 4780 8524 4808
rect 8444 4768 8450 4780
rect 6730 4749 6736 4752
rect 4856 4712 5764 4740
rect 4856 4700 4862 4712
rect 6724 4703 6736 4749
rect 6788 4740 6794 4752
rect 6788 4712 6824 4740
rect 6730 4700 6736 4703
rect 6788 4700 6794 4712
rect 5350 4672 5356 4684
rect 3528 4644 5356 4672
rect 3326 4604 3332 4616
rect 3239 4576 3332 4604
rect 3326 4564 3332 4576
rect 3384 4604 3390 4616
rect 3528 4613 3556 4644
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 5626 4632 5632 4684
rect 5684 4672 5690 4684
rect 5684 4644 5729 4672
rect 5684 4632 5690 4644
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 5868 4644 5948 4672
rect 5868 4632 5874 4644
rect 3513 4607 3571 4613
rect 3384 4576 3464 4604
rect 3384 4564 3390 4576
rect 2866 4536 2872 4548
rect 2827 4508 2872 4536
rect 2866 4496 2872 4508
rect 2924 4496 2930 4548
rect 3436 4536 3464 4576
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 3786 4564 3792 4616
rect 3844 4604 3850 4616
rect 5920 4613 5948 4644
rect 6270 4632 6276 4684
rect 6328 4672 6334 4684
rect 6457 4675 6515 4681
rect 6457 4672 6469 4675
rect 6328 4644 6469 4672
rect 6328 4632 6334 4644
rect 6457 4641 6469 4644
rect 6503 4672 6515 4675
rect 7006 4672 7012 4684
rect 6503 4644 7012 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 7006 4632 7012 4644
rect 7064 4632 7070 4684
rect 7834 4632 7840 4684
rect 7892 4672 7898 4684
rect 8294 4672 8300 4684
rect 7892 4644 8300 4672
rect 7892 4632 7898 4644
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8496 4672 8524 4780
rect 8570 4768 8576 4820
rect 8628 4808 8634 4820
rect 8757 4811 8815 4817
rect 8757 4808 8769 4811
rect 8628 4780 8769 4808
rect 8628 4768 8634 4780
rect 8757 4777 8769 4780
rect 8803 4777 8815 4811
rect 8757 4771 8815 4777
rect 9122 4768 9128 4820
rect 9180 4808 9186 4820
rect 9677 4811 9735 4817
rect 9677 4808 9689 4811
rect 9180 4780 9689 4808
rect 9180 4768 9186 4780
rect 9677 4777 9689 4780
rect 9723 4777 9735 4811
rect 10226 4808 10232 4820
rect 9677 4771 9735 4777
rect 9876 4780 10232 4808
rect 8665 4743 8723 4749
rect 8665 4709 8677 4743
rect 8711 4740 8723 4743
rect 9030 4740 9036 4752
rect 8711 4712 9036 4740
rect 8711 4709 8723 4712
rect 8665 4703 8723 4709
rect 9030 4700 9036 4712
rect 9088 4700 9094 4752
rect 8496 4644 8892 4672
rect 4617 4607 4675 4613
rect 4617 4604 4629 4607
rect 3844 4576 4629 4604
rect 3844 4564 3850 4576
rect 4617 4573 4629 4576
rect 4663 4573 4675 4607
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 4617 4567 4675 4573
rect 5552 4576 5733 4604
rect 5350 4536 5356 4548
rect 3436 4508 5356 4536
rect 5350 4496 5356 4508
rect 5408 4496 5414 4548
rect 3786 4428 3792 4480
rect 3844 4468 3850 4480
rect 4065 4471 4123 4477
rect 4065 4468 4077 4471
rect 3844 4440 4077 4468
rect 3844 4428 3850 4440
rect 4065 4437 4077 4440
rect 4111 4437 4123 4471
rect 5552 4468 5580 4576
rect 5721 4573 5733 4576
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 7558 4564 7564 4616
rect 7616 4604 7622 4616
rect 8754 4604 8760 4616
rect 7616 4576 8760 4604
rect 7616 4564 7622 4576
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 7392 4508 7963 4536
rect 5718 4468 5724 4480
rect 5552 4440 5724 4468
rect 4065 4431 4123 4437
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 7392 4468 7420 4508
rect 7834 4468 7840 4480
rect 5868 4440 7420 4468
rect 7795 4440 7840 4468
rect 5868 4428 5874 4440
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 7935 4468 7963 4508
rect 8018 4496 8024 4548
rect 8076 4536 8082 4548
rect 8662 4536 8668 4548
rect 8076 4508 8668 4536
rect 8076 4496 8082 4508
rect 8662 4496 8668 4508
rect 8720 4496 8726 4548
rect 8864 4536 8892 4644
rect 9214 4632 9220 4684
rect 9272 4672 9278 4684
rect 9876 4672 9904 4780
rect 10226 4768 10232 4780
rect 10284 4768 10290 4820
rect 11333 4811 11391 4817
rect 11333 4777 11345 4811
rect 11379 4808 11391 4811
rect 11885 4811 11943 4817
rect 11379 4780 11652 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 9950 4700 9956 4752
rect 10008 4740 10014 4752
rect 10594 4740 10600 4752
rect 10008 4712 10600 4740
rect 10008 4700 10014 4712
rect 10594 4700 10600 4712
rect 10652 4700 10658 4752
rect 11238 4700 11244 4752
rect 11296 4740 11302 4752
rect 11624 4740 11652 4780
rect 11885 4777 11897 4811
rect 11931 4808 11943 4811
rect 11974 4808 11980 4820
rect 11931 4780 11980 4808
rect 11931 4777 11943 4780
rect 11885 4771 11943 4777
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 12250 4768 12256 4820
rect 12308 4808 12314 4820
rect 12618 4808 12624 4820
rect 12308 4780 12624 4808
rect 12308 4768 12314 4780
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 12894 4768 12900 4820
rect 12952 4808 12958 4820
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 12952 4780 13645 4808
rect 12952 4768 12958 4780
rect 13633 4777 13645 4780
rect 13679 4777 13691 4811
rect 13633 4771 13691 4777
rect 12342 4740 12348 4752
rect 11296 4712 11341 4740
rect 11624 4712 12348 4740
rect 11296 4700 11302 4712
rect 12342 4700 12348 4712
rect 12400 4700 12406 4752
rect 12437 4743 12495 4749
rect 12437 4709 12449 4743
rect 12483 4709 12495 4743
rect 12437 4703 12495 4709
rect 9272 4644 9904 4672
rect 10045 4675 10103 4681
rect 9272 4632 9278 4644
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 11698 4672 11704 4684
rect 10091 4644 11192 4672
rect 11659 4644 11704 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 11164 4616 11192 4644
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 12452 4616 12480 4703
rect 13446 4700 13452 4752
rect 13504 4740 13510 4752
rect 13725 4743 13783 4749
rect 13725 4740 13737 4743
rect 13504 4712 13737 4740
rect 13504 4700 13510 4712
rect 13725 4709 13737 4712
rect 13771 4709 13783 4743
rect 13725 4703 13783 4709
rect 14090 4672 14096 4684
rect 12636 4644 14096 4672
rect 12636 4616 12664 4644
rect 14090 4632 14096 4644
rect 14148 4632 14154 4684
rect 14458 4672 14464 4684
rect 14419 4644 14464 4672
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4604 8999 4607
rect 9490 4604 9496 4616
rect 8987 4576 9496 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 10134 4604 10140 4616
rect 10095 4576 10140 4604
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 10244 4536 10272 4567
rect 11146 4564 11152 4616
rect 11204 4564 11210 4616
rect 11517 4607 11575 4613
rect 11517 4573 11529 4607
rect 11563 4604 11575 4607
rect 12066 4604 12072 4616
rect 11563 4576 12072 4604
rect 11563 4573 11575 4576
rect 11517 4567 11575 4573
rect 10870 4536 10876 4548
rect 8864 4508 10272 4536
rect 10336 4508 10640 4536
rect 10831 4508 10876 4536
rect 10336 4468 10364 4508
rect 7935 4440 10364 4468
rect 10612 4468 10640 4508
rect 10870 4496 10876 4508
rect 10928 4496 10934 4548
rect 10962 4496 10968 4548
rect 11020 4536 11026 4548
rect 11532 4536 11560 4567
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 12434 4564 12440 4616
rect 12492 4564 12498 4616
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4573 12587 4607
rect 12529 4567 12587 4573
rect 11020 4508 11560 4536
rect 11020 4496 11026 4508
rect 11882 4496 11888 4548
rect 11940 4536 11946 4548
rect 12544 4536 12572 4567
rect 12618 4564 12624 4616
rect 12676 4604 12682 4616
rect 12676 4576 12721 4604
rect 12676 4564 12682 4576
rect 12894 4564 12900 4616
rect 12952 4604 12958 4616
rect 13817 4607 13875 4613
rect 13817 4604 13829 4607
rect 12952 4576 13829 4604
rect 12952 4564 12958 4576
rect 13817 4573 13829 4576
rect 13863 4573 13875 4607
rect 13817 4567 13875 4573
rect 11940 4508 12572 4536
rect 11940 4496 11946 4508
rect 12069 4471 12127 4477
rect 12069 4468 12081 4471
rect 10612 4440 12081 4468
rect 12069 4437 12081 4440
rect 12115 4437 12127 4471
rect 12069 4431 12127 4437
rect 12250 4428 12256 4480
rect 12308 4468 12314 4480
rect 13265 4471 13323 4477
rect 13265 4468 13277 4471
rect 12308 4440 13277 4468
rect 12308 4428 12314 4440
rect 13265 4437 13277 4440
rect 13311 4437 13323 4471
rect 13265 4431 13323 4437
rect 14645 4471 14703 4477
rect 14645 4437 14657 4471
rect 14691 4468 14703 4471
rect 14918 4468 14924 4480
rect 14691 4440 14924 4468
rect 14691 4437 14703 4440
rect 14645 4431 14703 4437
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 3973 4267 4031 4273
rect 2832 4236 3648 4264
rect 2832 4224 2838 4236
rect 1026 4088 1032 4140
rect 1084 4128 1090 4140
rect 1578 4128 1584 4140
rect 1084 4100 1584 4128
rect 1084 4088 1090 4100
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4128 2283 4131
rect 2498 4128 2504 4140
rect 2271 4100 2504 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 3620 4128 3648 4236
rect 3973 4233 3985 4267
rect 4019 4264 4031 4267
rect 5166 4264 5172 4276
rect 4019 4236 5172 4264
rect 4019 4233 4031 4236
rect 3973 4227 4031 4233
rect 5166 4224 5172 4236
rect 5224 4224 5230 4276
rect 5534 4264 5540 4276
rect 5495 4236 5540 4264
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 5626 4224 5632 4276
rect 5684 4264 5690 4276
rect 6825 4267 6883 4273
rect 6825 4264 6837 4267
rect 5684 4236 6837 4264
rect 5684 4224 5690 4236
rect 6825 4233 6837 4236
rect 6871 4233 6883 4267
rect 6825 4227 6883 4233
rect 7834 4224 7840 4276
rect 7892 4264 7898 4276
rect 9122 4264 9128 4276
rect 7892 4236 9128 4264
rect 7892 4224 7898 4236
rect 9122 4224 9128 4236
rect 9180 4264 9186 4276
rect 9180 4236 10364 4264
rect 9180 4224 9186 4236
rect 4065 4199 4123 4205
rect 4065 4165 4077 4199
rect 4111 4196 4123 4199
rect 4154 4196 4160 4208
rect 4111 4168 4160 4196
rect 4111 4165 4123 4168
rect 4065 4159 4123 4165
rect 4154 4156 4160 4168
rect 4212 4156 4218 4208
rect 4338 4156 4344 4208
rect 4396 4196 4402 4208
rect 8202 4196 8208 4208
rect 4396 4168 5304 4196
rect 4396 4156 4402 4168
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 3620 4100 4721 4128
rect 4709 4097 4721 4100
rect 4755 4128 4767 4131
rect 5276 4128 5304 4168
rect 5644 4168 8208 4196
rect 5534 4128 5540 4140
rect 4755 4100 5212 4128
rect 5276 4100 5540 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 1394 4020 1400 4072
rect 1452 4060 1458 4072
rect 1946 4060 1952 4072
rect 1452 4032 1952 4060
rect 1452 4020 1458 4032
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 2590 4060 2596 4072
rect 2551 4032 2596 4060
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 4890 4060 4896 4072
rect 2700 4032 3096 4060
rect 4851 4032 4896 4060
rect 1596 3964 2268 3992
rect 1596 3933 1624 3964
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3893 1639 3927
rect 1946 3924 1952 3936
rect 1907 3896 1952 3924
rect 1581 3887 1639 3893
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 2038 3884 2044 3936
rect 2096 3924 2102 3936
rect 2240 3924 2268 3964
rect 2314 3952 2320 4004
rect 2372 3992 2378 4004
rect 2700 3992 2728 4032
rect 2372 3964 2728 3992
rect 2372 3952 2378 3964
rect 2774 3952 2780 4004
rect 2832 4001 2838 4004
rect 2832 3995 2896 4001
rect 2832 3961 2850 3995
rect 2884 3961 2896 3995
rect 3068 3992 3096 4032
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 5184 4060 5212 4100
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 5644 4060 5672 4168
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 8849 4199 8907 4205
rect 8849 4165 8861 4199
rect 8895 4196 8907 4199
rect 10042 4196 10048 4208
rect 8895 4168 10048 4196
rect 8895 4165 8907 4168
rect 8849 4159 8907 4165
rect 10042 4156 10048 4168
rect 10100 4156 10106 4208
rect 10336 4196 10364 4236
rect 11054 4224 11060 4276
rect 11112 4264 11118 4276
rect 11882 4264 11888 4276
rect 11112 4236 11888 4264
rect 11112 4224 11118 4236
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 11974 4224 11980 4276
rect 12032 4264 12038 4276
rect 15286 4264 15292 4276
rect 12032 4236 15292 4264
rect 12032 4224 12038 4236
rect 15286 4224 15292 4236
rect 15344 4224 15350 4276
rect 10336 4168 10732 4196
rect 6181 4131 6239 4137
rect 6181 4097 6193 4131
rect 6227 4097 6239 4131
rect 6181 4091 6239 4097
rect 5184 4032 5672 4060
rect 6196 4060 6224 4091
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 6972 4100 7389 4128
rect 6972 4088 6978 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 8570 4128 8576 4140
rect 7377 4091 7435 4097
rect 8220 4100 8576 4128
rect 8220 4060 8248 4100
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 9030 4088 9036 4140
rect 9088 4128 9094 4140
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 9088 4100 9321 4128
rect 9088 4088 9094 4100
rect 9309 4097 9321 4100
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 9493 4131 9551 4137
rect 9493 4097 9505 4131
rect 9539 4128 9551 4131
rect 10318 4128 10324 4140
rect 9539 4100 10324 4128
rect 9539 4097 9551 4100
rect 9493 4091 9551 4097
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 10410 4088 10416 4140
rect 10468 4128 10474 4140
rect 10704 4128 10732 4168
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 11241 4199 11299 4205
rect 11241 4196 11253 4199
rect 10928 4168 11253 4196
rect 10928 4156 10934 4168
rect 11241 4165 11253 4168
rect 11287 4165 11299 4199
rect 11241 4159 11299 4165
rect 11514 4156 11520 4208
rect 11572 4196 11578 4208
rect 12250 4196 12256 4208
rect 11572 4168 12256 4196
rect 11572 4156 11578 4168
rect 12250 4156 12256 4168
rect 12308 4156 12314 4208
rect 12437 4199 12495 4205
rect 12437 4165 12449 4199
rect 12483 4196 12495 4199
rect 12802 4196 12808 4208
rect 12483 4168 12808 4196
rect 12483 4165 12495 4168
rect 12437 4159 12495 4165
rect 12802 4156 12808 4168
rect 12860 4156 12866 4208
rect 13633 4199 13691 4205
rect 13633 4165 13645 4199
rect 13679 4196 13691 4199
rect 13722 4196 13728 4208
rect 13679 4168 13728 4196
rect 13679 4165 13691 4168
rect 13633 4159 13691 4165
rect 13722 4156 13728 4168
rect 13780 4156 13786 4208
rect 10962 4128 10968 4140
rect 10468 4100 10640 4128
rect 10704 4100 10968 4128
rect 10468 4088 10474 4100
rect 8478 4060 8484 4072
rect 6196 4032 8248 4060
rect 8439 4032 8484 4060
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 10502 4060 10508 4072
rect 10275 4032 10508 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 10612 4060 10640 4100
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 11054 4088 11060 4140
rect 11112 4128 11118 4140
rect 11839 4131 11897 4137
rect 11112 4100 11744 4128
rect 11112 4088 11118 4100
rect 10781 4063 10839 4069
rect 10781 4060 10793 4063
rect 10612 4032 10793 4060
rect 10781 4029 10793 4032
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 11330 4020 11336 4072
rect 11388 4060 11394 4072
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 11388 4032 11621 4060
rect 11388 4020 11394 4032
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 11716 4060 11744 4100
rect 11839 4097 11851 4131
rect 11885 4128 11897 4131
rect 12158 4128 12164 4140
rect 11885 4100 12164 4128
rect 11885 4097 11897 4100
rect 11839 4091 11897 4097
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12618 4088 12624 4140
rect 12676 4128 12682 4140
rect 12894 4128 12900 4140
rect 12676 4100 12900 4128
rect 12676 4088 12682 4100
rect 12894 4088 12900 4100
rect 12952 4128 12958 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12952 4100 13001 4128
rect 12952 4088 12958 4100
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 14185 4131 14243 4137
rect 14185 4128 14197 4131
rect 13596 4100 14197 4128
rect 13596 4088 13602 4100
rect 14185 4097 14197 4100
rect 14231 4097 14243 4131
rect 14185 4091 14243 4097
rect 12526 4060 12532 4072
rect 11716 4032 12532 4060
rect 11609 4023 11667 4029
rect 12526 4020 12532 4032
rect 12584 4020 12590 4072
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 12636 4032 14841 4060
rect 3068 3964 3832 3992
rect 2832 3955 2896 3961
rect 2832 3952 2838 3955
rect 3418 3924 3424 3936
rect 2096 3896 2141 3924
rect 2240 3896 3424 3924
rect 2096 3884 2102 3896
rect 3418 3884 3424 3896
rect 3476 3884 3482 3936
rect 3804 3924 3832 3964
rect 4154 3952 4160 4004
rect 4212 3992 4218 4004
rect 5169 3995 5227 4001
rect 5169 3992 5181 3995
rect 4212 3964 5181 3992
rect 4212 3952 4218 3964
rect 5169 3961 5181 3964
rect 5215 3961 5227 3995
rect 5169 3955 5227 3961
rect 5350 3952 5356 4004
rect 5408 3992 5414 4004
rect 5902 3992 5908 4004
rect 5408 3964 5908 3992
rect 5408 3952 5414 3964
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 5997 3995 6055 4001
rect 5997 3961 6009 3995
rect 6043 3992 6055 3995
rect 6546 3992 6552 4004
rect 6043 3964 6552 3992
rect 6043 3961 6055 3964
rect 5997 3955 6055 3961
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 6822 3992 6828 4004
rect 6728 3964 6828 3992
rect 4433 3927 4491 3933
rect 4433 3924 4445 3927
rect 3804 3896 4445 3924
rect 4433 3893 4445 3896
rect 4479 3893 4491 3927
rect 4433 3887 4491 3893
rect 4525 3927 4583 3933
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 6728 3924 6756 3964
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 7285 3995 7343 4001
rect 7285 3961 7297 3995
rect 7331 3992 7343 3995
rect 7466 3992 7472 4004
rect 7331 3964 7472 3992
rect 7331 3961 7343 3964
rect 7285 3955 7343 3961
rect 7466 3952 7472 3964
rect 7524 3952 7530 4004
rect 8110 3992 8116 4004
rect 7668 3964 8116 3992
rect 4571 3896 6756 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 7006 3884 7012 3936
rect 7064 3924 7070 3936
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 7064 3896 7205 3924
rect 7064 3884 7070 3896
rect 7193 3893 7205 3896
rect 7239 3924 7251 3927
rect 7668 3924 7696 3964
rect 8110 3952 8116 3964
rect 8168 3952 8174 4004
rect 8389 3995 8447 4001
rect 8389 3961 8401 3995
rect 8435 3992 8447 3995
rect 8846 3992 8852 4004
rect 8435 3964 8852 3992
rect 8435 3961 8447 3964
rect 8389 3955 8447 3961
rect 8846 3952 8852 3964
rect 8904 3952 8910 4004
rect 9217 3995 9275 4001
rect 9217 3961 9229 3995
rect 9263 3992 9275 3995
rect 10873 3995 10931 4001
rect 9263 3964 10824 3992
rect 9263 3961 9275 3964
rect 9217 3955 9275 3961
rect 7239 3896 7696 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 7742 3884 7748 3936
rect 7800 3924 7806 3936
rect 8021 3927 8079 3933
rect 8021 3924 8033 3927
rect 7800 3896 8033 3924
rect 7800 3884 7806 3896
rect 8021 3893 8033 3896
rect 8067 3893 8079 3927
rect 8021 3887 8079 3893
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 10045 3927 10103 3933
rect 10045 3924 10057 3927
rect 8352 3896 10057 3924
rect 8352 3884 8358 3896
rect 10045 3893 10057 3896
rect 10091 3893 10103 3927
rect 10410 3924 10416 3936
rect 10371 3896 10416 3924
rect 10045 3887 10103 3893
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 10796 3924 10824 3964
rect 10873 3961 10885 3995
rect 10919 3992 10931 3995
rect 11054 3992 11060 4004
rect 10919 3964 11060 3992
rect 10919 3961 10931 3964
rect 10873 3955 10931 3961
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 11514 3992 11520 4004
rect 11164 3964 11520 3992
rect 11164 3924 11192 3964
rect 11514 3952 11520 3964
rect 11572 3952 11578 4004
rect 11701 3995 11759 4001
rect 11701 3961 11713 3995
rect 11747 3992 11759 3995
rect 11882 3992 11888 4004
rect 11747 3964 11888 3992
rect 11747 3961 11759 3964
rect 11701 3955 11759 3961
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 10796 3896 11192 3924
rect 12066 3884 12072 3936
rect 12124 3924 12130 3936
rect 12636 3924 12664 4032
rect 14829 4029 14841 4032
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 13541 3995 13599 4001
rect 13541 3961 13553 3995
rect 13587 3992 13599 3995
rect 13630 3992 13636 4004
rect 13587 3964 13636 3992
rect 13587 3961 13599 3964
rect 13541 3955 13599 3961
rect 13630 3952 13636 3964
rect 13688 3992 13694 4004
rect 14001 3995 14059 4001
rect 14001 3992 14013 3995
rect 13688 3964 14013 3992
rect 13688 3952 13694 3964
rect 14001 3961 14013 3964
rect 14047 3961 14059 3995
rect 14001 3955 14059 3961
rect 14093 3995 14151 4001
rect 14093 3961 14105 3995
rect 14139 3992 14151 3995
rect 15470 3992 15476 4004
rect 14139 3964 15476 3992
rect 14139 3961 14151 3964
rect 14093 3955 14151 3961
rect 12802 3924 12808 3936
rect 12124 3896 12664 3924
rect 12763 3896 12808 3924
rect 12124 3884 12130 3896
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 12986 3924 12992 3936
rect 12943 3896 12992 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13262 3884 13268 3936
rect 13320 3924 13326 3936
rect 14108 3924 14136 3955
rect 15470 3952 15476 3964
rect 15528 3952 15534 4004
rect 15010 3924 15016 3936
rect 13320 3896 14136 3924
rect 14971 3896 15016 3924
rect 13320 3884 13326 3896
rect 15010 3884 15016 3896
rect 15068 3884 15074 3936
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 566 3680 572 3732
rect 624 3720 630 3732
rect 1486 3720 1492 3732
rect 624 3692 1492 3720
rect 624 3680 630 3692
rect 1486 3680 1492 3692
rect 1544 3680 1550 3732
rect 1854 3720 1860 3732
rect 1815 3692 1860 3720
rect 1854 3680 1860 3692
rect 1912 3680 1918 3732
rect 2869 3723 2927 3729
rect 2869 3689 2881 3723
rect 2915 3720 2927 3723
rect 3142 3720 3148 3732
rect 2915 3692 3148 3720
rect 2915 3689 2927 3692
rect 2869 3683 2927 3689
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 4154 3720 4160 3732
rect 3476 3692 4160 3720
rect 3476 3680 3482 3692
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 4433 3723 4491 3729
rect 4433 3689 4445 3723
rect 4479 3720 4491 3723
rect 5074 3720 5080 3732
rect 4479 3692 5080 3720
rect 4479 3689 4491 3692
rect 4433 3683 4491 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 6181 3723 6239 3729
rect 6181 3720 6193 3723
rect 5776 3692 6193 3720
rect 5776 3680 5782 3692
rect 6181 3689 6193 3692
rect 6227 3689 6239 3723
rect 7190 3720 7196 3732
rect 6181 3683 6239 3689
rect 6288 3692 7196 3720
rect 198 3612 204 3664
rect 256 3652 262 3664
rect 3694 3652 3700 3664
rect 256 3624 3700 3652
rect 256 3612 262 3624
rect 3694 3612 3700 3624
rect 3752 3612 3758 3664
rect 3878 3612 3884 3664
rect 3936 3652 3942 3664
rect 4525 3655 4583 3661
rect 4525 3652 4537 3655
rect 3936 3624 4537 3652
rect 3936 3612 3942 3624
rect 4525 3621 4537 3624
rect 4571 3621 4583 3655
rect 5902 3652 5908 3664
rect 4525 3615 4583 3621
rect 5184 3624 5908 3652
rect 934 3544 940 3596
rect 992 3584 998 3596
rect 1765 3587 1823 3593
rect 1765 3584 1777 3587
rect 992 3556 1777 3584
rect 992 3544 998 3556
rect 1765 3553 1777 3556
rect 1811 3553 1823 3587
rect 1765 3547 1823 3553
rect 2777 3587 2835 3593
rect 2777 3553 2789 3587
rect 2823 3584 2835 3587
rect 3234 3584 3240 3596
rect 2823 3556 3240 3584
rect 2823 3553 2835 3556
rect 2777 3547 2835 3553
rect 3234 3544 3240 3556
rect 3292 3544 3298 3596
rect 3329 3587 3387 3593
rect 3329 3553 3341 3587
rect 3375 3584 3387 3587
rect 3418 3584 3424 3596
rect 3375 3556 3424 3584
rect 3375 3553 3387 3556
rect 3329 3547 3387 3553
rect 3418 3544 3424 3556
rect 3476 3544 3482 3596
rect 3602 3544 3608 3596
rect 3660 3584 3666 3596
rect 5184 3584 5212 3624
rect 5902 3612 5908 3624
rect 5960 3612 5966 3664
rect 6086 3612 6092 3664
rect 6144 3652 6150 3664
rect 6288 3652 6316 3692
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 7377 3723 7435 3729
rect 7377 3689 7389 3723
rect 7423 3720 7435 3723
rect 8018 3720 8024 3732
rect 7423 3692 8024 3720
rect 7423 3689 7435 3692
rect 7377 3683 7435 3689
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 8205 3723 8263 3729
rect 8205 3689 8217 3723
rect 8251 3720 8263 3723
rect 9030 3720 9036 3732
rect 8251 3692 9036 3720
rect 8251 3689 8263 3692
rect 8205 3683 8263 3689
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9306 3680 9312 3732
rect 9364 3720 9370 3732
rect 10410 3720 10416 3732
rect 9364 3692 10416 3720
rect 9364 3680 9370 3692
rect 10410 3680 10416 3692
rect 10468 3680 10474 3732
rect 12802 3720 12808 3732
rect 12268 3692 12808 3720
rect 6144 3624 6316 3652
rect 6549 3655 6607 3661
rect 6144 3612 6150 3624
rect 6549 3621 6561 3655
rect 6595 3621 6607 3655
rect 6549 3615 6607 3621
rect 5350 3584 5356 3596
rect 3660 3556 5212 3584
rect 5311 3556 5356 3584
rect 3660 3544 3666 3556
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3584 5503 3587
rect 6178 3584 6184 3596
rect 5491 3556 6184 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 6564 3584 6592 3615
rect 7466 3612 7472 3664
rect 7524 3652 7530 3664
rect 7745 3655 7803 3661
rect 7745 3652 7757 3655
rect 7524 3624 7757 3652
rect 7524 3612 7530 3624
rect 7745 3621 7757 3624
rect 7791 3621 7803 3655
rect 7745 3615 7803 3621
rect 8110 3612 8116 3664
rect 8168 3652 8174 3664
rect 8665 3655 8723 3661
rect 8665 3652 8677 3655
rect 8168 3624 8677 3652
rect 8168 3612 8174 3624
rect 8665 3621 8677 3624
rect 8711 3621 8723 3655
rect 8665 3615 8723 3621
rect 10137 3655 10195 3661
rect 10137 3621 10149 3655
rect 10183 3652 10195 3655
rect 10226 3652 10232 3664
rect 10183 3624 10232 3652
rect 10183 3621 10195 3624
rect 10137 3615 10195 3621
rect 10226 3612 10232 3624
rect 10284 3612 10290 3664
rect 10318 3612 10324 3664
rect 10376 3652 10382 3664
rect 11054 3652 11060 3664
rect 10376 3624 11060 3652
rect 10376 3612 10382 3624
rect 11054 3612 11060 3624
rect 11112 3612 11118 3664
rect 11241 3655 11299 3661
rect 11241 3621 11253 3655
rect 11287 3652 11299 3655
rect 11606 3652 11612 3664
rect 11287 3624 11612 3652
rect 11287 3621 11299 3624
rect 11241 3615 11299 3621
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 7834 3584 7840 3596
rect 6288 3556 7840 3584
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 2406 3516 2412 3528
rect 2087 3488 2412 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 2406 3476 2412 3488
rect 2464 3476 2470 3528
rect 3510 3516 3516 3528
rect 3471 3488 3516 3516
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 4522 3476 4528 3528
rect 4580 3516 4586 3528
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 4580 3488 4721 3516
rect 4580 3476 4586 3488
rect 4709 3485 4721 3488
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 5166 3476 5172 3528
rect 5224 3516 5230 3528
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 5224 3488 5641 3516
rect 5224 3476 5230 3488
rect 5629 3485 5641 3488
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 1394 3448 1400 3460
rect 1355 3420 1400 3448
rect 1394 3408 1400 3420
rect 1452 3408 1458 3460
rect 1946 3408 1952 3460
rect 2004 3448 2010 3460
rect 4430 3448 4436 3460
rect 2004 3420 4436 3448
rect 2004 3408 2010 3420
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 4982 3408 4988 3460
rect 5040 3448 5046 3460
rect 5644 3448 5672 3479
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 6288 3516 6316 3556
rect 7834 3544 7840 3556
rect 7892 3584 7898 3596
rect 8573 3587 8631 3593
rect 8573 3584 8585 3587
rect 7892 3556 8585 3584
rect 7892 3544 7898 3556
rect 8573 3553 8585 3556
rect 8619 3553 8631 3587
rect 9033 3587 9091 3593
rect 9033 3584 9045 3587
rect 8573 3547 8631 3553
rect 8680 3556 9045 3584
rect 5776 3488 6316 3516
rect 5776 3476 5782 3488
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 6641 3519 6699 3525
rect 6641 3516 6653 3519
rect 6604 3488 6653 3516
rect 6604 3476 6610 3488
rect 6641 3485 6653 3488
rect 6687 3485 6699 3519
rect 6641 3479 6699 3485
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 6914 3516 6920 3528
rect 6871 3488 6920 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7374 3476 7380 3528
rect 7432 3516 7438 3528
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 7432 3488 7941 3516
rect 7432 3476 7438 3488
rect 7929 3485 7941 3488
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 8680 3516 8708 3556
rect 9033 3553 9045 3556
rect 9079 3553 9091 3587
rect 9033 3547 9091 3553
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 9548 3556 9812 3584
rect 9548 3544 9554 3556
rect 8168 3488 8708 3516
rect 8849 3519 8907 3525
rect 8168 3476 8174 3488
rect 8849 3485 8861 3519
rect 8895 3485 8907 3519
rect 8849 3479 8907 3485
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3485 9275 3519
rect 9674 3516 9680 3528
rect 9217 3479 9275 3485
rect 9600 3488 9680 3516
rect 6730 3448 6736 3460
rect 5040 3420 5085 3448
rect 5644 3420 6736 3448
rect 5040 3408 5046 3420
rect 6730 3408 6736 3420
rect 6788 3408 6794 3460
rect 8570 3408 8576 3460
rect 8628 3448 8634 3460
rect 8754 3448 8760 3460
rect 8628 3420 8760 3448
rect 8628 3408 8634 3420
rect 8754 3408 8760 3420
rect 8812 3408 8818 3460
rect 8864 3448 8892 3479
rect 9030 3448 9036 3460
rect 8864 3420 9036 3448
rect 9030 3408 9036 3420
rect 9088 3408 9094 3460
rect 4062 3380 4068 3392
rect 4023 3352 4068 3380
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 4614 3340 4620 3392
rect 4672 3380 4678 3392
rect 6086 3380 6092 3392
rect 4672 3352 6092 3380
rect 4672 3340 4678 3352
rect 6086 3340 6092 3352
rect 6144 3340 6150 3392
rect 6270 3340 6276 3392
rect 6328 3380 6334 3392
rect 9232 3380 9260 3479
rect 6328 3352 9260 3380
rect 9600 3380 9628 3488
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 9784 3516 9812 3556
rect 9950 3544 9956 3596
rect 10008 3584 10014 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 10008 3556 10057 3584
rect 10008 3544 10014 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10244 3584 10272 3612
rect 10244 3556 10548 3584
rect 10045 3547 10103 3553
rect 10318 3516 10324 3528
rect 9784 3488 10324 3516
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 10520 3516 10548 3556
rect 10594 3544 10600 3596
rect 10652 3584 10658 3596
rect 10962 3584 10968 3596
rect 10652 3556 10968 3584
rect 10652 3544 10658 3556
rect 10962 3544 10968 3556
rect 11020 3584 11026 3596
rect 11333 3587 11391 3593
rect 11333 3584 11345 3587
rect 11020 3556 11345 3584
rect 11020 3544 11026 3556
rect 11333 3553 11345 3556
rect 11379 3553 11391 3587
rect 11333 3547 11391 3553
rect 11701 3587 11759 3593
rect 11701 3553 11713 3587
rect 11747 3584 11759 3587
rect 11974 3584 11980 3596
rect 11747 3556 11980 3584
rect 11747 3553 11759 3556
rect 11701 3547 11759 3553
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 10686 3516 10692 3528
rect 10520 3488 10692 3516
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 10778 3476 10784 3528
rect 10836 3516 10842 3528
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 10836 3488 11437 3516
rect 10836 3476 10842 3488
rect 11425 3485 11437 3488
rect 11471 3485 11483 3519
rect 11425 3479 11483 3485
rect 11606 3476 11612 3528
rect 11664 3516 11670 3528
rect 12268 3516 12296 3692
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 13078 3680 13084 3732
rect 13136 3720 13142 3732
rect 13265 3723 13323 3729
rect 13265 3720 13277 3723
rect 13136 3692 13277 3720
rect 13136 3680 13142 3692
rect 13265 3689 13277 3692
rect 13311 3689 13323 3723
rect 13265 3683 13323 3689
rect 13630 3680 13636 3732
rect 13688 3720 13694 3732
rect 13725 3723 13783 3729
rect 13725 3720 13737 3723
rect 13688 3692 13737 3720
rect 13688 3680 13694 3692
rect 13725 3689 13737 3692
rect 13771 3689 13783 3723
rect 13725 3683 13783 3689
rect 12342 3612 12348 3664
rect 12400 3652 12406 3664
rect 12437 3655 12495 3661
rect 12437 3652 12449 3655
rect 12400 3624 12449 3652
rect 12400 3612 12406 3624
rect 12437 3621 12449 3624
rect 12483 3621 12495 3655
rect 12437 3615 12495 3621
rect 12526 3612 12532 3664
rect 12584 3652 12590 3664
rect 12894 3652 12900 3664
rect 12584 3624 12900 3652
rect 12584 3612 12590 3624
rect 12894 3612 12900 3624
rect 12952 3612 12958 3664
rect 13633 3587 13691 3593
rect 13633 3584 13645 3587
rect 12452 3556 13645 3584
rect 12452 3528 12480 3556
rect 13633 3553 13645 3556
rect 13679 3553 13691 3587
rect 13633 3547 13691 3553
rect 14274 3544 14280 3596
rect 14332 3584 14338 3596
rect 14461 3587 14519 3593
rect 14461 3584 14473 3587
rect 14332 3556 14473 3584
rect 14332 3544 14338 3556
rect 14461 3553 14473 3556
rect 14507 3553 14519 3587
rect 14461 3547 14519 3553
rect 11664 3488 12296 3516
rect 11664 3476 11670 3488
rect 12434 3476 12440 3528
rect 12492 3476 12498 3528
rect 12618 3516 12624 3528
rect 12579 3488 12624 3516
rect 12618 3476 12624 3488
rect 12676 3476 12682 3528
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13538 3516 13544 3528
rect 13044 3488 13544 3516
rect 13044 3476 13050 3488
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3485 13967 3519
rect 13909 3479 13967 3485
rect 10873 3451 10931 3457
rect 10873 3417 10885 3451
rect 10919 3448 10931 3451
rect 13814 3448 13820 3460
rect 10919 3420 12480 3448
rect 10919 3417 10931 3420
rect 10873 3411 10931 3417
rect 9677 3383 9735 3389
rect 9677 3380 9689 3383
rect 9600 3352 9689 3380
rect 6328 3340 6334 3352
rect 9677 3349 9689 3352
rect 9723 3349 9735 3383
rect 9677 3343 9735 3349
rect 10410 3340 10416 3392
rect 10468 3380 10474 3392
rect 11606 3380 11612 3392
rect 10468 3352 11612 3380
rect 10468 3340 10474 3352
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 11882 3380 11888 3392
rect 11843 3352 11888 3380
rect 11882 3340 11888 3352
rect 11940 3340 11946 3392
rect 12066 3380 12072 3392
rect 12027 3352 12072 3380
rect 12066 3340 12072 3352
rect 12124 3340 12130 3392
rect 12452 3380 12480 3420
rect 13096 3420 13820 3448
rect 13096 3380 13124 3420
rect 13814 3408 13820 3420
rect 13872 3408 13878 3460
rect 13924 3448 13952 3479
rect 14274 3448 14280 3460
rect 13924 3420 14280 3448
rect 14274 3408 14280 3420
rect 14332 3408 14338 3460
rect 12452 3352 13124 3380
rect 13722 3340 13728 3392
rect 13780 3380 13786 3392
rect 14645 3383 14703 3389
rect 14645 3380 14657 3383
rect 13780 3352 14657 3380
rect 13780 3340 13786 3352
rect 14645 3349 14657 3352
rect 14691 3349 14703 3383
rect 14645 3343 14703 3349
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 2406 3136 2412 3188
rect 2464 3176 2470 3188
rect 2777 3179 2835 3185
rect 2777 3176 2789 3179
rect 2464 3148 2789 3176
rect 2464 3136 2470 3148
rect 2777 3145 2789 3148
rect 2823 3145 2835 3179
rect 5074 3176 5080 3188
rect 2777 3139 2835 3145
rect 4172 3148 5080 3176
rect 2590 3000 2596 3052
rect 2648 3040 2654 3052
rect 2869 3043 2927 3049
rect 2869 3040 2881 3043
rect 2648 3012 2881 3040
rect 2648 3000 2654 3012
rect 2869 3009 2881 3012
rect 2915 3009 2927 3043
rect 2869 3003 2927 3009
rect 750 2932 756 2984
rect 808 2972 814 2984
rect 3136 2975 3194 2981
rect 808 2944 1808 2972
rect 808 2932 814 2944
rect 1664 2907 1722 2913
rect 1664 2873 1676 2907
rect 1710 2873 1722 2907
rect 1780 2904 1808 2944
rect 3136 2941 3148 2975
rect 3182 2972 3194 2975
rect 4172 2972 4200 3148
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5537 3179 5595 3185
rect 5537 3145 5549 3179
rect 5583 3176 5595 3179
rect 6546 3176 6552 3188
rect 5583 3148 6552 3176
rect 5583 3145 5595 3148
rect 5537 3139 5595 3145
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 6822 3176 6828 3188
rect 6783 3148 6828 3176
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7653 3179 7711 3185
rect 7653 3145 7665 3179
rect 7699 3176 7711 3179
rect 8018 3176 8024 3188
rect 7699 3148 8024 3176
rect 7699 3145 7711 3148
rect 7653 3139 7711 3145
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 9214 3176 9220 3188
rect 9175 3148 9220 3176
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 10042 3176 10048 3188
rect 9324 3148 10048 3176
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 5810 3108 5816 3120
rect 4387 3080 5816 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 5810 3068 5816 3080
rect 5868 3068 5874 3120
rect 7374 3108 7380 3120
rect 6012 3080 7380 3108
rect 4246 3000 4252 3052
rect 4304 3040 4310 3052
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4304 3012 4997 3040
rect 4304 3000 4310 3012
rect 4985 3009 4997 3012
rect 5031 3040 5043 3043
rect 5442 3040 5448 3052
rect 5031 3012 5448 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 5534 3000 5540 3052
rect 5592 3040 5598 3052
rect 6012 3049 6040 3080
rect 7374 3068 7380 3080
rect 7432 3108 7438 3120
rect 7432 3080 7871 3108
rect 7432 3068 7438 3080
rect 5997 3043 6055 3049
rect 5997 3040 6009 3043
rect 5592 3012 6009 3040
rect 5592 3000 5598 3012
rect 5997 3009 6009 3012
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 6181 3043 6239 3049
rect 6181 3009 6193 3043
rect 6227 3040 6239 3043
rect 6362 3040 6368 3052
rect 6227 3012 6368 3040
rect 6227 3009 6239 3012
rect 6181 3003 6239 3009
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 7282 3040 7288 3052
rect 7243 3012 7288 3040
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3040 7527 3043
rect 7558 3040 7564 3052
rect 7515 3012 7564 3040
rect 7515 3009 7527 3012
rect 7469 3003 7527 3009
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 7843 3040 7871 3080
rect 7926 3068 7932 3120
rect 7984 3108 7990 3120
rect 8849 3111 8907 3117
rect 8849 3108 8861 3111
rect 7984 3080 8861 3108
rect 7984 3068 7990 3080
rect 8849 3077 8861 3080
rect 8895 3077 8907 3111
rect 8849 3071 8907 3077
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 7843 3012 8125 3040
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 9324 3040 9352 3148
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 10318 3136 10324 3188
rect 10376 3176 10382 3188
rect 10778 3176 10784 3188
rect 10376 3148 10784 3176
rect 10376 3136 10382 3148
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 11241 3179 11299 3185
rect 11241 3176 11253 3179
rect 11204 3148 11253 3176
rect 11204 3136 11210 3148
rect 11241 3145 11253 3148
rect 11287 3145 11299 3179
rect 11241 3139 11299 3145
rect 11330 3136 11336 3188
rect 11388 3176 11394 3188
rect 11388 3148 12296 3176
rect 11388 3136 11394 3148
rect 9582 3068 9588 3120
rect 9640 3108 9646 3120
rect 10229 3111 10287 3117
rect 10229 3108 10241 3111
rect 9640 3080 10241 3108
rect 9640 3068 9646 3080
rect 10229 3077 10241 3080
rect 10275 3077 10287 3111
rect 12268 3108 12296 3148
rect 12710 3136 12716 3188
rect 12768 3176 12774 3188
rect 13265 3179 13323 3185
rect 13265 3176 13277 3179
rect 12768 3148 13277 3176
rect 12768 3136 12774 3148
rect 13265 3145 13277 3148
rect 13311 3145 13323 3179
rect 13265 3139 13323 3145
rect 16298 3108 16304 3120
rect 10229 3071 10287 3077
rect 10612 3080 12204 3108
rect 12268 3080 16304 3108
rect 8343 3012 9352 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 9398 3000 9404 3052
rect 9456 3040 9462 3052
rect 9766 3040 9772 3052
rect 9456 3012 9628 3040
rect 9727 3012 9772 3040
rect 9456 3000 9462 3012
rect 4522 2972 4528 2984
rect 3182 2944 4200 2972
rect 4264 2944 4528 2972
rect 3182 2941 3194 2944
rect 3136 2935 3194 2941
rect 4264 2904 4292 2944
rect 4522 2932 4528 2944
rect 4580 2932 4586 2984
rect 4614 2932 4620 2984
rect 4672 2972 4678 2984
rect 4709 2975 4767 2981
rect 4709 2972 4721 2975
rect 4672 2944 4721 2972
rect 4672 2932 4678 2944
rect 4709 2941 4721 2944
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 4801 2975 4859 2981
rect 4801 2941 4813 2975
rect 4847 2972 4859 2975
rect 5718 2972 5724 2984
rect 4847 2944 5724 2972
rect 4847 2941 4859 2944
rect 4801 2935 4859 2941
rect 5718 2932 5724 2944
rect 5776 2932 5782 2984
rect 5902 2972 5908 2984
rect 5863 2944 5908 2972
rect 5902 2932 5908 2944
rect 5960 2972 5966 2984
rect 7006 2972 7012 2984
rect 5960 2944 7012 2972
rect 5960 2932 5966 2944
rect 7006 2932 7012 2944
rect 7064 2932 7070 2984
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 8662 2972 8668 2984
rect 7239 2944 8668 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 8662 2932 8668 2944
rect 8720 2932 8726 2984
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 9600 2981 9628 3012
rect 9766 3000 9772 3012
rect 9824 3000 9830 3052
rect 10502 3040 10508 3052
rect 9968 3012 10508 3040
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 8996 2944 9045 2972
rect 8996 2932 9002 2944
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 9125 2975 9183 2981
rect 9125 2941 9137 2975
rect 9171 2972 9183 2975
rect 9585 2975 9643 2981
rect 9171 2944 9444 2972
rect 9171 2941 9183 2944
rect 9125 2935 9183 2941
rect 1780 2876 4292 2904
rect 1664 2867 1722 2873
rect 1679 2836 1707 2867
rect 4430 2864 4436 2916
rect 4488 2904 4494 2916
rect 9416 2904 9444 2944
rect 9585 2941 9597 2975
rect 9631 2941 9643 2975
rect 9585 2935 9643 2941
rect 9677 2975 9735 2981
rect 9677 2941 9689 2975
rect 9723 2972 9735 2975
rect 9968 2972 9996 3012
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 9723 2944 9996 2972
rect 9723 2941 9735 2944
rect 9677 2935 9735 2941
rect 10042 2932 10048 2984
rect 10100 2972 10106 2984
rect 10612 2972 10640 3080
rect 10686 3000 10692 3052
rect 10744 3040 10750 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10744 3012 10977 3040
rect 10744 3000 10750 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11793 3043 11851 3049
rect 11793 3040 11805 3043
rect 11112 3012 11805 3040
rect 11112 3000 11118 3012
rect 11793 3009 11805 3012
rect 11839 3009 11851 3043
rect 12066 3040 12072 3052
rect 11793 3003 11851 3009
rect 11900 3012 12072 3040
rect 10100 2944 10640 2972
rect 10781 2975 10839 2981
rect 10100 2932 10106 2944
rect 10781 2941 10793 2975
rect 10827 2972 10839 2975
rect 11422 2972 11428 2984
rect 10827 2944 11428 2972
rect 10827 2941 10839 2944
rect 10781 2935 10839 2941
rect 11422 2932 11428 2944
rect 11480 2932 11486 2984
rect 11606 2972 11612 2984
rect 11567 2944 11612 2972
rect 11606 2932 11612 2944
rect 11664 2932 11670 2984
rect 11701 2975 11759 2981
rect 11701 2941 11713 2975
rect 11747 2972 11759 2975
rect 11900 2972 11928 3012
rect 12066 3000 12072 3012
rect 12124 3000 12130 3052
rect 12176 3040 12204 3080
rect 16298 3068 16304 3080
rect 16356 3068 16362 3120
rect 12434 3040 12440 3052
rect 12176 3012 12440 3040
rect 12434 3000 12440 3012
rect 12492 3000 12498 3052
rect 12526 3000 12532 3052
rect 12584 3040 12590 3052
rect 12986 3040 12992 3052
rect 12584 3012 12992 3040
rect 12584 3000 12590 3012
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 13078 3000 13084 3052
rect 13136 3040 13142 3052
rect 13817 3043 13875 3049
rect 13817 3040 13829 3043
rect 13136 3012 13829 3040
rect 13136 3000 13142 3012
rect 13817 3009 13829 3012
rect 13863 3009 13875 3043
rect 13817 3003 13875 3009
rect 13906 3000 13912 3052
rect 13964 3040 13970 3052
rect 14366 3040 14372 3052
rect 13964 3012 14136 3040
rect 14327 3012 14372 3040
rect 13964 3000 13970 3012
rect 12618 2972 12624 2984
rect 11747 2944 11928 2972
rect 11992 2944 12624 2972
rect 11747 2941 11759 2944
rect 11701 2935 11759 2941
rect 9930 2904 9936 2916
rect 4488 2876 9352 2904
rect 9416 2876 9936 2904
rect 4488 2864 4494 2876
rect 2314 2836 2320 2848
rect 1679 2808 2320 2836
rect 2314 2796 2320 2808
rect 2372 2796 2378 2848
rect 4249 2839 4307 2845
rect 4249 2805 4261 2839
rect 4295 2836 4307 2839
rect 4798 2836 4804 2848
rect 4295 2808 4804 2836
rect 4295 2805 4307 2808
rect 4249 2799 4307 2805
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 5350 2796 5356 2848
rect 5408 2836 5414 2848
rect 6914 2836 6920 2848
rect 5408 2808 6920 2836
rect 5408 2796 5414 2808
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7006 2796 7012 2848
rect 7064 2836 7070 2848
rect 8021 2839 8079 2845
rect 8021 2836 8033 2839
rect 7064 2808 8033 2836
rect 7064 2796 7070 2808
rect 8021 2805 8033 2808
rect 8067 2836 8079 2839
rect 9125 2839 9183 2845
rect 9125 2836 9137 2839
rect 8067 2808 9137 2836
rect 8067 2805 8079 2808
rect 8021 2799 8079 2805
rect 9125 2805 9137 2808
rect 9171 2805 9183 2839
rect 9324 2836 9352 2876
rect 9930 2864 9936 2876
rect 9988 2864 9994 2916
rect 10962 2904 10968 2916
rect 10060 2876 10456 2904
rect 10060 2836 10088 2876
rect 10428 2845 10456 2876
rect 10520 2876 10968 2904
rect 10520 2848 10548 2876
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 11146 2864 11152 2916
rect 11204 2904 11210 2916
rect 11790 2904 11796 2916
rect 11204 2876 11796 2904
rect 11204 2864 11210 2876
rect 11790 2864 11796 2876
rect 11848 2864 11854 2916
rect 9324 2808 10088 2836
rect 10413 2839 10471 2845
rect 9125 2799 9183 2805
rect 10413 2805 10425 2839
rect 10459 2805 10471 2839
rect 10413 2799 10471 2805
rect 10502 2796 10508 2848
rect 10560 2796 10566 2848
rect 10594 2796 10600 2848
rect 10652 2836 10658 2848
rect 10873 2839 10931 2845
rect 10873 2836 10885 2839
rect 10652 2808 10885 2836
rect 10652 2796 10658 2808
rect 10873 2805 10885 2808
rect 10919 2805 10931 2839
rect 10873 2799 10931 2805
rect 11422 2796 11428 2848
rect 11480 2836 11486 2848
rect 11992 2836 12020 2944
rect 12618 2932 12624 2944
rect 12676 2932 12682 2984
rect 14108 2981 14136 3012
rect 14366 3000 14372 3012
rect 14424 3000 14430 3052
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 14608 3012 14688 3040
rect 14608 3000 14614 3012
rect 14660 2981 14688 3012
rect 14093 2975 14151 2981
rect 12820 2944 13952 2972
rect 12158 2864 12164 2916
rect 12216 2904 12222 2916
rect 12820 2913 12848 2944
rect 12805 2907 12863 2913
rect 12805 2904 12817 2907
rect 12216 2876 12817 2904
rect 12216 2864 12222 2876
rect 12805 2873 12817 2876
rect 12851 2873 12863 2907
rect 12805 2867 12863 2873
rect 13725 2907 13783 2913
rect 13725 2873 13737 2907
rect 13771 2904 13783 2907
rect 13814 2904 13820 2916
rect 13771 2876 13820 2904
rect 13771 2873 13783 2876
rect 13725 2867 13783 2873
rect 13814 2864 13820 2876
rect 13872 2864 13878 2916
rect 13924 2904 13952 2944
rect 14093 2941 14105 2975
rect 14139 2941 14151 2975
rect 14093 2935 14151 2941
rect 14645 2975 14703 2981
rect 14645 2941 14657 2975
rect 14691 2941 14703 2975
rect 14645 2935 14703 2941
rect 14550 2904 14556 2916
rect 13924 2876 14556 2904
rect 14550 2864 14556 2876
rect 14608 2904 14614 2916
rect 15194 2904 15200 2916
rect 14608 2876 15200 2904
rect 14608 2864 14614 2876
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 11480 2808 12020 2836
rect 11480 2796 11486 2808
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12897 2839 12955 2845
rect 12492 2808 12537 2836
rect 12492 2796 12498 2808
rect 12897 2805 12909 2839
rect 12943 2836 12955 2839
rect 13633 2839 13691 2845
rect 13633 2836 13645 2839
rect 12943 2808 13645 2836
rect 12943 2805 12955 2808
rect 12897 2799 12955 2805
rect 13633 2805 13645 2808
rect 13679 2836 13691 2839
rect 13998 2836 14004 2848
rect 13679 2808 14004 2836
rect 13679 2805 13691 2808
rect 13633 2799 13691 2805
rect 13998 2796 14004 2808
rect 14056 2796 14062 2848
rect 14090 2796 14096 2848
rect 14148 2836 14154 2848
rect 14829 2839 14887 2845
rect 14829 2836 14841 2839
rect 14148 2808 14841 2836
rect 14148 2796 14154 2808
rect 14829 2805 14841 2808
rect 14875 2805 14887 2839
rect 14829 2799 14887 2805
rect 15102 2796 15108 2848
rect 15160 2836 15166 2848
rect 16758 2836 16764 2848
rect 15160 2808 16764 2836
rect 15160 2796 15166 2808
rect 16758 2796 16764 2808
rect 16816 2796 16822 2848
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 2590 2632 2596 2644
rect 1412 2604 2596 2632
rect 1412 2505 1440 2604
rect 2590 2592 2596 2604
rect 2648 2592 2654 2644
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 3142 2632 3148 2644
rect 2915 2604 3148 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 3142 2592 3148 2604
rect 3200 2592 3206 2644
rect 3237 2635 3295 2641
rect 3237 2601 3249 2635
rect 3283 2632 3295 2635
rect 3326 2632 3332 2644
rect 3283 2604 3332 2632
rect 3283 2601 3295 2604
rect 3237 2595 3295 2601
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4212 2604 4292 2632
rect 4212 2592 4218 2604
rect 1762 2524 1768 2576
rect 1820 2564 1826 2576
rect 4264 2564 4292 2604
rect 4890 2592 4896 2644
rect 4948 2632 4954 2644
rect 5445 2635 5503 2641
rect 5445 2632 5457 2635
rect 4948 2604 5457 2632
rect 4948 2592 4954 2604
rect 5445 2601 5457 2604
rect 5491 2601 5503 2635
rect 5445 2595 5503 2601
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 5905 2635 5963 2641
rect 5905 2632 5917 2635
rect 5868 2604 5917 2632
rect 5868 2592 5874 2604
rect 5905 2601 5917 2604
rect 5951 2601 5963 2635
rect 5905 2595 5963 2601
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2601 6975 2635
rect 8570 2632 8576 2644
rect 8531 2604 8576 2632
rect 6917 2595 6975 2601
rect 6549 2567 6607 2573
rect 6549 2564 6561 2567
rect 1820 2536 2643 2564
rect 4264 2536 5856 2564
rect 1820 2524 1826 2536
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 1664 2499 1722 2505
rect 1664 2465 1676 2499
rect 1710 2496 1722 2499
rect 2406 2496 2412 2508
rect 1710 2468 2412 2496
rect 1710 2465 1722 2468
rect 1664 2459 1722 2465
rect 2406 2456 2412 2468
rect 2464 2456 2470 2508
rect 2615 2496 2643 2536
rect 4614 2496 4620 2508
rect 2615 2468 4476 2496
rect 4575 2468 4620 2496
rect 3326 2428 3332 2440
rect 3287 2400 3332 2428
rect 3326 2388 3332 2400
rect 3384 2388 3390 2440
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 4338 2428 4344 2440
rect 3559 2400 4344 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 4448 2428 4476 2468
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 4709 2499 4767 2505
rect 4709 2465 4721 2499
rect 4755 2496 4767 2499
rect 5626 2496 5632 2508
rect 4755 2468 5632 2496
rect 4755 2465 4767 2468
rect 4709 2459 4767 2465
rect 4724 2428 4752 2459
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 5828 2505 5856 2536
rect 5920 2536 6561 2564
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2465 5871 2499
rect 5813 2459 5871 2465
rect 4448 2400 4752 2428
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2428 4951 2431
rect 5166 2428 5172 2440
rect 4939 2400 5172 2428
rect 4939 2397 4951 2400
rect 4893 2391 4951 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5920 2428 5948 2536
rect 6549 2533 6561 2536
rect 6595 2533 6607 2567
rect 6549 2527 6607 2533
rect 6273 2499 6331 2505
rect 6273 2465 6285 2499
rect 6319 2496 6331 2499
rect 6932 2496 6960 2595
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 8938 2632 8944 2644
rect 8711 2604 8944 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 8938 2592 8944 2604
rect 8996 2592 9002 2644
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 10229 2635 10287 2641
rect 9088 2604 10088 2632
rect 9088 2592 9094 2604
rect 7285 2567 7343 2573
rect 7285 2533 7297 2567
rect 7331 2564 7343 2567
rect 9950 2564 9956 2576
rect 7331 2536 9956 2564
rect 7331 2533 7343 2536
rect 7285 2527 7343 2533
rect 9950 2524 9956 2536
rect 10008 2524 10014 2576
rect 6319 2468 6960 2496
rect 6319 2465 6331 2468
rect 6273 2459 6331 2465
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 7064 2468 7512 2496
rect 7064 2456 7070 2468
rect 5276 2400 5948 2428
rect 6089 2431 6147 2437
rect 3970 2360 3976 2372
rect 2424 2332 3976 2360
rect 1394 2252 1400 2304
rect 1452 2292 1458 2304
rect 2424 2292 2452 2332
rect 3970 2320 3976 2332
rect 4028 2320 4034 2372
rect 4430 2360 4436 2372
rect 4264 2332 4436 2360
rect 1452 2264 2452 2292
rect 1452 2252 1458 2264
rect 2498 2252 2504 2304
rect 2556 2292 2562 2304
rect 2777 2295 2835 2301
rect 2777 2292 2789 2295
rect 2556 2264 2789 2292
rect 2556 2252 2562 2264
rect 2777 2261 2789 2264
rect 2823 2292 2835 2295
rect 4154 2292 4160 2304
rect 2823 2264 4160 2292
rect 2823 2261 2835 2264
rect 2777 2255 2835 2261
rect 4154 2252 4160 2264
rect 4212 2252 4218 2304
rect 4264 2301 4292 2332
rect 4430 2320 4436 2332
rect 4488 2320 4494 2372
rect 4249 2295 4307 2301
rect 4249 2261 4261 2295
rect 4295 2261 4307 2295
rect 4249 2255 4307 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 5276 2292 5304 2400
rect 6089 2397 6101 2431
rect 6135 2428 6147 2431
rect 6454 2428 6460 2440
rect 6135 2400 6460 2428
rect 6135 2397 6147 2400
rect 6089 2391 6147 2397
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 7484 2437 7512 2468
rect 8202 2456 8208 2508
rect 8260 2496 8266 2508
rect 10060 2496 10088 2604
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 11146 2632 11152 2644
rect 10275 2604 11152 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11425 2635 11483 2641
rect 11425 2601 11437 2635
rect 11471 2632 11483 2635
rect 12434 2632 12440 2644
rect 11471 2604 12440 2632
rect 11471 2601 11483 2604
rect 11425 2595 11483 2601
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 12618 2632 12624 2644
rect 12579 2604 12624 2632
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 13078 2592 13084 2644
rect 13136 2632 13142 2644
rect 13262 2632 13268 2644
rect 13136 2604 13268 2632
rect 13136 2592 13142 2604
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 13909 2635 13967 2641
rect 13909 2632 13921 2635
rect 13872 2604 13921 2632
rect 13872 2592 13878 2604
rect 13909 2601 13921 2604
rect 13955 2601 13967 2635
rect 13909 2595 13967 2601
rect 14826 2592 14832 2644
rect 14884 2592 14890 2644
rect 10137 2567 10195 2573
rect 10137 2533 10149 2567
rect 10183 2564 10195 2567
rect 11054 2564 11060 2576
rect 10183 2536 11060 2564
rect 10183 2533 10195 2536
rect 10137 2527 10195 2533
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 11333 2567 11391 2573
rect 11333 2533 11345 2567
rect 11379 2564 11391 2567
rect 13630 2564 13636 2576
rect 11379 2536 13636 2564
rect 11379 2533 11391 2536
rect 11333 2527 11391 2533
rect 13630 2524 13636 2536
rect 13688 2524 13694 2576
rect 14844 2564 14872 2592
rect 15102 2564 15108 2576
rect 14108 2536 14872 2564
rect 15063 2536 15108 2564
rect 11422 2496 11428 2508
rect 8260 2468 9976 2496
rect 10060 2468 11428 2496
rect 8260 2456 8266 2468
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 8849 2431 8907 2437
rect 8849 2397 8861 2431
rect 8895 2428 8907 2431
rect 9122 2428 9128 2440
rect 8895 2400 9128 2428
rect 8895 2397 8907 2400
rect 8849 2391 8907 2397
rect 5442 2320 5448 2372
rect 5500 2360 5506 2372
rect 7392 2360 7420 2391
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 5500 2332 7420 2360
rect 8205 2363 8263 2369
rect 5500 2320 5506 2332
rect 8205 2329 8217 2363
rect 8251 2360 8263 2363
rect 9398 2360 9404 2372
rect 8251 2332 9404 2360
rect 8251 2329 8263 2332
rect 8205 2323 8263 2329
rect 9398 2320 9404 2332
rect 9456 2320 9462 2372
rect 9948 2360 9976 2468
rect 11422 2456 11428 2468
rect 11480 2456 11486 2508
rect 11974 2496 11980 2508
rect 11935 2468 11980 2496
rect 11974 2456 11980 2468
rect 12032 2456 12038 2508
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 12989 2499 13047 2505
rect 12989 2496 13001 2499
rect 12124 2468 13001 2496
rect 12124 2456 12130 2468
rect 12989 2465 13001 2468
rect 13035 2465 13047 2499
rect 12989 2459 13047 2465
rect 13817 2499 13875 2505
rect 13817 2465 13829 2499
rect 13863 2496 13875 2499
rect 13998 2496 14004 2508
rect 13863 2468 14004 2496
rect 13863 2465 13875 2468
rect 13817 2459 13875 2465
rect 13998 2456 14004 2468
rect 14056 2456 14062 2508
rect 10318 2428 10324 2440
rect 10279 2400 10324 2428
rect 10318 2388 10324 2400
rect 10376 2428 10382 2440
rect 10686 2428 10692 2440
rect 10376 2400 10692 2428
rect 10376 2388 10382 2400
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 11532 2360 11560 2391
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 12161 2431 12219 2437
rect 12161 2428 12173 2431
rect 11664 2400 12173 2428
rect 11664 2388 11670 2400
rect 12161 2397 12173 2400
rect 12207 2397 12219 2431
rect 12161 2391 12219 2397
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 12952 2400 13093 2428
rect 12952 2388 12958 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 13262 2388 13268 2440
rect 13320 2428 13326 2440
rect 14108 2437 14136 2536
rect 15102 2524 15108 2536
rect 15160 2524 15166 2576
rect 14274 2496 14280 2508
rect 14235 2468 14280 2496
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 14826 2496 14832 2508
rect 14787 2468 14832 2496
rect 14826 2456 14832 2468
rect 14884 2456 14890 2508
rect 14093 2431 14151 2437
rect 13320 2400 13365 2428
rect 13320 2388 13326 2400
rect 14093 2397 14105 2431
rect 14139 2397 14151 2431
rect 14458 2428 14464 2440
rect 14419 2400 14464 2428
rect 14093 2391 14151 2397
rect 14458 2388 14464 2400
rect 14516 2388 14522 2440
rect 9948 2332 11560 2360
rect 13449 2363 13507 2369
rect 13449 2329 13461 2363
rect 13495 2360 13507 2363
rect 14734 2360 14740 2372
rect 13495 2332 14740 2360
rect 13495 2329 13507 2332
rect 13449 2323 13507 2329
rect 14734 2320 14740 2332
rect 14792 2320 14798 2372
rect 4580 2264 5304 2292
rect 4580 2252 4586 2264
rect 6270 2252 6276 2304
rect 6328 2292 6334 2304
rect 9769 2295 9827 2301
rect 9769 2292 9781 2295
rect 6328 2264 9781 2292
rect 6328 2252 6334 2264
rect 9769 2261 9781 2264
rect 9815 2261 9827 2295
rect 9769 2255 9827 2261
rect 9950 2252 9956 2304
rect 10008 2292 10014 2304
rect 10965 2295 11023 2301
rect 10965 2292 10977 2295
rect 10008 2264 10977 2292
rect 10008 2252 10014 2264
rect 10965 2261 10977 2264
rect 11011 2261 11023 2295
rect 10965 2255 11023 2261
rect 11054 2252 11060 2304
rect 11112 2292 11118 2304
rect 11698 2292 11704 2304
rect 11112 2264 11704 2292
rect 11112 2252 11118 2264
rect 11698 2252 11704 2264
rect 11756 2292 11762 2304
rect 15470 2292 15476 2304
rect 11756 2264 15476 2292
rect 11756 2252 11762 2264
rect 15470 2252 15476 2264
rect 15528 2252 15534 2304
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 842 2048 848 2100
rect 900 2088 906 2100
rect 11606 2088 11612 2100
rect 900 2060 11612 2088
rect 900 2048 906 2060
rect 11606 2048 11612 2060
rect 11664 2048 11670 2100
rect 12158 2048 12164 2100
rect 12216 2088 12222 2100
rect 13906 2088 13912 2100
rect 12216 2060 13912 2088
rect 12216 2048 12222 2060
rect 13906 2048 13912 2060
rect 13964 2048 13970 2100
rect 3326 1980 3332 2032
rect 3384 2020 3390 2032
rect 9674 2020 9680 2032
rect 3384 1992 9680 2020
rect 3384 1980 3390 1992
rect 9674 1980 9680 1992
rect 9732 1980 9738 2032
rect 9769 2023 9827 2029
rect 9769 1989 9781 2023
rect 9815 2020 9827 2023
rect 14458 2020 14464 2032
rect 9815 1992 14464 2020
rect 9815 1989 9827 1992
rect 9769 1983 9827 1989
rect 14458 1980 14464 1992
rect 14516 1980 14522 2032
rect 3786 1912 3792 1964
rect 3844 1952 3850 1964
rect 11974 1952 11980 1964
rect 3844 1924 11980 1952
rect 3844 1912 3850 1924
rect 11974 1912 11980 1924
rect 12032 1912 12038 1964
rect 12342 1912 12348 1964
rect 12400 1952 12406 1964
rect 15378 1952 15384 1964
rect 12400 1924 15384 1952
rect 12400 1912 12406 1924
rect 15378 1912 15384 1924
rect 15436 1952 15442 1964
rect 15930 1952 15936 1964
rect 15436 1924 15936 1952
rect 15436 1912 15442 1924
rect 15930 1912 15936 1924
rect 15988 1912 15994 1964
rect 1210 1844 1216 1896
rect 1268 1884 1274 1896
rect 5994 1884 6000 1896
rect 1268 1856 6000 1884
rect 1268 1844 1274 1856
rect 5994 1844 6000 1856
rect 6052 1844 6058 1896
rect 7374 1844 7380 1896
rect 7432 1884 7438 1896
rect 8478 1884 8484 1896
rect 7432 1856 8484 1884
rect 7432 1844 7438 1856
rect 8478 1844 8484 1856
rect 8536 1884 8542 1896
rect 8754 1884 8760 1896
rect 8536 1856 8760 1884
rect 8536 1844 8542 1856
rect 8754 1844 8760 1856
rect 8812 1844 8818 1896
rect 10134 1844 10140 1896
rect 10192 1884 10198 1896
rect 14182 1884 14188 1896
rect 10192 1856 14188 1884
rect 10192 1844 10198 1856
rect 14182 1844 14188 1856
rect 14240 1844 14246 1896
rect 4430 1776 4436 1828
rect 4488 1816 4494 1828
rect 11238 1816 11244 1828
rect 4488 1788 11244 1816
rect 4488 1776 4494 1788
rect 11238 1776 11244 1788
rect 11296 1776 11302 1828
rect 2406 1708 2412 1760
rect 2464 1748 2470 1760
rect 10318 1748 10324 1760
rect 2464 1720 10324 1748
rect 2464 1708 2470 1720
rect 10318 1708 10324 1720
rect 10376 1708 10382 1760
rect 10410 1708 10416 1760
rect 10468 1748 10474 1760
rect 14918 1748 14924 1760
rect 10468 1720 14924 1748
rect 10468 1708 10474 1720
rect 14918 1708 14924 1720
rect 14976 1708 14982 1760
rect 2038 1640 2044 1692
rect 2096 1680 2102 1692
rect 6270 1680 6276 1692
rect 2096 1652 6276 1680
rect 2096 1640 2102 1652
rect 6270 1640 6276 1652
rect 6328 1640 6334 1692
rect 7926 1640 7932 1692
rect 7984 1680 7990 1692
rect 9582 1680 9588 1692
rect 7984 1652 9588 1680
rect 7984 1640 7990 1652
rect 9582 1640 9588 1652
rect 9640 1640 9646 1692
rect 3970 1572 3976 1624
rect 4028 1612 4034 1624
rect 11882 1612 11888 1624
rect 4028 1584 11888 1612
rect 4028 1572 4034 1584
rect 11882 1572 11888 1584
rect 11940 1572 11946 1624
rect 2866 1504 2872 1556
rect 2924 1544 2930 1556
rect 9769 1547 9827 1553
rect 9769 1544 9781 1547
rect 2924 1516 9781 1544
rect 2924 1504 2930 1516
rect 9769 1513 9781 1516
rect 9815 1513 9827 1547
rect 9769 1507 9827 1513
rect 5350 1436 5356 1488
rect 5408 1476 5414 1488
rect 14826 1476 14832 1488
rect 5408 1448 14832 1476
rect 5408 1436 5414 1448
rect 14826 1436 14832 1448
rect 14884 1436 14890 1488
rect 8662 1368 8668 1420
rect 8720 1408 8726 1420
rect 12618 1408 12624 1420
rect 8720 1380 12624 1408
rect 8720 1368 8726 1380
rect 12618 1368 12624 1380
rect 12676 1368 12682 1420
rect 7834 1300 7840 1352
rect 7892 1340 7898 1352
rect 9306 1340 9312 1352
rect 7892 1312 9312 1340
rect 7892 1300 7898 1312
rect 9306 1300 9312 1312
rect 9364 1300 9370 1352
rect 7098 1232 7104 1284
rect 7156 1272 7162 1284
rect 10962 1272 10968 1284
rect 7156 1244 10968 1272
rect 7156 1232 7162 1244
rect 10962 1232 10968 1244
rect 11020 1232 11026 1284
rect 8846 1164 8852 1216
rect 8904 1204 8910 1216
rect 10226 1204 10232 1216
rect 8904 1176 10232 1204
rect 8904 1164 8910 1176
rect 10226 1164 10232 1176
rect 10284 1164 10290 1216
<< via1 >>
rect 572 18368 624 18420
rect 9128 18368 9180 18420
rect 8208 18164 8260 18216
rect 8760 18164 8812 18216
rect 1768 18096 1820 18148
rect 9680 18096 9732 18148
rect 11060 18096 11112 18148
rect 7472 18028 7524 18080
rect 10600 18028 10652 18080
rect 4068 17960 4120 18012
rect 12992 17960 13044 18012
rect 12808 17892 12860 17944
rect 7840 17824 7892 17876
rect 12624 17824 12676 17876
rect 3424 17756 3476 17808
rect 9404 17756 9456 17808
rect 12532 17756 12584 17808
rect 2228 17688 2280 17740
rect 8300 17688 8352 17740
rect 8944 17688 8996 17740
rect 7012 17620 7064 17672
rect 12164 17620 12216 17672
rect 13544 17620 13596 17672
rect 14464 17620 14516 17672
rect 1308 17552 1360 17604
rect 5448 17552 5500 17604
rect 8668 17552 8720 17604
rect 15200 17552 15252 17604
rect 15936 17552 15988 17604
rect 1400 17484 1452 17536
rect 7288 17484 7340 17536
rect 7564 17484 7616 17536
rect 10324 17484 10376 17536
rect 10784 17484 10836 17536
rect 11244 17484 11296 17536
rect 3447 17382 3499 17434
rect 3511 17382 3563 17434
rect 3575 17382 3627 17434
rect 3639 17382 3691 17434
rect 8378 17382 8430 17434
rect 8442 17382 8494 17434
rect 8506 17382 8558 17434
rect 8570 17382 8622 17434
rect 13308 17382 13360 17434
rect 13372 17382 13424 17434
rect 13436 17382 13488 17434
rect 13500 17382 13552 17434
rect 7288 17280 7340 17332
rect 10784 17280 10836 17332
rect 11244 17280 11296 17332
rect 12624 17280 12676 17332
rect 3608 17144 3660 17196
rect 5540 17212 5592 17264
rect 7380 17212 7432 17264
rect 2136 17051 2188 17060
rect 2136 17017 2145 17051
rect 2145 17017 2179 17051
rect 2179 17017 2188 17051
rect 2136 17008 2188 17017
rect 5356 17076 5408 17128
rect 7656 17144 7708 17196
rect 8116 17212 8168 17264
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 12072 17212 12124 17264
rect 6736 17076 6788 17128
rect 7012 17076 7064 17128
rect 9128 17076 9180 17128
rect 10508 17076 10560 17128
rect 11980 17144 12032 17196
rect 12992 17144 13044 17196
rect 13728 17144 13780 17196
rect 3056 17051 3108 17060
rect 3056 17017 3065 17051
rect 3065 17017 3099 17051
rect 3099 17017 3108 17051
rect 3056 17008 3108 17017
rect 4344 17008 4396 17060
rect 6368 17008 6420 17060
rect 7564 17051 7616 17060
rect 7564 17017 7573 17051
rect 7573 17017 7607 17051
rect 7607 17017 7616 17051
rect 7564 17008 7616 17017
rect 4712 16940 4764 16992
rect 5632 16983 5684 16992
rect 5632 16949 5641 16983
rect 5641 16949 5675 16983
rect 5675 16949 5684 16983
rect 5632 16940 5684 16949
rect 6552 16940 6604 16992
rect 7932 16940 7984 16992
rect 8392 16983 8444 16992
rect 8392 16949 8401 16983
rect 8401 16949 8435 16983
rect 8435 16949 8444 16983
rect 8392 16940 8444 16949
rect 9864 17008 9916 17060
rect 10048 17008 10100 17060
rect 13176 17076 13228 17128
rect 13636 17051 13688 17060
rect 13636 17017 13645 17051
rect 13645 17017 13679 17051
rect 13679 17017 13688 17051
rect 13636 17008 13688 17017
rect 9588 16940 9640 16992
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 10416 16940 10468 16992
rect 10600 16940 10652 16992
rect 5912 16838 5964 16890
rect 5976 16838 6028 16890
rect 6040 16838 6092 16890
rect 6104 16838 6156 16890
rect 10843 16838 10895 16890
rect 10907 16838 10959 16890
rect 10971 16838 11023 16890
rect 11035 16838 11087 16890
rect 4620 16736 4672 16788
rect 5264 16736 5316 16788
rect 6276 16736 6328 16788
rect 7288 16779 7340 16788
rect 7288 16745 7297 16779
rect 7297 16745 7331 16779
rect 7331 16745 7340 16779
rect 7288 16736 7340 16745
rect 7564 16736 7616 16788
rect 8392 16736 8444 16788
rect 8668 16736 8720 16788
rect 8944 16736 8996 16788
rect 12532 16779 12584 16788
rect 10508 16668 10560 16720
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 12808 16736 12860 16788
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 2504 16643 2556 16652
rect 2504 16609 2513 16643
rect 2513 16609 2547 16643
rect 2547 16609 2556 16643
rect 2504 16600 2556 16609
rect 3332 16600 3384 16652
rect 3608 16643 3660 16652
rect 3608 16609 3617 16643
rect 3617 16609 3651 16643
rect 3651 16609 3660 16643
rect 3608 16600 3660 16609
rect 4436 16600 4488 16652
rect 7196 16600 7248 16652
rect 6644 16532 6696 16584
rect 8208 16532 8260 16584
rect 9036 16600 9088 16652
rect 9220 16600 9272 16652
rect 10048 16643 10100 16652
rect 10048 16609 10057 16643
rect 10057 16609 10091 16643
rect 10091 16609 10100 16643
rect 10048 16600 10100 16609
rect 10416 16600 10468 16652
rect 11244 16600 11296 16652
rect 11612 16643 11664 16652
rect 11612 16609 11621 16643
rect 11621 16609 11655 16643
rect 11655 16609 11664 16643
rect 11612 16600 11664 16609
rect 11704 16600 11756 16652
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 8576 16532 8628 16584
rect 3148 16464 3200 16516
rect 204 16396 256 16448
rect 4068 16396 4120 16448
rect 4252 16396 4304 16448
rect 4712 16396 4764 16448
rect 4988 16396 5040 16448
rect 9312 16532 9364 16584
rect 10140 16575 10192 16584
rect 10140 16541 10149 16575
rect 10149 16541 10183 16575
rect 10183 16541 10192 16575
rect 10140 16532 10192 16541
rect 10968 16532 11020 16584
rect 14004 16532 14056 16584
rect 5816 16396 5868 16448
rect 5908 16396 5960 16448
rect 6920 16396 6972 16448
rect 8208 16396 8260 16448
rect 11612 16464 11664 16516
rect 8852 16396 8904 16448
rect 11152 16396 11204 16448
rect 11888 16396 11940 16448
rect 12164 16396 12216 16448
rect 14280 16396 14332 16448
rect 14556 16396 14608 16448
rect 3447 16294 3499 16346
rect 3511 16294 3563 16346
rect 3575 16294 3627 16346
rect 3639 16294 3691 16346
rect 8378 16294 8430 16346
rect 8442 16294 8494 16346
rect 8506 16294 8558 16346
rect 8570 16294 8622 16346
rect 13308 16294 13360 16346
rect 13372 16294 13424 16346
rect 13436 16294 13488 16346
rect 13500 16294 13552 16346
rect 2872 16192 2924 16244
rect 5724 16192 5776 16244
rect 7012 16192 7064 16244
rect 7104 16192 7156 16244
rect 8852 16192 8904 16244
rect 2780 16056 2832 16108
rect 3976 16124 4028 16176
rect 5172 16124 5224 16176
rect 5264 16124 5316 16176
rect 4620 16056 4672 16108
rect 4804 16099 4856 16108
rect 4804 16065 4813 16099
rect 4813 16065 4847 16099
rect 4847 16065 4856 16099
rect 4804 16056 4856 16065
rect 4988 16099 5040 16108
rect 4988 16065 4997 16099
rect 4997 16065 5031 16099
rect 5031 16065 5040 16099
rect 4988 16056 5040 16065
rect 5908 16056 5960 16108
rect 7196 16056 7248 16108
rect 7472 16056 7524 16108
rect 5080 15988 5132 16040
rect 2320 15920 2372 15972
rect 2780 15852 2832 15904
rect 3240 15852 3292 15904
rect 4896 15852 4948 15904
rect 5080 15852 5132 15904
rect 7472 15920 7524 15972
rect 7564 15920 7616 15972
rect 7748 16056 7800 16108
rect 9772 16192 9824 16244
rect 10968 16192 11020 16244
rect 11336 16192 11388 16244
rect 9680 16124 9732 16176
rect 11888 16124 11940 16176
rect 9128 16056 9180 16108
rect 9496 16056 9548 16108
rect 10968 16099 11020 16108
rect 8024 15988 8076 16040
rect 8300 15988 8352 16040
rect 9220 15988 9272 16040
rect 10968 16065 10977 16099
rect 10977 16065 11011 16099
rect 11011 16065 11020 16099
rect 10968 16056 11020 16065
rect 12716 16056 12768 16108
rect 11428 15988 11480 16040
rect 11704 15988 11756 16040
rect 12992 16056 13044 16108
rect 16764 16056 16816 16108
rect 7104 15852 7156 15904
rect 7288 15895 7340 15904
rect 7288 15861 7297 15895
rect 7297 15861 7331 15895
rect 7331 15861 7340 15895
rect 7288 15852 7340 15861
rect 9128 15920 9180 15972
rect 8484 15852 8536 15904
rect 9588 15852 9640 15904
rect 9772 15852 9824 15904
rect 10140 15852 10192 15904
rect 12900 15988 12952 16040
rect 14648 16031 14700 16040
rect 14648 15997 14657 16031
rect 14657 15997 14691 16031
rect 14691 15997 14700 16031
rect 14648 15988 14700 15997
rect 11244 15852 11296 15904
rect 12808 15852 12860 15904
rect 13636 15852 13688 15904
rect 5912 15750 5964 15802
rect 5976 15750 6028 15802
rect 6040 15750 6092 15802
rect 6104 15750 6156 15802
rect 10843 15750 10895 15802
rect 10907 15750 10959 15802
rect 10971 15750 11023 15802
rect 11035 15750 11087 15802
rect 5080 15648 5132 15700
rect 5356 15691 5408 15700
rect 5356 15657 5365 15691
rect 5365 15657 5399 15691
rect 5399 15657 5408 15691
rect 5356 15648 5408 15657
rect 6920 15691 6972 15700
rect 6920 15657 6929 15691
rect 6929 15657 6963 15691
rect 6963 15657 6972 15691
rect 6920 15648 6972 15657
rect 9772 15648 9824 15700
rect 10416 15648 10468 15700
rect 10692 15648 10744 15700
rect 12256 15648 12308 15700
rect 13452 15691 13504 15700
rect 1216 15512 1268 15564
rect 4160 15512 4212 15564
rect 2964 15444 3016 15496
rect 2872 15376 2924 15428
rect 6092 15580 6144 15632
rect 4528 15555 4580 15564
rect 4528 15521 4537 15555
rect 4537 15521 4571 15555
rect 4571 15521 4580 15555
rect 4528 15512 4580 15521
rect 4620 15555 4672 15564
rect 4620 15521 4629 15555
rect 4629 15521 4663 15555
rect 4663 15521 4672 15555
rect 10968 15580 11020 15632
rect 11428 15580 11480 15632
rect 12072 15580 12124 15632
rect 4620 15512 4672 15521
rect 5264 15444 5316 15496
rect 5816 15487 5868 15496
rect 5816 15453 5825 15487
rect 5825 15453 5859 15487
rect 5859 15453 5868 15487
rect 5816 15444 5868 15453
rect 6460 15444 6512 15496
rect 7472 15512 7524 15564
rect 7104 15444 7156 15496
rect 3240 15376 3292 15428
rect 7012 15376 7064 15428
rect 7472 15376 7524 15428
rect 7840 15444 7892 15496
rect 8116 15444 8168 15496
rect 8668 15512 8720 15564
rect 8852 15512 8904 15564
rect 9312 15512 9364 15564
rect 11060 15512 11112 15564
rect 8852 15376 8904 15428
rect 3976 15308 4028 15360
rect 4160 15351 4212 15360
rect 4160 15317 4169 15351
rect 4169 15317 4203 15351
rect 4203 15317 4212 15351
rect 4160 15308 4212 15317
rect 6552 15351 6604 15360
rect 6552 15317 6561 15351
rect 6561 15317 6595 15351
rect 6595 15317 6604 15351
rect 6552 15308 6604 15317
rect 7564 15308 7616 15360
rect 8116 15308 8168 15360
rect 10416 15444 10468 15496
rect 10876 15444 10928 15496
rect 11888 15444 11940 15496
rect 12440 15555 12492 15564
rect 12440 15521 12449 15555
rect 12449 15521 12483 15555
rect 12483 15521 12492 15555
rect 12440 15512 12492 15521
rect 12532 15487 12584 15496
rect 12532 15453 12541 15487
rect 12541 15453 12575 15487
rect 12575 15453 12584 15487
rect 12532 15444 12584 15453
rect 12808 15512 12860 15564
rect 13452 15657 13461 15691
rect 13461 15657 13495 15691
rect 13495 15657 13504 15691
rect 13452 15648 13504 15657
rect 14188 15691 14240 15700
rect 14188 15657 14197 15691
rect 14197 15657 14231 15691
rect 14231 15657 14240 15691
rect 14188 15648 14240 15657
rect 14096 15512 14148 15564
rect 15292 15444 15344 15496
rect 9220 15376 9272 15428
rect 9680 15376 9732 15428
rect 10048 15376 10100 15428
rect 10968 15376 11020 15428
rect 12348 15376 12400 15428
rect 9128 15308 9180 15360
rect 12072 15351 12124 15360
rect 12072 15317 12081 15351
rect 12081 15317 12115 15351
rect 12115 15317 12124 15351
rect 12072 15308 12124 15317
rect 3447 15206 3499 15258
rect 3511 15206 3563 15258
rect 3575 15206 3627 15258
rect 3639 15206 3691 15258
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 13308 15206 13360 15258
rect 13372 15206 13424 15258
rect 13436 15206 13488 15258
rect 13500 15206 13552 15258
rect 2504 15104 2556 15156
rect 4344 15104 4396 15156
rect 3884 15036 3936 15088
rect 2872 14968 2924 15020
rect 3792 15011 3844 15020
rect 3792 14977 3801 15011
rect 3801 14977 3835 15011
rect 3835 14977 3844 15011
rect 3792 14968 3844 14977
rect 5356 15104 5408 15156
rect 5816 15104 5868 15156
rect 7380 15104 7432 15156
rect 9588 15104 9640 15156
rect 10692 15104 10744 15156
rect 4712 15036 4764 15088
rect 8944 15036 8996 15088
rect 9864 15079 9916 15088
rect 4988 15011 5040 15020
rect 1676 14832 1728 14884
rect 2688 14832 2740 14884
rect 2780 14832 2832 14884
rect 1768 14764 1820 14816
rect 2872 14764 2924 14816
rect 4988 14977 4997 15011
rect 4997 14977 5031 15011
rect 5031 14977 5040 15011
rect 4988 14968 5040 14977
rect 5356 14968 5408 15020
rect 4068 14900 4120 14952
rect 4620 14900 4672 14952
rect 4344 14807 4396 14816
rect 4344 14773 4353 14807
rect 4353 14773 4387 14807
rect 4387 14773 4396 14807
rect 4344 14764 4396 14773
rect 4804 14807 4856 14816
rect 4804 14773 4813 14807
rect 4813 14773 4847 14807
rect 4847 14773 4856 14807
rect 4804 14764 4856 14773
rect 5632 14900 5684 14952
rect 5816 14968 5868 15020
rect 6092 15011 6144 15020
rect 6092 14977 6101 15011
rect 6101 14977 6135 15011
rect 6135 14977 6144 15011
rect 6092 14968 6144 14977
rect 7564 14968 7616 15020
rect 7932 14968 7984 15020
rect 9220 15011 9272 15020
rect 9220 14977 9229 15011
rect 9229 14977 9263 15011
rect 9263 14977 9272 15011
rect 9220 14968 9272 14977
rect 9864 15045 9873 15079
rect 9873 15045 9907 15079
rect 9907 15045 9916 15079
rect 9864 15036 9916 15045
rect 10048 15036 10100 15088
rect 13084 15036 13136 15088
rect 13820 15036 13872 15088
rect 11888 14968 11940 15020
rect 6368 14900 6420 14952
rect 7748 14900 7800 14952
rect 8484 14900 8536 14952
rect 6920 14832 6972 14884
rect 10876 14900 10928 14952
rect 12072 14900 12124 14952
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 13084 14900 13136 14952
rect 15200 14900 15252 14952
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 8024 14807 8076 14816
rect 8024 14773 8033 14807
rect 8033 14773 8067 14807
rect 8067 14773 8076 14807
rect 8024 14764 8076 14773
rect 8668 14807 8720 14816
rect 8668 14773 8677 14807
rect 8677 14773 8711 14807
rect 8711 14773 8720 14807
rect 8668 14764 8720 14773
rect 8852 14764 8904 14816
rect 14464 14832 14516 14884
rect 10140 14764 10192 14816
rect 11520 14764 11572 14816
rect 5912 14662 5964 14714
rect 5976 14662 6028 14714
rect 6040 14662 6092 14714
rect 6104 14662 6156 14714
rect 10843 14662 10895 14714
rect 10907 14662 10959 14714
rect 10971 14662 11023 14714
rect 11035 14662 11087 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 2688 14560 2740 14612
rect 3240 14560 3292 14612
rect 4252 14560 4304 14612
rect 6552 14492 6604 14544
rect 7288 14560 7340 14612
rect 12348 14560 12400 14612
rect 10508 14492 10560 14544
rect 13084 14492 13136 14544
rect 13176 14492 13228 14544
rect 14924 14492 14976 14544
rect 3148 14467 3200 14476
rect 3148 14433 3157 14467
rect 3157 14433 3191 14467
rect 3191 14433 3200 14467
rect 3148 14424 3200 14433
rect 4712 14424 4764 14476
rect 2044 14399 2096 14408
rect 2044 14365 2053 14399
rect 2053 14365 2087 14399
rect 2087 14365 2096 14399
rect 2044 14356 2096 14365
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 3240 14399 3292 14408
rect 2136 14356 2188 14365
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 4436 14356 4488 14408
rect 5908 14424 5960 14476
rect 7840 14424 7892 14476
rect 8208 14424 8260 14476
rect 9312 14424 9364 14476
rect 3792 14288 3844 14340
rect 4896 14356 4948 14408
rect 5356 14399 5408 14408
rect 5356 14365 5365 14399
rect 5365 14365 5399 14399
rect 5399 14365 5408 14399
rect 5356 14356 5408 14365
rect 6828 14356 6880 14408
rect 9772 14356 9824 14408
rect 10140 14399 10192 14408
rect 10140 14365 10149 14399
rect 10149 14365 10183 14399
rect 10183 14365 10192 14399
rect 10140 14356 10192 14365
rect 8576 14331 8628 14340
rect 6736 14263 6788 14272
rect 6736 14229 6745 14263
rect 6745 14229 6779 14263
rect 6779 14229 6788 14263
rect 6736 14220 6788 14229
rect 7012 14220 7064 14272
rect 8576 14297 8585 14331
rect 8585 14297 8619 14331
rect 8619 14297 8628 14331
rect 8576 14288 8628 14297
rect 9680 14331 9732 14340
rect 9680 14297 9689 14331
rect 9689 14297 9723 14331
rect 9723 14297 9732 14331
rect 9680 14288 9732 14297
rect 10048 14288 10100 14340
rect 8208 14220 8260 14272
rect 8944 14220 8996 14272
rect 9864 14220 9916 14272
rect 11060 14424 11112 14476
rect 11612 14424 11664 14476
rect 12716 14424 12768 14476
rect 13544 14424 13596 14476
rect 11888 14356 11940 14408
rect 12348 14356 12400 14408
rect 13820 14399 13872 14408
rect 13820 14365 13829 14399
rect 13829 14365 13863 14399
rect 13863 14365 13872 14399
rect 13820 14356 13872 14365
rect 13176 14220 13228 14272
rect 3447 14118 3499 14170
rect 3511 14118 3563 14170
rect 3575 14118 3627 14170
rect 3639 14118 3691 14170
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 13308 14118 13360 14170
rect 13372 14118 13424 14170
rect 13436 14118 13488 14170
rect 13500 14118 13552 14170
rect 2504 14059 2556 14068
rect 2504 14025 2513 14059
rect 2513 14025 2547 14059
rect 2547 14025 2556 14059
rect 2504 14016 2556 14025
rect 4068 14016 4120 14068
rect 2596 13948 2648 14000
rect 6644 13948 6696 14000
rect 8116 13948 8168 14000
rect 8576 13948 8628 14000
rect 3792 13880 3844 13932
rect 4160 13923 4212 13932
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 2872 13812 2924 13864
rect 4252 13812 4304 13864
rect 4896 13855 4948 13864
rect 4896 13821 4905 13855
rect 4905 13821 4939 13855
rect 4939 13821 4948 13855
rect 4896 13812 4948 13821
rect 6368 13880 6420 13932
rect 6552 13880 6604 13932
rect 8484 13880 8536 13932
rect 9312 14016 9364 14068
rect 9404 14016 9456 14068
rect 10508 14059 10560 14068
rect 10508 14025 10517 14059
rect 10517 14025 10551 14059
rect 10551 14025 10560 14059
rect 10508 14016 10560 14025
rect 9956 13948 10008 14000
rect 10140 13948 10192 14000
rect 13820 14016 13872 14068
rect 12716 13948 12768 14000
rect 13360 13948 13412 14000
rect 11336 13880 11388 13932
rect 11612 13880 11664 13932
rect 6276 13812 6328 13864
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 6368 13744 6420 13796
rect 6460 13744 6512 13796
rect 7380 13744 7432 13796
rect 7748 13744 7800 13796
rect 9680 13812 9732 13864
rect 9956 13812 10008 13864
rect 10048 13812 10100 13864
rect 10692 13812 10744 13864
rect 11888 13855 11940 13864
rect 11888 13821 11897 13855
rect 11897 13821 11931 13855
rect 11931 13821 11940 13855
rect 11888 13812 11940 13821
rect 12348 13880 12400 13932
rect 13268 13812 13320 13864
rect 15568 13880 15620 13932
rect 13636 13812 13688 13864
rect 9312 13744 9364 13796
rect 9588 13744 9640 13796
rect 12256 13744 12308 13796
rect 2320 13676 2372 13728
rect 9956 13676 10008 13728
rect 10692 13676 10744 13728
rect 16396 13744 16448 13796
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 13820 13676 13872 13728
rect 5912 13574 5964 13626
rect 5976 13574 6028 13626
rect 6040 13574 6092 13626
rect 6104 13574 6156 13626
rect 10843 13574 10895 13626
rect 10907 13574 10959 13626
rect 10971 13574 11023 13626
rect 11035 13574 11087 13626
rect 2228 13404 2280 13456
rect 4620 13472 4672 13524
rect 5080 13472 5132 13524
rect 5356 13472 5408 13524
rect 6368 13515 6420 13524
rect 6368 13481 6377 13515
rect 6377 13481 6411 13515
rect 6411 13481 6420 13515
rect 6368 13472 6420 13481
rect 6920 13472 6972 13524
rect 7104 13472 7156 13524
rect 7840 13472 7892 13524
rect 8208 13515 8260 13524
rect 8208 13481 8217 13515
rect 8217 13481 8251 13515
rect 8251 13481 8260 13515
rect 8208 13472 8260 13481
rect 9496 13472 9548 13524
rect 10508 13472 10560 13524
rect 11980 13472 12032 13524
rect 12256 13472 12308 13524
rect 3792 13404 3844 13456
rect 2504 13336 2556 13388
rect 2688 13336 2740 13388
rect 12624 13404 12676 13456
rect 4620 13336 4672 13388
rect 7104 13379 7156 13388
rect 7104 13345 7138 13379
rect 7138 13345 7156 13379
rect 7104 13336 7156 13345
rect 8300 13336 8352 13388
rect 9588 13336 9640 13388
rect 9772 13336 9824 13388
rect 10508 13336 10560 13388
rect 1492 13268 1544 13320
rect 4252 13311 4304 13320
rect 2412 13200 2464 13252
rect 2780 13243 2832 13252
rect 2780 13209 2789 13243
rect 2789 13209 2823 13243
rect 2823 13209 2832 13243
rect 2780 13200 2832 13209
rect 1860 13132 1912 13184
rect 3240 13132 3292 13184
rect 4252 13277 4261 13311
rect 4261 13277 4295 13311
rect 4295 13277 4304 13311
rect 4252 13268 4304 13277
rect 4896 13268 4948 13320
rect 6828 13311 6880 13320
rect 6828 13277 6837 13311
rect 6837 13277 6871 13311
rect 6871 13277 6880 13311
rect 6828 13268 6880 13277
rect 8852 13311 8904 13320
rect 8852 13277 8861 13311
rect 8861 13277 8895 13311
rect 8895 13277 8904 13311
rect 8852 13268 8904 13277
rect 11520 13336 11572 13388
rect 13912 13472 13964 13524
rect 14832 13472 14884 13524
rect 13820 13447 13872 13456
rect 13820 13413 13829 13447
rect 13829 13413 13863 13447
rect 13863 13413 13872 13447
rect 13820 13404 13872 13413
rect 13268 13336 13320 13388
rect 12348 13268 12400 13320
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 14004 13311 14056 13320
rect 14004 13277 14013 13311
rect 14013 13277 14047 13311
rect 14047 13277 14056 13311
rect 14004 13268 14056 13277
rect 7840 13200 7892 13252
rect 9680 13200 9732 13252
rect 11060 13243 11112 13252
rect 11060 13209 11069 13243
rect 11069 13209 11103 13243
rect 11103 13209 11112 13243
rect 11060 13200 11112 13209
rect 6644 13132 6696 13184
rect 7196 13132 7248 13184
rect 13820 13200 13872 13252
rect 11520 13175 11572 13184
rect 11520 13141 11529 13175
rect 11529 13141 11563 13175
rect 11563 13141 11572 13175
rect 11520 13132 11572 13141
rect 3447 13030 3499 13082
rect 3511 13030 3563 13082
rect 3575 13030 3627 13082
rect 3639 13030 3691 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 13308 13030 13360 13082
rect 13372 13030 13424 13082
rect 13436 13030 13488 13082
rect 13500 13030 13552 13082
rect 1860 12971 1912 12980
rect 1860 12937 1869 12971
rect 1869 12937 1903 12971
rect 1903 12937 1912 12971
rect 1860 12928 1912 12937
rect 2228 12928 2280 12980
rect 4160 12928 4212 12980
rect 4436 12971 4488 12980
rect 4436 12937 4445 12971
rect 4445 12937 4479 12971
rect 4479 12937 4488 12971
rect 4436 12928 4488 12937
rect 4528 12928 4580 12980
rect 3056 12835 3108 12844
rect 3056 12801 3065 12835
rect 3065 12801 3099 12835
rect 3099 12801 3108 12835
rect 3056 12792 3108 12801
rect 4712 12792 4764 12844
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 4436 12724 4488 12776
rect 5448 12724 5500 12776
rect 9128 12928 9180 12980
rect 9588 12928 9640 12980
rect 7656 12860 7708 12912
rect 8300 12860 8352 12912
rect 8392 12860 8444 12912
rect 9772 12860 9824 12912
rect 9956 12928 10008 12980
rect 11060 12928 11112 12980
rect 12992 12928 13044 12980
rect 13084 12928 13136 12980
rect 12624 12860 12676 12912
rect 7840 12792 7892 12844
rect 7932 12792 7984 12844
rect 9036 12835 9088 12844
rect 7380 12724 7432 12776
rect 8392 12767 8444 12776
rect 8392 12733 8401 12767
rect 8401 12733 8435 12767
rect 8435 12733 8444 12767
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 10876 12792 10928 12844
rect 11520 12792 11572 12844
rect 13820 12792 13872 12844
rect 8392 12724 8444 12733
rect 9588 12724 9640 12776
rect 9680 12724 9732 12776
rect 10600 12724 10652 12776
rect 3424 12656 3476 12708
rect 3792 12656 3844 12708
rect 7932 12656 7984 12708
rect 1952 12588 2004 12640
rect 4344 12588 4396 12640
rect 5724 12588 5776 12640
rect 6920 12588 6972 12640
rect 8944 12656 8996 12708
rect 8208 12588 8260 12640
rect 9220 12588 9272 12640
rect 9772 12588 9824 12640
rect 9956 12588 10008 12640
rect 10692 12656 10744 12708
rect 12072 12724 12124 12776
rect 12348 12724 12400 12776
rect 12440 12724 12492 12776
rect 13636 12656 13688 12708
rect 11520 12588 11572 12640
rect 13084 12588 13136 12640
rect 5912 12486 5964 12538
rect 5976 12486 6028 12538
rect 6040 12486 6092 12538
rect 6104 12486 6156 12538
rect 10843 12486 10895 12538
rect 10907 12486 10959 12538
rect 10971 12486 11023 12538
rect 11035 12486 11087 12538
rect 1584 12384 1636 12436
rect 5724 12384 5776 12436
rect 6460 12384 6512 12436
rect 6368 12316 6420 12368
rect 6920 12384 6972 12436
rect 7196 12384 7248 12436
rect 7380 12384 7432 12436
rect 8484 12384 8536 12436
rect 8852 12384 8904 12436
rect 2688 12291 2740 12300
rect 2688 12257 2697 12291
rect 2697 12257 2731 12291
rect 2731 12257 2740 12291
rect 2688 12248 2740 12257
rect 4712 12291 4764 12300
rect 4712 12257 4721 12291
rect 4721 12257 4755 12291
rect 4755 12257 4764 12291
rect 4712 12248 4764 12257
rect 5264 12248 5316 12300
rect 8208 12316 8260 12368
rect 8668 12359 8720 12368
rect 8668 12325 8677 12359
rect 8677 12325 8711 12359
rect 8711 12325 8720 12359
rect 9312 12384 9364 12436
rect 10048 12384 10100 12436
rect 10692 12384 10744 12436
rect 15200 12384 15252 12436
rect 8668 12316 8720 12325
rect 9220 12316 9272 12368
rect 6736 12291 6788 12300
rect 6736 12257 6745 12291
rect 6745 12257 6779 12291
rect 6779 12257 6788 12291
rect 6736 12248 6788 12257
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 6552 12180 6604 12232
rect 8576 12248 8628 12300
rect 8760 12248 8812 12300
rect 9772 12248 9824 12300
rect 10048 12248 10100 12300
rect 10232 12248 10284 12300
rect 10968 12316 11020 12368
rect 11336 12291 11388 12300
rect 11336 12257 11345 12291
rect 11345 12257 11379 12291
rect 11379 12257 11388 12291
rect 11336 12248 11388 12257
rect 4160 12044 4212 12096
rect 7012 12044 7064 12096
rect 7472 12044 7524 12096
rect 7840 12180 7892 12232
rect 7748 12044 7800 12096
rect 8300 12180 8352 12232
rect 8024 12112 8076 12164
rect 8208 12044 8260 12096
rect 9128 12044 9180 12096
rect 11888 12248 11940 12300
rect 12164 12316 12216 12368
rect 13268 12316 13320 12368
rect 12808 12248 12860 12300
rect 14280 12248 14332 12300
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 12900 12180 12952 12232
rect 12256 12044 12308 12096
rect 12808 12112 12860 12164
rect 3447 11942 3499 11994
rect 3511 11942 3563 11994
rect 3575 11942 3627 11994
rect 3639 11942 3691 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 13308 11942 13360 11994
rect 13372 11942 13424 11994
rect 13436 11942 13488 11994
rect 13500 11942 13552 11994
rect 2320 11611 2372 11620
rect 2320 11577 2329 11611
rect 2329 11577 2363 11611
rect 2363 11577 2372 11611
rect 2320 11568 2372 11577
rect 2780 11704 2832 11756
rect 3240 11840 3292 11892
rect 7840 11840 7892 11892
rect 4712 11704 4764 11756
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 10508 11840 10560 11892
rect 10876 11840 10928 11892
rect 12716 11840 12768 11892
rect 9864 11772 9916 11824
rect 6644 11636 6696 11688
rect 3424 11568 3476 11620
rect 5356 11568 5408 11620
rect 5632 11568 5684 11620
rect 7196 11568 7248 11620
rect 2044 11500 2096 11552
rect 2688 11500 2740 11552
rect 4620 11500 4672 11552
rect 7104 11500 7156 11552
rect 8300 11636 8352 11688
rect 11612 11704 11664 11756
rect 14740 11704 14792 11756
rect 15476 11704 15528 11756
rect 10876 11679 10928 11688
rect 7656 11568 7708 11620
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 8484 11568 8536 11620
rect 9864 11568 9916 11620
rect 10876 11645 10885 11679
rect 10885 11645 10919 11679
rect 10919 11645 10928 11679
rect 10876 11636 10928 11645
rect 12440 11636 12492 11688
rect 14464 11636 14516 11688
rect 16396 11636 16448 11688
rect 10784 11568 10836 11620
rect 11428 11568 11480 11620
rect 12624 11568 12676 11620
rect 12716 11568 12768 11620
rect 12992 11568 13044 11620
rect 14740 11568 14792 11620
rect 13452 11500 13504 11552
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 14096 11543 14148 11552
rect 14096 11509 14105 11543
rect 14105 11509 14139 11543
rect 14139 11509 14148 11543
rect 15016 11543 15068 11552
rect 14096 11500 14148 11509
rect 15016 11509 15025 11543
rect 15025 11509 15059 11543
rect 15059 11509 15068 11543
rect 15016 11500 15068 11509
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 6104 11398 6156 11450
rect 10843 11398 10895 11450
rect 10907 11398 10959 11450
rect 10971 11398 11023 11450
rect 11035 11398 11087 11450
rect 11336 11296 11388 11348
rect 11520 11339 11572 11348
rect 11520 11305 11529 11339
rect 11529 11305 11563 11339
rect 11563 11305 11572 11339
rect 11520 11296 11572 11305
rect 11704 11296 11756 11348
rect 12532 11296 12584 11348
rect 12808 11296 12860 11348
rect 12992 11296 13044 11348
rect 14096 11296 14148 11348
rect 1860 11271 1912 11280
rect 1860 11237 1869 11271
rect 1869 11237 1903 11271
rect 1903 11237 1912 11271
rect 1860 11228 1912 11237
rect 2780 11228 2832 11280
rect 4896 11228 4948 11280
rect 4712 11160 4764 11212
rect 6552 11160 6604 11212
rect 7380 11228 7432 11280
rect 8208 11228 8260 11280
rect 9404 11228 9456 11280
rect 10508 11228 10560 11280
rect 10784 11228 10836 11280
rect 13176 11228 13228 11280
rect 11520 11160 11572 11212
rect 6828 11092 6880 11144
rect 8760 11135 8812 11144
rect 8760 11101 8769 11135
rect 8769 11101 8803 11135
rect 8803 11101 8812 11135
rect 8760 11092 8812 11101
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 10692 11092 10744 11144
rect 11796 11092 11848 11144
rect 3240 11024 3292 11076
rect 3424 11024 3476 11076
rect 3792 11024 3844 11076
rect 4068 11024 4120 11076
rect 5080 11024 5132 11076
rect 5540 11024 5592 11076
rect 8024 11024 8076 11076
rect 9496 11024 9548 11076
rect 10784 11024 10836 11076
rect 12440 11160 12492 11212
rect 13084 11203 13136 11212
rect 13084 11169 13093 11203
rect 13093 11169 13127 11203
rect 13127 11169 13136 11203
rect 13084 11160 13136 11169
rect 12072 11135 12124 11144
rect 12072 11101 12081 11135
rect 12081 11101 12115 11135
rect 12115 11101 12124 11135
rect 12072 11092 12124 11101
rect 13544 11160 13596 11212
rect 14096 11160 14148 11212
rect 14280 11203 14332 11212
rect 14280 11169 14289 11203
rect 14289 11169 14323 11203
rect 14323 11169 14332 11203
rect 14280 11160 14332 11169
rect 13268 11135 13320 11144
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 14004 11024 14056 11076
rect 2504 10956 2556 11008
rect 4252 10956 4304 11008
rect 5356 10956 5408 11008
rect 14648 11092 14700 11144
rect 3447 10854 3499 10906
rect 3511 10854 3563 10906
rect 3575 10854 3627 10906
rect 3639 10854 3691 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 13308 10854 13360 10906
rect 13372 10854 13424 10906
rect 13436 10854 13488 10906
rect 13500 10854 13552 10906
rect 1308 10752 1360 10804
rect 2136 10752 2188 10804
rect 2228 10752 2280 10804
rect 6276 10795 6328 10804
rect 6276 10761 6285 10795
rect 6285 10761 6319 10795
rect 6319 10761 6328 10795
rect 6276 10752 6328 10761
rect 6552 10752 6604 10804
rect 11244 10752 11296 10804
rect 11704 10752 11756 10804
rect 12900 10752 12952 10804
rect 13636 10795 13688 10804
rect 13636 10761 13645 10795
rect 13645 10761 13679 10795
rect 13679 10761 13688 10795
rect 13636 10752 13688 10761
rect 13912 10752 13964 10804
rect 14096 10752 14148 10804
rect 4160 10684 4212 10736
rect 7932 10684 7984 10736
rect 11796 10684 11848 10736
rect 2504 10659 2556 10668
rect 2504 10625 2513 10659
rect 2513 10625 2547 10659
rect 2547 10625 2556 10659
rect 2504 10616 2556 10625
rect 4068 10616 4120 10668
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 9680 10616 9732 10668
rect 10140 10616 10192 10668
rect 11520 10616 11572 10668
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 2780 10548 2832 10600
rect 8024 10548 8076 10600
rect 8208 10548 8260 10600
rect 8300 10548 8352 10600
rect 1860 10480 1912 10532
rect 2228 10455 2280 10464
rect 2228 10421 2237 10455
rect 2237 10421 2271 10455
rect 2271 10421 2280 10455
rect 2228 10412 2280 10421
rect 5080 10480 5132 10532
rect 4344 10412 4396 10464
rect 4988 10412 5040 10464
rect 11612 10548 11664 10600
rect 11796 10548 11848 10600
rect 13452 10684 13504 10736
rect 14924 10684 14976 10736
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 13176 10616 13228 10668
rect 14096 10548 14148 10600
rect 14372 10548 14424 10600
rect 14556 10548 14608 10600
rect 5448 10412 5500 10464
rect 11152 10480 11204 10532
rect 13268 10480 13320 10532
rect 13912 10480 13964 10532
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 11520 10412 11572 10464
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 12900 10412 12952 10464
rect 13084 10412 13136 10464
rect 15016 10455 15068 10464
rect 15016 10421 15025 10455
rect 15025 10421 15059 10455
rect 15059 10421 15068 10455
rect 15016 10412 15068 10421
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 6104 10310 6156 10362
rect 10843 10310 10895 10362
rect 10907 10310 10959 10362
rect 10971 10310 11023 10362
rect 11035 10310 11087 10362
rect 2412 10183 2464 10192
rect 2412 10149 2446 10183
rect 2446 10149 2464 10183
rect 2412 10140 2464 10149
rect 4620 10208 4672 10260
rect 4436 10140 4488 10192
rect 5448 10140 5500 10192
rect 2780 10072 2832 10124
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 5816 10208 5868 10260
rect 6552 10208 6604 10260
rect 7380 10208 7432 10260
rect 7748 10208 7800 10260
rect 8208 10208 8260 10260
rect 8852 10208 8904 10260
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 9312 10208 9364 10260
rect 9496 10208 9548 10260
rect 10508 10208 10560 10260
rect 11612 10208 11664 10260
rect 12164 10208 12216 10260
rect 12440 10208 12492 10260
rect 13820 10208 13872 10260
rect 6276 10140 6328 10192
rect 7840 10140 7892 10192
rect 8116 10140 8168 10192
rect 5264 10004 5316 10056
rect 8300 10072 8352 10124
rect 3424 9936 3476 9988
rect 5356 9936 5408 9988
rect 4252 9868 4304 9920
rect 10508 10072 10560 10124
rect 8852 10004 8904 10056
rect 9312 10004 9364 10056
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 10784 9936 10836 9988
rect 11152 9936 11204 9988
rect 11520 10072 11572 10124
rect 11704 10004 11756 10056
rect 12440 10072 12492 10124
rect 13084 10115 13136 10124
rect 13084 10081 13093 10115
rect 13093 10081 13127 10115
rect 13127 10081 13136 10115
rect 13084 10072 13136 10081
rect 13636 10072 13688 10124
rect 13820 10072 13872 10124
rect 12440 9936 12492 9988
rect 8852 9868 8904 9920
rect 9036 9868 9088 9920
rect 9220 9868 9272 9920
rect 12164 9868 12216 9920
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 14464 10047 14516 10056
rect 14464 10013 14473 10047
rect 14473 10013 14507 10047
rect 14507 10013 14516 10047
rect 14464 10004 14516 10013
rect 13912 9868 13964 9920
rect 3447 9766 3499 9818
rect 3511 9766 3563 9818
rect 3575 9766 3627 9818
rect 3639 9766 3691 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 13308 9766 13360 9818
rect 13372 9766 13424 9818
rect 13436 9766 13488 9818
rect 13500 9766 13552 9818
rect 1860 9707 1912 9716
rect 1860 9673 1869 9707
rect 1869 9673 1903 9707
rect 1903 9673 1912 9707
rect 1860 9664 1912 9673
rect 4436 9707 4488 9716
rect 4436 9673 4445 9707
rect 4445 9673 4479 9707
rect 4479 9673 4488 9707
rect 4436 9664 4488 9673
rect 4160 9596 4212 9648
rect 6552 9664 6604 9716
rect 10048 9664 10100 9716
rect 11152 9664 11204 9716
rect 11612 9664 11664 9716
rect 11888 9664 11940 9716
rect 12164 9664 12216 9716
rect 13084 9664 13136 9716
rect 7288 9596 7340 9648
rect 8024 9596 8076 9648
rect 9036 9596 9088 9648
rect 5080 9528 5132 9580
rect 5264 9571 5316 9580
rect 5264 9537 5273 9571
rect 5273 9537 5307 9571
rect 5307 9537 5316 9571
rect 5264 9528 5316 9537
rect 6276 9528 6328 9580
rect 7104 9528 7156 9580
rect 7748 9528 7800 9580
rect 2136 9460 2188 9512
rect 2872 9460 2924 9512
rect 6736 9460 6788 9512
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 10048 9528 10100 9580
rect 9588 9460 9640 9512
rect 9680 9460 9732 9512
rect 11612 9460 11664 9512
rect 2688 9392 2740 9444
rect 4988 9392 5040 9444
rect 6828 9392 6880 9444
rect 7012 9392 7064 9444
rect 7288 9392 7340 9444
rect 8392 9392 8444 9444
rect 9404 9392 9456 9444
rect 10600 9392 10652 9444
rect 11520 9392 11572 9444
rect 2320 9367 2372 9376
rect 2320 9333 2329 9367
rect 2329 9333 2363 9367
rect 2363 9333 2372 9367
rect 2320 9324 2372 9333
rect 2596 9324 2648 9376
rect 6644 9367 6696 9376
rect 6644 9333 6653 9367
rect 6653 9333 6687 9367
rect 6687 9333 6696 9367
rect 6644 9324 6696 9333
rect 6920 9324 6972 9376
rect 9680 9324 9732 9376
rect 9956 9324 10008 9376
rect 13636 9596 13688 9648
rect 15384 9596 15436 9648
rect 12992 9528 13044 9580
rect 12624 9460 12676 9512
rect 13268 9460 13320 9512
rect 14004 9460 14056 9512
rect 14924 9460 14976 9512
rect 12440 9392 12492 9444
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 11980 9324 12032 9376
rect 12992 9324 13044 9376
rect 13636 9367 13688 9376
rect 13636 9333 13645 9367
rect 13645 9333 13679 9367
rect 13679 9333 13688 9367
rect 13636 9324 13688 9333
rect 14004 9367 14056 9376
rect 14004 9333 14013 9367
rect 14013 9333 14047 9367
rect 14047 9333 14056 9367
rect 14004 9324 14056 9333
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 6104 9222 6156 9274
rect 10843 9222 10895 9274
rect 10907 9222 10959 9274
rect 10971 9222 11023 9274
rect 11035 9222 11087 9274
rect 2320 9120 2372 9172
rect 9220 9120 9272 9172
rect 9588 9120 9640 9172
rect 14004 9120 14056 9172
rect 15108 9120 15160 9172
rect 5080 9052 5132 9104
rect 11888 9052 11940 9104
rect 1308 8916 1360 8968
rect 1584 8916 1636 8968
rect 1216 8780 1268 8832
rect 2136 9027 2188 9036
rect 2136 8993 2145 9027
rect 2145 8993 2179 9027
rect 2179 8993 2188 9027
rect 2136 8984 2188 8993
rect 4344 8984 4396 9036
rect 5356 8984 5408 9036
rect 5816 8984 5868 9036
rect 7012 8984 7064 9036
rect 7104 8984 7156 9036
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 3516 8891 3568 8900
rect 3516 8857 3525 8891
rect 3525 8857 3559 8891
rect 3559 8857 3568 8891
rect 3516 8848 3568 8857
rect 5632 8891 5684 8900
rect 5632 8857 5641 8891
rect 5641 8857 5675 8891
rect 5675 8857 5684 8891
rect 5632 8848 5684 8857
rect 6828 8848 6880 8900
rect 7196 8848 7248 8900
rect 4252 8780 4304 8832
rect 4436 8780 4488 8832
rect 6920 8780 6972 8832
rect 7104 8823 7156 8832
rect 7104 8789 7113 8823
rect 7113 8789 7147 8823
rect 7147 8789 7156 8823
rect 7104 8780 7156 8789
rect 8760 8984 8812 9036
rect 9404 8984 9456 9036
rect 13176 9052 13228 9104
rect 9036 8916 9088 8968
rect 9680 8959 9732 8968
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 11428 8916 11480 8968
rect 12532 8916 12584 8968
rect 12716 8916 12768 8968
rect 13176 8916 13228 8968
rect 13820 8916 13872 8968
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 8576 8848 8628 8900
rect 9220 8848 9272 8900
rect 9496 8848 9548 8900
rect 7932 8780 7984 8832
rect 8668 8780 8720 8832
rect 9036 8780 9088 8832
rect 9128 8780 9180 8832
rect 9956 8780 10008 8832
rect 11244 8780 11296 8832
rect 11336 8780 11388 8832
rect 13084 8848 13136 8900
rect 13360 8891 13412 8900
rect 13360 8857 13369 8891
rect 13369 8857 13403 8891
rect 13403 8857 13412 8891
rect 13360 8848 13412 8857
rect 14188 8780 14240 8832
rect 3447 8678 3499 8730
rect 3511 8678 3563 8730
rect 3575 8678 3627 8730
rect 3639 8678 3691 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 13308 8678 13360 8730
rect 13372 8678 13424 8730
rect 13436 8678 13488 8730
rect 13500 8678 13552 8730
rect 2596 8440 2648 8492
rect 2872 8440 2924 8492
rect 4344 8576 4396 8628
rect 4436 8551 4488 8560
rect 4436 8517 4445 8551
rect 4445 8517 4479 8551
rect 4479 8517 4488 8551
rect 4436 8508 4488 8517
rect 7840 8576 7892 8628
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 13636 8619 13688 8628
rect 12440 8576 12492 8585
rect 13636 8585 13645 8619
rect 13645 8585 13679 8619
rect 13679 8585 13688 8619
rect 13636 8576 13688 8585
rect 10048 8551 10100 8560
rect 1952 8415 2004 8424
rect 1952 8381 1961 8415
rect 1961 8381 1995 8415
rect 1995 8381 2004 8415
rect 1952 8372 2004 8381
rect 4160 8372 4212 8424
rect 4528 8372 4580 8424
rect 4896 8415 4948 8424
rect 4896 8381 4905 8415
rect 4905 8381 4939 8415
rect 4939 8381 4948 8415
rect 4896 8372 4948 8381
rect 6000 8440 6052 8492
rect 6368 8440 6420 8492
rect 10048 8517 10057 8551
rect 10057 8517 10091 8551
rect 10091 8517 10100 8551
rect 10048 8508 10100 8517
rect 11612 8508 11664 8560
rect 12716 8508 12768 8560
rect 15016 8551 15068 8560
rect 15016 8517 15025 8551
rect 15025 8517 15059 8551
rect 15059 8517 15068 8551
rect 15016 8508 15068 8517
rect 3240 8304 3292 8356
rect 2320 8236 2372 8288
rect 4988 8304 5040 8356
rect 5540 8304 5592 8356
rect 5908 8372 5960 8424
rect 6828 8415 6880 8424
rect 6184 8304 6236 8356
rect 4252 8236 4304 8288
rect 6368 8236 6420 8288
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 8024 8440 8076 8492
rect 8392 8440 8444 8492
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 9772 8440 9824 8492
rect 9956 8440 10008 8492
rect 11520 8440 11572 8492
rect 13820 8440 13872 8492
rect 14464 8440 14516 8492
rect 9220 8372 9272 8424
rect 9680 8372 9732 8424
rect 12348 8372 12400 8424
rect 13084 8372 13136 8424
rect 7196 8304 7248 8356
rect 6920 8236 6972 8288
rect 7932 8236 7984 8288
rect 8208 8304 8260 8356
rect 10600 8304 10652 8356
rect 10692 8304 10744 8356
rect 11428 8304 11480 8356
rect 13820 8304 13872 8356
rect 8760 8236 8812 8288
rect 9036 8236 9088 8288
rect 11612 8236 11664 8288
rect 12164 8236 12216 8288
rect 12348 8236 12400 8288
rect 14004 8279 14056 8288
rect 14004 8245 14013 8279
rect 14013 8245 14047 8279
rect 14047 8245 14056 8279
rect 14004 8236 14056 8245
rect 15476 8372 15528 8424
rect 14464 8236 14516 8288
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 6104 8134 6156 8186
rect 10843 8134 10895 8186
rect 10907 8134 10959 8186
rect 10971 8134 11023 8186
rect 11035 8134 11087 8186
rect 5080 7964 5132 8016
rect 2688 7896 2740 7948
rect 5632 7896 5684 7948
rect 6368 8032 6420 8084
rect 6920 8032 6972 8084
rect 6000 8007 6052 8016
rect 6000 7973 6034 8007
rect 6034 7973 6052 8007
rect 6000 7964 6052 7973
rect 6736 7964 6788 8016
rect 7748 8032 7800 8084
rect 8208 8032 8260 8084
rect 8392 8032 8444 8084
rect 11796 8032 11848 8084
rect 14004 8032 14056 8084
rect 8668 8007 8720 8016
rect 1492 7692 1544 7744
rect 5264 7828 5316 7880
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 6920 7896 6972 7948
rect 8668 7973 8677 8007
rect 8677 7973 8711 8007
rect 8711 7973 8720 8007
rect 8668 7964 8720 7973
rect 7748 7896 7800 7948
rect 8024 7896 8076 7948
rect 8852 7871 8904 7880
rect 4252 7760 4304 7812
rect 2872 7692 2924 7744
rect 4528 7735 4580 7744
rect 4528 7701 4537 7735
rect 4537 7701 4571 7735
rect 4571 7701 4580 7735
rect 4528 7692 4580 7701
rect 8024 7760 8076 7812
rect 8852 7837 8861 7871
rect 8861 7837 8895 7871
rect 8895 7837 8904 7871
rect 8852 7828 8904 7837
rect 9588 7896 9640 7948
rect 10324 7896 10376 7948
rect 10876 7896 10928 7948
rect 11980 7939 12032 7948
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 12900 7896 12952 7948
rect 10968 7828 11020 7880
rect 11520 7828 11572 7880
rect 12072 7871 12124 7880
rect 12072 7837 12081 7871
rect 12081 7837 12115 7871
rect 12115 7837 12124 7871
rect 12072 7828 12124 7837
rect 12164 7828 12216 7880
rect 13728 7896 13780 7948
rect 14280 7828 14332 7880
rect 8668 7692 8720 7744
rect 8760 7692 8812 7744
rect 9036 7692 9088 7744
rect 10048 7692 10100 7744
rect 14188 7760 14240 7812
rect 10784 7692 10836 7744
rect 12532 7692 12584 7744
rect 3447 7590 3499 7642
rect 3511 7590 3563 7642
rect 3575 7590 3627 7642
rect 3639 7590 3691 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 13308 7590 13360 7642
rect 13372 7590 13424 7642
rect 13436 7590 13488 7642
rect 13500 7590 13552 7642
rect 2872 7488 2924 7540
rect 3240 7488 3292 7540
rect 5264 7488 5316 7540
rect 5632 7488 5684 7540
rect 7564 7488 7616 7540
rect 7840 7488 7892 7540
rect 5908 7420 5960 7472
rect 2596 7352 2648 7404
rect 2872 7352 2924 7404
rect 3056 7395 3108 7404
rect 3056 7361 3065 7395
rect 3065 7361 3099 7395
rect 3099 7361 3108 7395
rect 3056 7352 3108 7361
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 8300 7420 8352 7472
rect 9588 7488 9640 7540
rect 9956 7488 10008 7540
rect 1124 7284 1176 7336
rect 3792 7284 3844 7336
rect 4620 7216 4672 7268
rect 5356 7216 5408 7268
rect 5632 7284 5684 7336
rect 6644 7284 6696 7336
rect 6835 7327 6887 7336
rect 6835 7293 6844 7327
rect 6844 7293 6878 7327
rect 6878 7293 6887 7327
rect 6835 7284 6887 7293
rect 8392 7284 8444 7336
rect 9404 7284 9456 7336
rect 2228 7191 2280 7200
rect 2228 7157 2237 7191
rect 2237 7157 2271 7191
rect 2271 7157 2280 7191
rect 2228 7148 2280 7157
rect 5632 7148 5684 7200
rect 6276 7191 6328 7200
rect 6276 7157 6285 7191
rect 6285 7157 6319 7191
rect 6319 7157 6328 7191
rect 6276 7148 6328 7157
rect 7380 7216 7432 7268
rect 7564 7216 7616 7268
rect 8668 7216 8720 7268
rect 9036 7216 9088 7268
rect 9128 7216 9180 7268
rect 9588 7216 9640 7268
rect 7932 7148 7984 7200
rect 10968 7420 11020 7472
rect 11980 7488 12032 7540
rect 14372 7488 14424 7540
rect 9956 7352 10008 7404
rect 10784 7352 10836 7404
rect 13084 7420 13136 7472
rect 11336 7284 11388 7336
rect 10784 7216 10836 7268
rect 11060 7216 11112 7268
rect 11980 7352 12032 7404
rect 12072 7352 12124 7404
rect 14188 7395 14240 7404
rect 11612 7284 11664 7336
rect 12072 7216 12124 7268
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 14832 7327 14884 7336
rect 14832 7293 14841 7327
rect 14841 7293 14875 7327
rect 14875 7293 14884 7327
rect 14832 7284 14884 7293
rect 13912 7216 13964 7268
rect 10140 7148 10192 7200
rect 10232 7148 10284 7200
rect 10600 7148 10652 7200
rect 11336 7148 11388 7200
rect 11428 7148 11480 7200
rect 11980 7148 12032 7200
rect 14004 7191 14056 7200
rect 14004 7157 14013 7191
rect 14013 7157 14047 7191
rect 14047 7157 14056 7191
rect 14004 7148 14056 7157
rect 14372 7148 14424 7200
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 6104 7046 6156 7098
rect 10843 7046 10895 7098
rect 10907 7046 10959 7098
rect 10971 7046 11023 7098
rect 11035 7046 11087 7098
rect 2228 6944 2280 6996
rect 6736 6944 6788 6996
rect 7196 6987 7248 6996
rect 7196 6953 7205 6987
rect 7205 6953 7239 6987
rect 7239 6953 7248 6987
rect 7196 6944 7248 6953
rect 7564 6944 7616 6996
rect 8116 6944 8168 6996
rect 8392 6944 8444 6996
rect 10416 6944 10468 6996
rect 10600 6944 10652 6996
rect 12164 6944 12216 6996
rect 12624 6944 12676 6996
rect 14188 6944 14240 6996
rect 1308 6808 1360 6860
rect 2596 6876 2648 6928
rect 10232 6876 10284 6928
rect 3792 6808 3844 6860
rect 4068 6808 4120 6860
rect 6920 6808 6972 6860
rect 9128 6808 9180 6860
rect 9404 6808 9456 6860
rect 11060 6876 11112 6928
rect 11612 6808 11664 6860
rect 12164 6808 12216 6860
rect 12716 6876 12768 6928
rect 12900 6808 12952 6860
rect 13636 6851 13688 6860
rect 13636 6817 13645 6851
rect 13645 6817 13679 6851
rect 13679 6817 13688 6851
rect 13636 6808 13688 6817
rect 14096 6808 14148 6860
rect 4988 6783 5040 6792
rect 4988 6749 4997 6783
rect 4997 6749 5031 6783
rect 5031 6749 5040 6783
rect 4988 6740 5040 6749
rect 5172 6783 5224 6792
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 5172 6740 5224 6749
rect 5632 6672 5684 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 4896 6604 4948 6656
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 7656 6783 7708 6792
rect 5816 6740 5868 6749
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 8668 6740 8720 6792
rect 6920 6672 6972 6724
rect 7104 6604 7156 6656
rect 8852 6672 8904 6724
rect 9772 6740 9824 6792
rect 9312 6672 9364 6724
rect 9680 6715 9732 6724
rect 9680 6681 9689 6715
rect 9689 6681 9723 6715
rect 9723 6681 9732 6715
rect 10048 6740 10100 6792
rect 10600 6740 10652 6792
rect 11704 6740 11756 6792
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 13912 6783 13964 6792
rect 13912 6749 13921 6783
rect 13921 6749 13955 6783
rect 13955 6749 13964 6783
rect 13912 6740 13964 6749
rect 9680 6672 9732 6681
rect 12256 6672 12308 6724
rect 12992 6672 13044 6724
rect 14004 6672 14056 6724
rect 11980 6604 12032 6656
rect 12808 6604 12860 6656
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 1860 6443 1912 6452
rect 1860 6409 1869 6443
rect 1869 6409 1903 6443
rect 1903 6409 1912 6443
rect 1860 6400 1912 6409
rect 3792 6400 3844 6452
rect 3056 6332 3108 6384
rect 5908 6332 5960 6384
rect 6276 6332 6328 6384
rect 7932 6400 7984 6452
rect 8392 6332 8444 6384
rect 8576 6332 8628 6384
rect 10232 6400 10284 6452
rect 13636 6400 13688 6452
rect 10324 6332 10376 6384
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 1768 6196 1820 6248
rect 2596 6128 2648 6180
rect 4436 6196 4488 6248
rect 4804 6196 4856 6248
rect 5724 6196 5776 6248
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 11060 6264 11112 6316
rect 12164 6332 12216 6384
rect 13268 6332 13320 6384
rect 14280 6332 14332 6384
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 12348 6264 12400 6316
rect 13084 6264 13136 6316
rect 7380 6196 7432 6248
rect 7564 6196 7616 6248
rect 7656 6196 7708 6248
rect 7840 6196 7892 6248
rect 6460 6128 6512 6180
rect 7748 6128 7800 6180
rect 9404 6196 9456 6248
rect 9956 6196 10008 6248
rect 10232 6196 10284 6248
rect 12624 6196 12676 6248
rect 12808 6239 12860 6248
rect 12808 6205 12817 6239
rect 12817 6205 12851 6239
rect 12851 6205 12860 6239
rect 12808 6196 12860 6205
rect 15292 6196 15344 6248
rect 4344 6060 4396 6112
rect 4436 6060 4488 6112
rect 5816 6060 5868 6112
rect 6368 6060 6420 6112
rect 7012 6060 7064 6112
rect 8484 6060 8536 6112
rect 8576 6060 8628 6112
rect 13084 6128 13136 6180
rect 13912 6128 13964 6180
rect 9220 6060 9272 6112
rect 9680 6060 9732 6112
rect 12624 6060 12676 6112
rect 13544 6060 13596 6112
rect 13728 6060 13780 6112
rect 14648 6060 14700 6112
rect 14832 6060 14884 6112
rect 15016 6103 15068 6112
rect 15016 6069 15025 6103
rect 15025 6069 15059 6103
rect 15059 6069 15068 6103
rect 15016 6060 15068 6069
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 1400 5899 1452 5908
rect 1400 5865 1409 5899
rect 1409 5865 1443 5899
rect 1443 5865 1452 5899
rect 1400 5856 1452 5865
rect 4436 5856 4488 5908
rect 4896 5899 4948 5908
rect 4896 5865 4905 5899
rect 4905 5865 4939 5899
rect 4939 5865 4948 5899
rect 4896 5856 4948 5865
rect 4988 5856 5040 5908
rect 11336 5856 11388 5908
rect 12624 5856 12676 5908
rect 14556 5856 14608 5908
rect 14648 5899 14700 5908
rect 14648 5865 14657 5899
rect 14657 5865 14691 5899
rect 14691 5865 14700 5899
rect 14648 5856 14700 5865
rect 1308 5788 1360 5840
rect 2044 5788 2096 5840
rect 2780 5788 2832 5840
rect 2412 5720 2464 5772
rect 5448 5788 5500 5840
rect 6276 5788 6328 5840
rect 7748 5720 7800 5772
rect 9772 5788 9824 5840
rect 10692 5788 10744 5840
rect 9220 5720 9272 5772
rect 9588 5720 9640 5772
rect 11980 5788 12032 5840
rect 1768 5652 1820 5704
rect 4620 5652 4672 5704
rect 4988 5695 5040 5704
rect 4988 5661 4997 5695
rect 4997 5661 5031 5695
rect 5031 5661 5040 5695
rect 4988 5652 5040 5661
rect 5448 5652 5500 5704
rect 5632 5652 5684 5704
rect 2228 5584 2280 5636
rect 5356 5584 5408 5636
rect 4436 5516 4488 5568
rect 4896 5516 4948 5568
rect 7380 5652 7432 5704
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 10324 5695 10376 5704
rect 6736 5584 6788 5636
rect 6000 5516 6052 5568
rect 6460 5516 6512 5568
rect 7012 5516 7064 5568
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 11704 5720 11756 5772
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 11980 5652 12032 5704
rect 12164 5652 12216 5704
rect 12348 5720 12400 5772
rect 14924 5788 14976 5840
rect 12992 5720 13044 5772
rect 12348 5584 12400 5636
rect 9036 5559 9088 5568
rect 9036 5525 9045 5559
rect 9045 5525 9079 5559
rect 9079 5525 9088 5559
rect 9036 5516 9088 5525
rect 9588 5516 9640 5568
rect 11244 5516 11296 5568
rect 11520 5516 11572 5568
rect 11704 5516 11756 5568
rect 14188 5720 14240 5772
rect 12716 5584 12768 5636
rect 13268 5652 13320 5704
rect 13084 5584 13136 5636
rect 13544 5584 13596 5636
rect 12992 5516 13044 5568
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 4804 5312 4856 5364
rect 3332 5244 3384 5296
rect 3608 5244 3660 5296
rect 6092 5312 6144 5364
rect 7564 5312 7616 5364
rect 7656 5312 7708 5364
rect 9220 5355 9272 5364
rect 1676 5108 1728 5160
rect 2872 5176 2924 5228
rect 4068 5176 4120 5228
rect 4620 5176 4672 5228
rect 7380 5219 7432 5228
rect 3516 5108 3568 5160
rect 2780 5040 2832 5092
rect 4528 5108 4580 5160
rect 4896 5151 4948 5160
rect 4896 5117 4905 5151
rect 4905 5117 4939 5151
rect 4939 5117 4948 5151
rect 4896 5108 4948 5117
rect 7380 5185 7389 5219
rect 7389 5185 7423 5219
rect 7423 5185 7432 5219
rect 7380 5176 7432 5185
rect 9220 5321 9229 5355
rect 9229 5321 9263 5355
rect 9263 5321 9272 5355
rect 9220 5312 9272 5321
rect 9680 5312 9732 5364
rect 10508 5312 10560 5364
rect 12440 5312 12492 5364
rect 12532 5312 12584 5364
rect 13820 5312 13872 5364
rect 14096 5312 14148 5364
rect 14556 5312 14608 5364
rect 9496 5176 9548 5228
rect 10140 5176 10192 5228
rect 12164 5244 12216 5296
rect 12256 5244 12308 5296
rect 7932 5108 7984 5160
rect 8576 5108 8628 5160
rect 4804 5040 4856 5092
rect 5172 5083 5224 5092
rect 5172 5049 5206 5083
rect 5206 5049 5224 5083
rect 5172 5040 5224 5049
rect 5816 5040 5868 5092
rect 6460 5040 6512 5092
rect 7012 5040 7064 5092
rect 7196 5040 7248 5092
rect 7380 5040 7432 5092
rect 8300 5040 8352 5092
rect 1400 5015 1452 5024
rect 1400 4981 1409 5015
rect 1409 4981 1443 5015
rect 1443 4981 1452 5015
rect 1400 4972 1452 4981
rect 3240 4972 3292 5024
rect 3700 5015 3752 5024
rect 3700 4981 3709 5015
rect 3709 4981 3743 5015
rect 3743 4981 3752 5015
rect 3700 4972 3752 4981
rect 5540 4972 5592 5024
rect 5632 4972 5684 5024
rect 9036 5040 9088 5092
rect 8760 4972 8812 5024
rect 10416 5108 10468 5160
rect 11520 5108 11572 5160
rect 12624 5176 12676 5228
rect 14004 5244 14056 5296
rect 13360 5176 13412 5228
rect 13912 5176 13964 5228
rect 14096 5176 14148 5228
rect 12256 5108 12308 5160
rect 13084 5108 13136 5160
rect 13820 5108 13872 5160
rect 9680 5015 9732 5024
rect 9680 4981 9689 5015
rect 9689 4981 9723 5015
rect 9723 4981 9732 5015
rect 9680 4972 9732 4981
rect 10968 5040 11020 5092
rect 11520 4972 11572 5024
rect 11704 4972 11756 5024
rect 13912 5040 13964 5092
rect 13636 5015 13688 5024
rect 13636 4981 13645 5015
rect 13645 4981 13679 5015
rect 13679 4981 13688 5015
rect 13636 4972 13688 4981
rect 13820 4972 13872 5024
rect 14188 4972 14240 5024
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 2964 4768 3016 4820
rect 3608 4768 3660 4820
rect 3700 4768 3752 4820
rect 4988 4768 5040 4820
rect 5356 4768 5408 4820
rect 5632 4768 5684 4820
rect 1676 4743 1728 4752
rect 1676 4709 1710 4743
rect 1710 4709 1728 4743
rect 1676 4700 1728 4709
rect 4436 4743 4488 4752
rect 4436 4709 4445 4743
rect 4445 4709 4479 4743
rect 4479 4709 4488 4743
rect 4436 4700 4488 4709
rect 4804 4700 4856 4752
rect 8392 4768 8444 4820
rect 6736 4743 6788 4752
rect 6736 4709 6770 4743
rect 6770 4709 6788 4743
rect 6736 4700 6788 4709
rect 3332 4607 3384 4616
rect 3332 4573 3341 4607
rect 3341 4573 3375 4607
rect 3375 4573 3384 4607
rect 5356 4632 5408 4684
rect 5632 4675 5684 4684
rect 5632 4641 5641 4675
rect 5641 4641 5675 4675
rect 5675 4641 5684 4675
rect 5632 4632 5684 4641
rect 5816 4632 5868 4684
rect 3332 4564 3384 4573
rect 2872 4539 2924 4548
rect 2872 4505 2881 4539
rect 2881 4505 2915 4539
rect 2915 4505 2924 4539
rect 2872 4496 2924 4505
rect 3792 4564 3844 4616
rect 6276 4632 6328 4684
rect 7012 4632 7064 4684
rect 7840 4632 7892 4684
rect 8300 4632 8352 4684
rect 8576 4768 8628 4820
rect 9128 4768 9180 4820
rect 9036 4700 9088 4752
rect 5356 4496 5408 4548
rect 3792 4428 3844 4480
rect 7564 4564 7616 4616
rect 8760 4564 8812 4616
rect 5724 4428 5776 4480
rect 5816 4428 5868 4480
rect 7840 4471 7892 4480
rect 7840 4437 7849 4471
rect 7849 4437 7883 4471
rect 7883 4437 7892 4471
rect 7840 4428 7892 4437
rect 8024 4496 8076 4548
rect 8668 4496 8720 4548
rect 9220 4632 9272 4684
rect 10232 4768 10284 4820
rect 9956 4700 10008 4752
rect 10600 4700 10652 4752
rect 11244 4743 11296 4752
rect 11244 4709 11253 4743
rect 11253 4709 11287 4743
rect 11287 4709 11296 4743
rect 11980 4768 12032 4820
rect 12256 4768 12308 4820
rect 12624 4768 12676 4820
rect 12900 4768 12952 4820
rect 11244 4700 11296 4709
rect 12348 4700 12400 4752
rect 11704 4675 11756 4684
rect 11704 4641 11713 4675
rect 11713 4641 11747 4675
rect 11747 4641 11756 4675
rect 11704 4632 11756 4641
rect 13452 4700 13504 4752
rect 14096 4632 14148 4684
rect 14464 4675 14516 4684
rect 14464 4641 14473 4675
rect 14473 4641 14507 4675
rect 14507 4641 14516 4675
rect 14464 4632 14516 4641
rect 9496 4564 9548 4616
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 11152 4564 11204 4616
rect 10876 4539 10928 4548
rect 10876 4505 10885 4539
rect 10885 4505 10919 4539
rect 10919 4505 10928 4539
rect 10876 4496 10928 4505
rect 10968 4496 11020 4548
rect 12072 4564 12124 4616
rect 12440 4564 12492 4616
rect 11888 4496 11940 4548
rect 12624 4607 12676 4616
rect 12624 4573 12633 4607
rect 12633 4573 12667 4607
rect 12667 4573 12676 4607
rect 12624 4564 12676 4573
rect 12900 4564 12952 4616
rect 12256 4428 12308 4480
rect 14924 4428 14976 4480
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 2780 4224 2832 4276
rect 1032 4088 1084 4140
rect 1584 4088 1636 4140
rect 2504 4088 2556 4140
rect 5172 4224 5224 4276
rect 5540 4267 5592 4276
rect 5540 4233 5549 4267
rect 5549 4233 5583 4267
rect 5583 4233 5592 4267
rect 5540 4224 5592 4233
rect 5632 4224 5684 4276
rect 7840 4224 7892 4276
rect 9128 4224 9180 4276
rect 4160 4156 4212 4208
rect 4344 4156 4396 4208
rect 1400 4020 1452 4072
rect 1952 4020 2004 4072
rect 2596 4063 2648 4072
rect 2596 4029 2605 4063
rect 2605 4029 2639 4063
rect 2639 4029 2648 4063
rect 2596 4020 2648 4029
rect 4896 4063 4948 4072
rect 1952 3927 2004 3936
rect 1952 3893 1961 3927
rect 1961 3893 1995 3927
rect 1995 3893 2004 3927
rect 1952 3884 2004 3893
rect 2044 3927 2096 3936
rect 2044 3893 2053 3927
rect 2053 3893 2087 3927
rect 2087 3893 2096 3927
rect 2320 3952 2372 4004
rect 2780 3952 2832 4004
rect 4896 4029 4905 4063
rect 4905 4029 4939 4063
rect 4939 4029 4948 4063
rect 4896 4020 4948 4029
rect 5540 4088 5592 4140
rect 8208 4156 8260 4208
rect 10048 4156 10100 4208
rect 11060 4224 11112 4276
rect 11888 4224 11940 4276
rect 11980 4224 12032 4276
rect 15292 4224 15344 4276
rect 6920 4088 6972 4140
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 9036 4088 9088 4140
rect 10324 4088 10376 4140
rect 10416 4088 10468 4140
rect 10876 4156 10928 4208
rect 11520 4156 11572 4208
rect 12256 4156 12308 4208
rect 12808 4156 12860 4208
rect 13728 4156 13780 4208
rect 10968 4131 11020 4140
rect 8484 4063 8536 4072
rect 8484 4029 8493 4063
rect 8493 4029 8527 4063
rect 8527 4029 8536 4063
rect 8484 4020 8536 4029
rect 10508 4020 10560 4072
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 11060 4088 11112 4140
rect 11336 4020 11388 4072
rect 12164 4088 12216 4140
rect 12624 4088 12676 4140
rect 12900 4088 12952 4140
rect 13544 4088 13596 4140
rect 12532 4020 12584 4072
rect 2044 3884 2096 3893
rect 3424 3884 3476 3936
rect 4160 3952 4212 4004
rect 5356 3952 5408 4004
rect 5908 3995 5960 4004
rect 5908 3961 5917 3995
rect 5917 3961 5951 3995
rect 5951 3961 5960 3995
rect 5908 3952 5960 3961
rect 6552 3952 6604 4004
rect 6828 3952 6880 4004
rect 7472 3952 7524 4004
rect 7012 3884 7064 3936
rect 8116 3952 8168 4004
rect 8852 3952 8904 4004
rect 7748 3884 7800 3936
rect 8300 3884 8352 3936
rect 10416 3927 10468 3936
rect 10416 3893 10425 3927
rect 10425 3893 10459 3927
rect 10459 3893 10468 3927
rect 10416 3884 10468 3893
rect 11060 3952 11112 4004
rect 11520 3952 11572 4004
rect 11888 3952 11940 4004
rect 12072 3884 12124 3936
rect 13636 3952 13688 4004
rect 12808 3927 12860 3936
rect 12808 3893 12817 3927
rect 12817 3893 12851 3927
rect 12851 3893 12860 3927
rect 12808 3884 12860 3893
rect 12992 3884 13044 3936
rect 13268 3884 13320 3936
rect 15476 3952 15528 4004
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 572 3680 624 3732
rect 1492 3680 1544 3732
rect 1860 3723 1912 3732
rect 1860 3689 1869 3723
rect 1869 3689 1903 3723
rect 1903 3689 1912 3723
rect 1860 3680 1912 3689
rect 3148 3680 3200 3732
rect 3424 3680 3476 3732
rect 4160 3680 4212 3732
rect 5080 3680 5132 3732
rect 5724 3680 5776 3732
rect 204 3612 256 3664
rect 3700 3612 3752 3664
rect 3884 3612 3936 3664
rect 940 3544 992 3596
rect 3240 3587 3292 3596
rect 3240 3553 3249 3587
rect 3249 3553 3283 3587
rect 3283 3553 3292 3587
rect 3240 3544 3292 3553
rect 3424 3544 3476 3596
rect 3608 3544 3660 3596
rect 5908 3612 5960 3664
rect 6092 3612 6144 3664
rect 7196 3680 7248 3732
rect 8024 3680 8076 3732
rect 9036 3680 9088 3732
rect 9312 3680 9364 3732
rect 10416 3680 10468 3732
rect 5356 3587 5408 3596
rect 5356 3553 5365 3587
rect 5365 3553 5399 3587
rect 5399 3553 5408 3587
rect 5356 3544 5408 3553
rect 6184 3544 6236 3596
rect 7472 3612 7524 3664
rect 8116 3612 8168 3664
rect 10232 3612 10284 3664
rect 10324 3612 10376 3664
rect 11060 3612 11112 3664
rect 11612 3612 11664 3664
rect 7840 3587 7892 3596
rect 2412 3476 2464 3528
rect 3516 3519 3568 3528
rect 3516 3485 3525 3519
rect 3525 3485 3559 3519
rect 3559 3485 3568 3519
rect 3516 3476 3568 3485
rect 4528 3476 4580 3528
rect 5172 3476 5224 3528
rect 1400 3451 1452 3460
rect 1400 3417 1409 3451
rect 1409 3417 1443 3451
rect 1443 3417 1452 3451
rect 1400 3408 1452 3417
rect 1952 3408 2004 3460
rect 4436 3408 4488 3460
rect 4988 3451 5040 3460
rect 4988 3417 4997 3451
rect 4997 3417 5031 3451
rect 5031 3417 5040 3451
rect 5724 3476 5776 3528
rect 7840 3553 7849 3587
rect 7849 3553 7883 3587
rect 7883 3553 7892 3587
rect 7840 3544 7892 3553
rect 6552 3476 6604 3528
rect 6920 3476 6972 3528
rect 7380 3476 7432 3528
rect 8116 3476 8168 3528
rect 9496 3544 9548 3596
rect 4988 3408 5040 3417
rect 6736 3408 6788 3460
rect 8576 3408 8628 3460
rect 8760 3408 8812 3460
rect 9036 3408 9088 3460
rect 4068 3383 4120 3392
rect 4068 3349 4077 3383
rect 4077 3349 4111 3383
rect 4111 3349 4120 3383
rect 4068 3340 4120 3349
rect 4620 3340 4672 3392
rect 6092 3340 6144 3392
rect 6276 3340 6328 3392
rect 9680 3476 9732 3528
rect 9956 3544 10008 3596
rect 10324 3519 10376 3528
rect 10324 3485 10333 3519
rect 10333 3485 10367 3519
rect 10367 3485 10376 3519
rect 10324 3476 10376 3485
rect 10600 3544 10652 3596
rect 10968 3544 11020 3596
rect 11980 3544 12032 3596
rect 10692 3476 10744 3528
rect 10784 3476 10836 3528
rect 11612 3476 11664 3528
rect 12808 3680 12860 3732
rect 13084 3680 13136 3732
rect 13636 3680 13688 3732
rect 12348 3612 12400 3664
rect 12532 3655 12584 3664
rect 12532 3621 12541 3655
rect 12541 3621 12575 3655
rect 12575 3621 12584 3655
rect 12532 3612 12584 3621
rect 12900 3612 12952 3664
rect 14280 3544 14332 3596
rect 12440 3476 12492 3528
rect 12624 3519 12676 3528
rect 12624 3485 12633 3519
rect 12633 3485 12667 3519
rect 12667 3485 12676 3519
rect 12624 3476 12676 3485
rect 12992 3476 13044 3528
rect 13544 3476 13596 3528
rect 10416 3340 10468 3392
rect 11612 3340 11664 3392
rect 11888 3383 11940 3392
rect 11888 3349 11897 3383
rect 11897 3349 11931 3383
rect 11931 3349 11940 3383
rect 11888 3340 11940 3349
rect 12072 3383 12124 3392
rect 12072 3349 12081 3383
rect 12081 3349 12115 3383
rect 12115 3349 12124 3383
rect 12072 3340 12124 3349
rect 13820 3408 13872 3460
rect 14280 3408 14332 3460
rect 13728 3340 13780 3392
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 2412 3136 2464 3188
rect 2596 3000 2648 3052
rect 756 2932 808 2984
rect 5080 3136 5132 3188
rect 6552 3136 6604 3188
rect 6828 3179 6880 3188
rect 6828 3145 6837 3179
rect 6837 3145 6871 3179
rect 6871 3145 6880 3179
rect 6828 3136 6880 3145
rect 8024 3136 8076 3188
rect 9220 3179 9272 3188
rect 9220 3145 9229 3179
rect 9229 3145 9263 3179
rect 9263 3145 9272 3179
rect 9220 3136 9272 3145
rect 5816 3068 5868 3120
rect 4252 3000 4304 3052
rect 5448 3000 5500 3052
rect 5540 3000 5592 3052
rect 7380 3068 7432 3120
rect 6368 3000 6420 3052
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 7564 3000 7616 3052
rect 7932 3068 7984 3120
rect 10048 3136 10100 3188
rect 10324 3136 10376 3188
rect 10784 3136 10836 3188
rect 11152 3136 11204 3188
rect 11336 3136 11388 3188
rect 9588 3068 9640 3120
rect 12716 3136 12768 3188
rect 9404 3000 9456 3052
rect 9772 3043 9824 3052
rect 4528 2932 4580 2984
rect 4620 2932 4672 2984
rect 5724 2932 5776 2984
rect 5908 2975 5960 2984
rect 5908 2941 5917 2975
rect 5917 2941 5951 2975
rect 5951 2941 5960 2975
rect 5908 2932 5960 2941
rect 7012 2932 7064 2984
rect 8668 2932 8720 2984
rect 8944 2932 8996 2984
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 4436 2864 4488 2916
rect 10508 3000 10560 3052
rect 10048 2975 10100 2984
rect 10048 2941 10057 2975
rect 10057 2941 10091 2975
rect 10091 2941 10100 2975
rect 10692 3000 10744 3052
rect 11060 3000 11112 3052
rect 10048 2932 10100 2941
rect 11428 2932 11480 2984
rect 11612 2975 11664 2984
rect 11612 2941 11621 2975
rect 11621 2941 11655 2975
rect 11655 2941 11664 2975
rect 11612 2932 11664 2941
rect 12072 3000 12124 3052
rect 16304 3068 16356 3120
rect 12440 3000 12492 3052
rect 12532 3000 12584 3052
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 13084 3000 13136 3052
rect 13912 3000 13964 3052
rect 14372 3043 14424 3052
rect 2320 2796 2372 2848
rect 4804 2796 4856 2848
rect 5356 2796 5408 2848
rect 6920 2796 6972 2848
rect 7012 2796 7064 2848
rect 9936 2864 9988 2916
rect 10968 2864 11020 2916
rect 11152 2864 11204 2916
rect 11796 2864 11848 2916
rect 10508 2796 10560 2848
rect 10600 2796 10652 2848
rect 11428 2796 11480 2848
rect 12624 2932 12676 2984
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 14556 3000 14608 3052
rect 12164 2864 12216 2916
rect 13820 2864 13872 2916
rect 14556 2864 14608 2916
rect 15200 2864 15252 2916
rect 12440 2839 12492 2848
rect 12440 2805 12449 2839
rect 12449 2805 12483 2839
rect 12483 2805 12492 2839
rect 12440 2796 12492 2805
rect 14004 2796 14056 2848
rect 14096 2796 14148 2848
rect 15108 2796 15160 2848
rect 16764 2796 16816 2848
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 2596 2592 2648 2644
rect 3148 2592 3200 2644
rect 3332 2592 3384 2644
rect 4160 2592 4212 2644
rect 1768 2524 1820 2576
rect 4896 2592 4948 2644
rect 5816 2592 5868 2644
rect 8576 2635 8628 2644
rect 2412 2456 2464 2508
rect 4620 2499 4672 2508
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 4344 2388 4396 2440
rect 4620 2465 4629 2499
rect 4629 2465 4663 2499
rect 4663 2465 4672 2499
rect 4620 2456 4672 2465
rect 5632 2456 5684 2508
rect 5172 2388 5224 2440
rect 8576 2601 8585 2635
rect 8585 2601 8619 2635
rect 8619 2601 8628 2635
rect 8576 2592 8628 2601
rect 8944 2592 8996 2644
rect 9036 2592 9088 2644
rect 9956 2524 10008 2576
rect 7012 2456 7064 2508
rect 1400 2252 1452 2304
rect 3976 2320 4028 2372
rect 2504 2252 2556 2304
rect 4160 2252 4212 2304
rect 4436 2320 4488 2372
rect 4528 2252 4580 2304
rect 6460 2388 6512 2440
rect 8208 2456 8260 2508
rect 11152 2592 11204 2644
rect 12440 2592 12492 2644
rect 12624 2635 12676 2644
rect 12624 2601 12633 2635
rect 12633 2601 12667 2635
rect 12667 2601 12676 2635
rect 12624 2592 12676 2601
rect 13084 2592 13136 2644
rect 13268 2592 13320 2644
rect 13820 2592 13872 2644
rect 14832 2592 14884 2644
rect 11060 2524 11112 2576
rect 13636 2524 13688 2576
rect 15108 2567 15160 2576
rect 5448 2320 5500 2372
rect 9128 2388 9180 2440
rect 9404 2320 9456 2372
rect 11428 2456 11480 2508
rect 11980 2499 12032 2508
rect 11980 2465 11989 2499
rect 11989 2465 12023 2499
rect 12023 2465 12032 2499
rect 11980 2456 12032 2465
rect 12072 2456 12124 2508
rect 14004 2456 14056 2508
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 10692 2388 10744 2440
rect 11612 2388 11664 2440
rect 12900 2388 12952 2440
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 15108 2533 15117 2567
rect 15117 2533 15151 2567
rect 15151 2533 15160 2567
rect 15108 2524 15160 2533
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 14832 2499 14884 2508
rect 14832 2465 14841 2499
rect 14841 2465 14875 2499
rect 14875 2465 14884 2499
rect 14832 2456 14884 2465
rect 13268 2388 13320 2397
rect 14464 2431 14516 2440
rect 14464 2397 14473 2431
rect 14473 2397 14507 2431
rect 14507 2397 14516 2431
rect 14464 2388 14516 2397
rect 14740 2320 14792 2372
rect 6276 2252 6328 2304
rect 9956 2252 10008 2304
rect 11060 2252 11112 2304
rect 11704 2252 11756 2304
rect 15476 2252 15528 2304
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 848 2048 900 2100
rect 11612 2048 11664 2100
rect 12164 2048 12216 2100
rect 13912 2048 13964 2100
rect 3332 1980 3384 2032
rect 9680 1980 9732 2032
rect 14464 1980 14516 2032
rect 3792 1912 3844 1964
rect 11980 1912 12032 1964
rect 12348 1912 12400 1964
rect 15384 1912 15436 1964
rect 15936 1912 15988 1964
rect 1216 1844 1268 1896
rect 6000 1844 6052 1896
rect 7380 1844 7432 1896
rect 8484 1844 8536 1896
rect 8760 1844 8812 1896
rect 10140 1844 10192 1896
rect 14188 1844 14240 1896
rect 4436 1776 4488 1828
rect 11244 1776 11296 1828
rect 2412 1708 2464 1760
rect 10324 1708 10376 1760
rect 10416 1708 10468 1760
rect 14924 1708 14976 1760
rect 2044 1640 2096 1692
rect 6276 1640 6328 1692
rect 7932 1640 7984 1692
rect 9588 1640 9640 1692
rect 3976 1572 4028 1624
rect 11888 1572 11940 1624
rect 2872 1504 2924 1556
rect 5356 1436 5408 1488
rect 14832 1436 14884 1488
rect 8668 1368 8720 1420
rect 12624 1368 12676 1420
rect 7840 1300 7892 1352
rect 9312 1300 9364 1352
rect 7104 1232 7156 1284
rect 10968 1232 11020 1284
rect 8852 1164 8904 1216
rect 10232 1164 10284 1216
<< metal2 >>
rect 202 19520 258 20000
rect 570 19520 626 20000
rect 938 19520 994 20000
rect 1398 19520 1454 20000
rect 1766 19520 1822 20000
rect 2226 19520 2282 20000
rect 2594 19520 2650 20000
rect 2870 19544 2926 19553
rect 216 16454 244 19520
rect 584 18426 612 19520
rect 572 18420 624 18426
rect 572 18362 624 18368
rect 204 16448 256 16454
rect 204 16390 256 16396
rect 952 16017 980 19520
rect 1308 17604 1360 17610
rect 1308 17546 1360 17552
rect 938 16008 994 16017
rect 938 15943 994 15952
rect 1216 15564 1268 15570
rect 1216 15506 1268 15512
rect 1228 9897 1256 15506
rect 1320 10810 1348 17546
rect 1412 17542 1440 19520
rect 1780 18154 1808 19520
rect 1768 18148 1820 18154
rect 1768 18090 1820 18096
rect 2240 17746 2268 19520
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 1400 17536 1452 17542
rect 1400 17478 1452 17484
rect 2136 17060 2188 17066
rect 2136 17002 2188 17008
rect 2148 16697 2176 17002
rect 2134 16688 2190 16697
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1860 16652 1912 16658
rect 2134 16623 2190 16632
rect 2504 16652 2556 16658
rect 1860 16594 1912 16600
rect 2504 16594 2556 16600
rect 1596 14618 1624 16594
rect 1872 15745 1900 16594
rect 2320 15972 2372 15978
rect 2320 15914 2372 15920
rect 1858 15736 1914 15745
rect 1858 15671 1914 15680
rect 1676 14884 1728 14890
rect 1676 14826 1728 14832
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1504 12617 1532 13262
rect 1490 12608 1546 12617
rect 1490 12543 1546 12552
rect 1308 10804 1360 10810
rect 1308 10746 1360 10752
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1214 9888 1270 9897
rect 1214 9823 1270 9832
rect 1308 8968 1360 8974
rect 1308 8910 1360 8916
rect 1216 8832 1268 8838
rect 1216 8774 1268 8780
rect 938 7984 994 7993
rect 938 7919 994 7928
rect 754 7168 810 7177
rect 754 7103 810 7112
rect 572 3732 624 3738
rect 572 3674 624 3680
rect 204 3664 256 3670
rect 204 3606 256 3612
rect 216 480 244 3606
rect 584 480 612 3674
rect 768 2990 796 7103
rect 846 5264 902 5273
rect 846 5199 902 5208
rect 756 2984 808 2990
rect 756 2926 808 2932
rect 860 2106 888 5199
rect 952 3602 980 7919
rect 1124 7336 1176 7342
rect 1124 7278 1176 7284
rect 1032 4140 1084 4146
rect 1032 4082 1084 4088
rect 940 3596 992 3602
rect 940 3538 992 3544
rect 848 2100 900 2106
rect 848 2042 900 2048
rect 1044 480 1072 4082
rect 1136 513 1164 7278
rect 1228 1902 1256 8774
rect 1320 6866 1348 8910
rect 1412 7993 1440 10542
rect 1504 8650 1532 12543
rect 1596 12442 1624 13806
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1688 11914 1716 14826
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1596 11886 1716 11914
rect 1596 8974 1624 11886
rect 1780 11257 1808 14758
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1872 12986 1900 13126
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1858 11928 1914 11937
rect 1858 11863 1914 11872
rect 1872 11286 1900 11863
rect 1860 11280 1912 11286
rect 1766 11248 1822 11257
rect 1860 11222 1912 11228
rect 1766 11183 1822 11192
rect 1766 11112 1822 11121
rect 1766 11047 1822 11056
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1504 8622 1716 8650
rect 1398 7984 1454 7993
rect 1398 7919 1454 7928
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1308 6860 1360 6866
rect 1308 6802 1360 6808
rect 1320 5846 1348 6802
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1308 5840 1360 5846
rect 1412 5817 1440 5850
rect 1308 5782 1360 5788
rect 1398 5808 1454 5817
rect 1320 2553 1348 5782
rect 1398 5743 1454 5752
rect 1398 5128 1454 5137
rect 1398 5063 1454 5072
rect 1412 5030 1440 5063
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 1412 3466 1440 4014
rect 1504 3738 1532 7686
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 4146 1624 6598
rect 1688 5166 1716 8622
rect 1780 6254 1808 11047
rect 1860 10532 1912 10538
rect 1860 10474 1912 10480
rect 1872 9722 1900 10474
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1964 8650 1992 12582
rect 2056 12322 2084 14350
rect 2148 12481 2176 14350
rect 2332 13734 2360 15914
rect 2516 15314 2544 16594
rect 2608 15473 2636 19520
rect 2962 19520 3018 20000
rect 3422 19520 3478 20000
rect 3790 19520 3846 20000
rect 4250 19520 4306 20000
rect 4618 19520 4674 20000
rect 4986 19520 5042 20000
rect 5446 19520 5502 20000
rect 5814 19520 5870 20000
rect 6274 19520 6330 20000
rect 6642 19520 6698 20000
rect 7010 19520 7066 20000
rect 7470 19520 7526 20000
rect 7838 19520 7894 20000
rect 8298 19520 8354 20000
rect 8666 19520 8722 20000
rect 9034 19520 9090 20000
rect 9494 19520 9550 20000
rect 9862 19520 9918 20000
rect 10322 19520 10378 20000
rect 10690 19520 10746 20000
rect 11058 19520 11114 20000
rect 11518 19520 11574 20000
rect 11886 19520 11942 20000
rect 12346 19520 12402 20000
rect 12714 19520 12770 20000
rect 13082 19520 13138 20000
rect 13542 19520 13598 20000
rect 13910 19520 13966 20000
rect 14370 19520 14426 20000
rect 14738 19520 14794 20000
rect 15106 19520 15162 20000
rect 15566 19520 15622 20000
rect 15934 19520 15990 20000
rect 16394 19520 16450 20000
rect 16762 19520 16818 20000
rect 2870 19479 2926 19488
rect 2778 17640 2834 17649
rect 2778 17575 2834 17584
rect 2792 16114 2820 17575
rect 2884 16250 2912 19479
rect 2976 17649 3004 19520
rect 3436 17814 3464 19520
rect 3424 17808 3476 17814
rect 3424 17750 3476 17756
rect 2962 17640 3018 17649
rect 2962 17575 3018 17584
rect 3421 17436 3717 17456
rect 3477 17434 3501 17436
rect 3557 17434 3581 17436
rect 3637 17434 3661 17436
rect 3499 17382 3501 17434
rect 3563 17382 3575 17434
rect 3637 17382 3639 17434
rect 3477 17380 3501 17382
rect 3557 17380 3581 17382
rect 3637 17380 3661 17382
rect 3421 17360 3717 17380
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 3056 17060 3108 17066
rect 3056 17002 3108 17008
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2686 15736 2742 15745
rect 2686 15671 2742 15680
rect 2594 15464 2650 15473
rect 2594 15399 2650 15408
rect 2516 15286 2636 15314
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2516 14074 2544 15098
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 2608 14006 2636 15286
rect 2700 14890 2728 15671
rect 2792 15065 2820 15846
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2872 15428 2924 15434
rect 2872 15370 2924 15376
rect 2778 15056 2834 15065
rect 2884 15026 2912 15370
rect 2778 14991 2834 15000
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2596 14000 2648 14006
rect 2596 13942 2648 13948
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2240 12986 2268 13398
rect 2700 13394 2728 14554
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2410 13288 2466 13297
rect 2410 13223 2412 13232
rect 2464 13223 2466 13232
rect 2412 13194 2464 13200
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2134 12472 2190 12481
rect 2134 12407 2190 12416
rect 2056 12294 2268 12322
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1872 8622 1992 8650
rect 1872 7562 1900 8622
rect 1950 8528 2006 8537
rect 1950 8463 2006 8472
rect 1964 8430 1992 8463
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1872 7534 1992 7562
rect 1858 7304 1914 7313
rect 1858 7239 1914 7248
rect 1872 6458 1900 7239
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1768 6248 1820 6254
rect 1820 6208 1900 6236
rect 1768 6190 1820 6196
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1674 4856 1730 4865
rect 1674 4791 1730 4800
rect 1688 4758 1716 4791
rect 1676 4752 1728 4758
rect 1676 4694 1728 4700
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1674 4040 1730 4049
rect 1674 3975 1730 3984
rect 1492 3732 1544 3738
rect 1492 3674 1544 3680
rect 1400 3460 1452 3466
rect 1400 3402 1452 3408
rect 1688 3369 1716 3975
rect 1674 3360 1730 3369
rect 1674 3295 1730 3304
rect 1780 2582 1808 5646
rect 1872 4185 1900 6208
rect 1858 4176 1914 4185
rect 1858 4111 1914 4120
rect 1964 4078 1992 7534
rect 2056 5846 2084 11494
rect 2148 10810 2176 12174
rect 2240 10810 2268 12294
rect 2318 11656 2374 11665
rect 2318 11591 2320 11600
rect 2372 11591 2374 11600
rect 2320 11562 2372 11568
rect 2516 11121 2544 13330
rect 2792 13258 2820 14826
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2884 13977 2912 14758
rect 2870 13968 2926 13977
rect 2870 13903 2926 13912
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2700 11801 2728 12242
rect 2686 11792 2742 11801
rect 2686 11727 2742 11736
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2688 11552 2740 11558
rect 2688 11494 2740 11500
rect 2502 11112 2558 11121
rect 2502 11047 2558 11056
rect 2504 11008 2556 11014
rect 2502 10976 2504 10985
rect 2556 10976 2558 10985
rect 2502 10911 2558 10920
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2502 10704 2558 10713
rect 2502 10639 2504 10648
rect 2556 10639 2558 10648
rect 2504 10610 2556 10616
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2136 9512 2188 9518
rect 2240 9489 2268 10406
rect 2412 10192 2464 10198
rect 2516 10180 2544 10610
rect 2464 10152 2544 10180
rect 2412 10134 2464 10140
rect 2502 9888 2558 9897
rect 2502 9823 2558 9832
rect 2136 9454 2188 9460
rect 2226 9480 2282 9489
rect 2148 9042 2176 9454
rect 2226 9415 2282 9424
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2332 9178 2360 9318
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2134 7848 2190 7857
rect 2134 7783 2190 7792
rect 2044 5840 2096 5846
rect 2044 5782 2096 5788
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1952 3936 2004 3942
rect 1858 3904 1914 3913
rect 1952 3878 2004 3884
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 2148 3890 2176 7783
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2240 7002 2268 7142
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2226 6896 2282 6905
rect 2226 6831 2282 6840
rect 2240 5642 2268 6831
rect 2228 5636 2280 5642
rect 2228 5578 2280 5584
rect 2332 4010 2360 8230
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2424 6089 2452 6258
rect 2410 6080 2466 6089
rect 2410 6015 2466 6024
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 1858 3839 1914 3848
rect 1872 3738 1900 3839
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 1964 3466 1992 3878
rect 1952 3460 2004 3466
rect 1952 3402 2004 3408
rect 1768 2576 1820 2582
rect 1306 2544 1362 2553
rect 1768 2518 1820 2524
rect 1306 2479 1362 2488
rect 1400 2304 1452 2310
rect 1400 2246 1452 2252
rect 1216 1896 1268 1902
rect 1216 1838 1268 1844
rect 1122 504 1178 513
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1412 480 1440 2246
rect 1858 2000 1914 2009
rect 1858 1935 1914 1944
rect 1872 480 1900 1935
rect 2056 1698 2084 3878
rect 2148 3862 2360 3890
rect 2332 2854 2360 3862
rect 2424 3534 2452 5714
rect 2516 5273 2544 9823
rect 2700 9625 2728 11494
rect 2792 11286 2820 11698
rect 2780 11280 2832 11286
rect 2780 11222 2832 11228
rect 2792 10606 2820 11222
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2792 10130 2820 10542
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2884 10033 2912 13806
rect 2976 12594 3004 15438
rect 3068 14793 3096 17002
rect 3620 16658 3648 17138
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 3608 16652 3660 16658
rect 3608 16594 3660 16600
rect 3148 16516 3200 16522
rect 3148 16458 3200 16464
rect 3054 14784 3110 14793
rect 3054 14719 3110 14728
rect 3160 14600 3188 16458
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3252 15434 3280 15846
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 3252 14618 3280 15370
rect 3068 14572 3188 14600
rect 3240 14612 3292 14618
rect 3068 12850 3096 14572
rect 3240 14554 3292 14560
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3068 12753 3096 12786
rect 3054 12744 3110 12753
rect 3054 12679 3110 12688
rect 2976 12566 3096 12594
rect 2962 12472 3018 12481
rect 2962 12407 3018 12416
rect 2870 10024 2926 10033
rect 2870 9959 2926 9968
rect 2686 9616 2742 9625
rect 2686 9551 2742 9560
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 8498 2636 9318
rect 2700 8945 2728 9386
rect 2778 9072 2834 9081
rect 2778 9007 2834 9016
rect 2686 8936 2742 8945
rect 2686 8871 2742 8880
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2594 7576 2650 7585
rect 2594 7511 2650 7520
rect 2608 7410 2636 7511
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2596 6928 2648 6934
rect 2596 6870 2648 6876
rect 2608 6186 2636 6870
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2502 5264 2558 5273
rect 2502 5199 2558 5208
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2424 3194 2452 3470
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 2412 2508 2464 2514
rect 2412 2450 2464 2456
rect 2424 1766 2452 2450
rect 2516 2310 2544 4082
rect 2608 4078 2636 6122
rect 2700 4264 2728 7890
rect 2792 5846 2820 9007
rect 2884 8498 2912 9454
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2884 7750 2912 8434
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2884 7546 2912 7686
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2778 5672 2834 5681
rect 2778 5607 2834 5616
rect 2792 5098 2820 5607
rect 2884 5234 2912 7346
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2976 4826 3004 12407
rect 3068 8129 3096 12566
rect 3054 8120 3110 8129
rect 3054 8055 3110 8064
rect 3054 7440 3110 7449
rect 3054 7375 3056 7384
rect 3108 7375 3110 7384
rect 3056 7346 3108 7352
rect 3054 6488 3110 6497
rect 3054 6423 3110 6432
rect 3068 6390 3096 6423
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2870 4584 2926 4593
rect 2870 4519 2872 4528
rect 2924 4519 2926 4528
rect 2872 4490 2924 4496
rect 2870 4312 2926 4321
rect 2780 4276 2832 4282
rect 2700 4236 2780 4264
rect 2870 4247 2926 4256
rect 2780 4218 2832 4224
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2608 3058 2636 4014
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2608 2650 2636 2994
rect 2686 2952 2742 2961
rect 2686 2887 2742 2896
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2412 1760 2464 1766
rect 2412 1702 2464 1708
rect 2044 1692 2096 1698
rect 2044 1634 2096 1640
rect 2226 1320 2282 1329
rect 2226 1255 2282 1264
rect 2240 480 2268 1255
rect 2700 480 2728 2887
rect 2792 1465 2820 3946
rect 2884 1562 2912 4247
rect 3160 3738 3188 14418
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3252 13190 3280 14350
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3344 12889 3372 16594
rect 3421 16348 3717 16368
rect 3477 16346 3501 16348
rect 3557 16346 3581 16348
rect 3637 16346 3661 16348
rect 3499 16294 3501 16346
rect 3563 16294 3575 16346
rect 3637 16294 3639 16346
rect 3477 16292 3501 16294
rect 3557 16292 3581 16294
rect 3637 16292 3661 16294
rect 3421 16272 3717 16292
rect 3804 16096 3832 19520
rect 4066 18592 4122 18601
rect 4066 18527 4122 18536
rect 4080 18018 4108 18527
rect 4068 18012 4120 18018
rect 4068 17954 4120 17960
rect 4264 17218 4292 19520
rect 4264 17190 4568 17218
rect 4344 17060 4396 17066
rect 4344 17002 4396 17008
rect 3974 16688 4030 16697
rect 3974 16623 4030 16632
rect 3988 16182 4016 16623
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 3976 16176 4028 16182
rect 4080 16153 4108 16390
rect 3976 16118 4028 16124
rect 4066 16144 4122 16153
rect 3804 16068 3924 16096
rect 3790 15872 3846 15881
rect 3790 15807 3846 15816
rect 3421 15260 3717 15280
rect 3477 15258 3501 15260
rect 3557 15258 3581 15260
rect 3637 15258 3661 15260
rect 3499 15206 3501 15258
rect 3563 15206 3575 15258
rect 3637 15206 3639 15258
rect 3477 15204 3501 15206
rect 3557 15204 3581 15206
rect 3637 15204 3661 15206
rect 3421 15184 3717 15204
rect 3804 15026 3832 15807
rect 3896 15201 3924 16068
rect 3988 15450 4016 16118
rect 4066 16079 4122 16088
rect 4158 15600 4214 15609
rect 4158 15535 4160 15544
rect 4212 15535 4214 15544
rect 4160 15506 4212 15512
rect 3988 15422 4108 15450
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3882 15192 3938 15201
rect 3882 15127 3938 15136
rect 3884 15088 3936 15094
rect 3884 15030 3936 15036
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3792 14340 3844 14346
rect 3792 14282 3844 14288
rect 3421 14172 3717 14192
rect 3477 14170 3501 14172
rect 3557 14170 3581 14172
rect 3637 14170 3661 14172
rect 3499 14118 3501 14170
rect 3563 14118 3575 14170
rect 3637 14118 3639 14170
rect 3477 14116 3501 14118
rect 3557 14116 3581 14118
rect 3637 14116 3661 14118
rect 3421 14096 3717 14116
rect 3804 13938 3832 14282
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3792 13456 3844 13462
rect 3792 13398 3844 13404
rect 3421 13084 3717 13104
rect 3477 13082 3501 13084
rect 3557 13082 3581 13084
rect 3637 13082 3661 13084
rect 3499 13030 3501 13082
rect 3563 13030 3575 13082
rect 3637 13030 3639 13082
rect 3477 13028 3501 13030
rect 3557 13028 3581 13030
rect 3637 13028 3661 13030
rect 3421 13008 3717 13028
rect 3330 12880 3386 12889
rect 3330 12815 3386 12824
rect 3238 12744 3294 12753
rect 3804 12714 3832 13398
rect 3238 12679 3294 12688
rect 3424 12708 3476 12714
rect 3252 11898 3280 12679
rect 3424 12650 3476 12656
rect 3792 12708 3844 12714
rect 3792 12650 3844 12656
rect 3330 12336 3386 12345
rect 3330 12271 3386 12280
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3252 8362 3280 11018
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3238 7576 3294 7585
rect 3238 7511 3240 7520
rect 3292 7511 3294 7520
rect 3240 7482 3292 7488
rect 3344 5302 3372 12271
rect 3436 12209 3464 12650
rect 3422 12200 3478 12209
rect 3422 12135 3478 12144
rect 3421 11996 3717 12016
rect 3477 11994 3501 11996
rect 3557 11994 3581 11996
rect 3637 11994 3661 11996
rect 3499 11942 3501 11994
rect 3563 11942 3575 11994
rect 3637 11942 3639 11994
rect 3477 11940 3501 11942
rect 3557 11940 3581 11942
rect 3637 11940 3661 11942
rect 3421 11920 3717 11940
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3436 11082 3464 11562
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3421 10908 3717 10928
rect 3477 10906 3501 10908
rect 3557 10906 3581 10908
rect 3637 10906 3661 10908
rect 3499 10854 3501 10906
rect 3563 10854 3575 10906
rect 3637 10854 3639 10906
rect 3477 10852 3501 10854
rect 3557 10852 3581 10854
rect 3637 10852 3661 10854
rect 3421 10832 3717 10852
rect 3422 10024 3478 10033
rect 3422 9959 3424 9968
rect 3476 9959 3478 9968
rect 3424 9930 3476 9936
rect 3421 9820 3717 9840
rect 3477 9818 3501 9820
rect 3557 9818 3581 9820
rect 3637 9818 3661 9820
rect 3499 9766 3501 9818
rect 3563 9766 3575 9818
rect 3637 9766 3639 9818
rect 3477 9764 3501 9766
rect 3557 9764 3581 9766
rect 3637 9764 3661 9766
rect 3421 9744 3717 9764
rect 3514 9208 3570 9217
rect 3514 9143 3570 9152
rect 3528 8906 3556 9143
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3421 8732 3717 8752
rect 3477 8730 3501 8732
rect 3557 8730 3581 8732
rect 3637 8730 3661 8732
rect 3499 8678 3501 8730
rect 3563 8678 3575 8730
rect 3637 8678 3639 8730
rect 3477 8676 3501 8678
rect 3557 8676 3581 8678
rect 3637 8676 3661 8678
rect 3421 8656 3717 8676
rect 3421 7644 3717 7664
rect 3477 7642 3501 7644
rect 3557 7642 3581 7644
rect 3637 7642 3661 7644
rect 3499 7590 3501 7642
rect 3563 7590 3575 7642
rect 3637 7590 3639 7642
rect 3477 7588 3501 7590
rect 3557 7588 3581 7590
rect 3637 7588 3661 7590
rect 3421 7568 3717 7588
rect 3804 7342 3832 11018
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 3804 6458 3832 6802
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3790 6352 3846 6361
rect 3790 6287 3846 6296
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 3332 5296 3384 5302
rect 3332 5238 3384 5244
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 3516 5160 3568 5166
rect 3514 5128 3516 5137
rect 3568 5128 3570 5137
rect 3514 5063 3570 5072
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3252 3777 3280 4966
rect 3620 4826 3648 5238
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3712 4826 3740 4966
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3804 4622 3832 6287
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3238 3768 3294 3777
rect 3148 3732 3200 3738
rect 3238 3703 3294 3712
rect 3148 3674 3200 3680
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3252 3505 3280 3538
rect 3238 3496 3294 3505
rect 3238 3431 3294 3440
rect 3054 2816 3110 2825
rect 3054 2751 3110 2760
rect 2872 1556 2924 1562
rect 2872 1498 2924 1504
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 3068 480 3096 2751
rect 3146 2680 3202 2689
rect 3344 2650 3372 4558
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3514 4176 3570 4185
rect 3698 4176 3754 4185
rect 3570 4134 3648 4162
rect 3514 4111 3570 4120
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3436 3738 3464 3878
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3514 3632 3570 3641
rect 3424 3596 3476 3602
rect 3620 3602 3648 4134
rect 3698 4111 3754 4120
rect 3712 3670 3740 4111
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3514 3567 3570 3576
rect 3608 3596 3660 3602
rect 3424 3538 3476 3544
rect 3436 3505 3464 3538
rect 3528 3534 3556 3567
rect 3608 3538 3660 3544
rect 3516 3528 3568 3534
rect 3422 3496 3478 3505
rect 3516 3470 3568 3476
rect 3422 3431 3478 3440
rect 3421 3292 3717 3312
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3514 3088 3570 3097
rect 3514 3023 3570 3032
rect 3528 2836 3556 3023
rect 3436 2825 3556 2836
rect 3422 2816 3556 2825
rect 3478 2808 3556 2816
rect 3422 2751 3478 2760
rect 3146 2615 3148 2624
rect 3200 2615 3202 2624
rect 3332 2644 3384 2650
rect 3148 2586 3200 2592
rect 3332 2586 3384 2592
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 3344 2038 3372 2382
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3421 2128 3717 2148
rect 3332 2032 3384 2038
rect 3332 1974 3384 1980
rect 3804 1970 3832 4422
rect 3896 3670 3924 15030
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3882 3224 3938 3233
rect 3882 3159 3938 3168
rect 3792 1964 3844 1970
rect 3792 1906 3844 1912
rect 3514 1728 3570 1737
rect 3514 1663 3570 1672
rect 3528 480 3556 1663
rect 3896 480 3924 3159
rect 3988 2825 4016 15302
rect 4080 14958 4108 15422
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4080 13841 4108 14010
rect 4172 13938 4200 15302
rect 4264 14618 4292 16390
rect 4356 15162 4384 17002
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4344 14816 4396 14822
rect 4448 14793 4476 16594
rect 4540 16289 4568 17190
rect 4632 16794 4660 19520
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4724 16454 4752 16934
rect 4802 16552 4858 16561
rect 4802 16487 4858 16496
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4526 16280 4582 16289
rect 4526 16215 4582 16224
rect 4816 16114 4844 16487
rect 5000 16454 5028 19520
rect 5460 17610 5488 19520
rect 5828 17785 5856 19520
rect 5814 17776 5870 17785
rect 5814 17711 5870 17720
rect 5448 17604 5500 17610
rect 5448 17546 5500 17552
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 5276 16182 5304 16730
rect 5172 16176 5224 16182
rect 5172 16118 5224 16124
rect 5264 16176 5316 16182
rect 5264 16118 5316 16124
rect 4620 16108 4672 16114
rect 4804 16108 4856 16114
rect 4672 16068 4752 16096
rect 4620 16050 4672 16056
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4344 14758 4396 14764
rect 4434 14784 4490 14793
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4252 13864 4304 13870
rect 4066 13832 4122 13841
rect 4066 13767 4122 13776
rect 4250 13832 4252 13841
rect 4304 13832 4306 13841
rect 4250 13767 4306 13776
rect 4066 13560 4122 13569
rect 4066 13495 4122 13504
rect 4080 11082 4108 13495
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4158 13016 4214 13025
rect 4158 12951 4160 12960
rect 4212 12951 4214 12960
rect 4160 12922 4212 12928
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4172 10826 4200 12038
rect 4264 11014 4292 13262
rect 4356 12646 4384 14758
rect 4434 14719 4490 14728
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4448 12986 4476 14350
rect 4540 12986 4568 15506
rect 4632 15337 4660 15506
rect 4618 15328 4674 15337
rect 4618 15263 4674 15272
rect 4724 15178 4752 16068
rect 4804 16050 4856 16056
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 4816 15745 4844 16050
rect 4896 15904 4948 15910
rect 5000 15881 5028 16050
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 5092 15910 5120 15982
rect 5080 15904 5132 15910
rect 4896 15846 4948 15852
rect 4986 15872 5042 15881
rect 4802 15736 4858 15745
rect 4802 15671 4858 15680
rect 4908 15473 4936 15846
rect 5080 15846 5132 15852
rect 4986 15807 5042 15816
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 4894 15464 4950 15473
rect 4894 15399 4950 15408
rect 4986 15328 5042 15337
rect 4986 15263 5042 15272
rect 4724 15150 4844 15178
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4632 13530 4660 14894
rect 4724 14482 4752 15030
rect 4816 14906 4844 15150
rect 5000 15026 5028 15263
rect 5092 15201 5120 15642
rect 5078 15192 5134 15201
rect 5078 15127 5134 15136
rect 4988 15020 5040 15026
rect 5040 14980 5120 15008
rect 4988 14962 5040 14968
rect 4816 14878 5028 14906
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4894 14784 4950 14793
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4448 12782 4476 12922
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4632 12481 4660 13330
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4618 12472 4674 12481
rect 4618 12407 4674 12416
rect 4724 12306 4752 12786
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4618 12200 4674 12209
rect 4618 12135 4674 12144
rect 4632 11558 4660 12135
rect 4724 11762 4752 12242
rect 4816 12209 4844 14758
rect 4894 14719 4950 14728
rect 4908 14414 4936 14719
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4908 13870 4936 14350
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 4908 13326 4936 13806
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4908 12850 4936 13262
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4802 12200 4858 12209
rect 4802 12135 4858 12144
rect 4802 12064 4858 12073
rect 4802 11999 4858 12008
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4712 11212 4764 11218
rect 4816 11200 4844 11999
rect 4896 11280 4948 11286
rect 4896 11222 4948 11228
rect 4764 11172 4844 11200
rect 4712 11154 4764 11160
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4172 10798 4292 10826
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4080 10130 4108 10610
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4172 10010 4200 10678
rect 4080 9982 4200 10010
rect 4080 7018 4108 9982
rect 4264 9926 4292 10798
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4356 10180 4384 10406
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4436 10192 4488 10198
rect 4356 10152 4436 10180
rect 4632 10169 4660 10202
rect 4436 10134 4488 10140
rect 4618 10160 4674 10169
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4448 9722 4476 10134
rect 4618 10095 4674 10104
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 4618 9616 4674 9625
rect 4172 8430 4200 9590
rect 4618 9551 4674 9560
rect 4264 9132 4568 9160
rect 4264 8974 4292 9132
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 4264 8294 4292 8774
rect 4356 8634 4384 8978
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4448 8566 4476 8774
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4540 8430 4568 9132
rect 4632 9081 4660 9551
rect 4618 9072 4674 9081
rect 4618 9007 4674 9016
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 4080 6990 4200 7018
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4080 5234 4108 6802
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4172 5114 4200 6990
rect 4080 5086 4200 5114
rect 4080 3398 4108 5086
rect 4158 4312 4214 4321
rect 4158 4247 4214 4256
rect 4172 4214 4200 4247
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 4158 4040 4214 4049
rect 4158 3975 4160 3984
rect 4212 3975 4214 3984
rect 4160 3946 4212 3952
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 3974 2816 4030 2825
rect 3974 2751 4030 2760
rect 4172 2650 4200 3674
rect 4264 3233 4292 7754
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4436 6248 4488 6254
rect 4434 6216 4436 6225
rect 4488 6216 4490 6225
rect 4434 6151 4490 6160
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4356 4214 4384 6054
rect 4448 5914 4476 6054
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4448 4758 4476 5510
rect 4540 5166 4568 7686
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4632 5710 4660 7210
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4632 5234 4660 5646
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4724 5012 4752 11154
rect 4908 10577 4936 11222
rect 4894 10568 4950 10577
rect 4894 10503 4950 10512
rect 4908 8514 4936 10503
rect 5000 10470 5028 14878
rect 5092 13530 5120 14980
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 5078 12880 5134 12889
rect 5078 12815 5134 12824
rect 5092 11082 5120 12815
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 5092 10538 5120 11018
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 4986 9616 5042 9625
rect 4986 9551 5042 9560
rect 5080 9580 5132 9586
rect 5000 9450 5028 9551
rect 5080 9522 5132 9528
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 5092 9110 5120 9522
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 5078 8664 5134 8673
rect 5078 8599 5134 8608
rect 4816 8486 4936 8514
rect 4986 8528 5042 8537
rect 4816 7585 4844 8486
rect 4986 8463 5042 8472
rect 4896 8424 4948 8430
rect 4894 8392 4896 8401
rect 4948 8392 4950 8401
rect 5000 8362 5028 8463
rect 4894 8327 4950 8336
rect 4988 8356 5040 8362
rect 4802 7576 4858 7585
rect 4802 7511 4858 7520
rect 4908 7449 4936 8327
rect 4988 8298 5040 8304
rect 5092 8022 5120 8599
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 4894 7440 4950 7449
rect 4894 7375 4896 7384
rect 4948 7375 4950 7384
rect 4896 7346 4948 7352
rect 4908 6769 4936 7346
rect 5184 6882 5212 16118
rect 5368 15706 5396 17070
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5276 12889 5304 15438
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5368 15026 5396 15098
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5552 14906 5580 17206
rect 6288 17184 6316 19520
rect 6656 17218 6684 19520
rect 7024 17678 7052 19520
rect 7484 18086 7512 19520
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7852 17882 7880 19520
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7300 17338 7328 17478
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7380 17264 7432 17270
rect 7286 17232 7342 17241
rect 6656 17190 6868 17218
rect 6288 17156 6500 17184
rect 6368 17060 6420 17066
rect 6368 17002 6420 17008
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5644 14958 5672 16934
rect 5886 16892 6182 16912
rect 5942 16890 5966 16892
rect 6022 16890 6046 16892
rect 6102 16890 6126 16892
rect 5964 16838 5966 16890
rect 6028 16838 6040 16890
rect 6102 16838 6104 16890
rect 5942 16836 5966 16838
rect 6022 16836 6046 16838
rect 6102 16836 6126 16838
rect 5886 16816 6182 16836
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 5736 15042 5764 16186
rect 5828 15586 5856 16390
rect 5920 16114 5948 16390
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5886 15804 6182 15824
rect 5942 15802 5966 15804
rect 6022 15802 6046 15804
rect 6102 15802 6126 15804
rect 5964 15750 5966 15802
rect 6028 15750 6040 15802
rect 6102 15750 6104 15802
rect 5942 15748 5966 15750
rect 6022 15748 6046 15750
rect 6102 15748 6126 15750
rect 5886 15728 6182 15748
rect 6092 15632 6144 15638
rect 5828 15558 5948 15586
rect 6092 15574 6144 15580
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5828 15162 5856 15438
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 5736 15026 5856 15042
rect 5736 15020 5868 15026
rect 5736 15014 5816 15020
rect 5816 14962 5868 14968
rect 5460 14878 5580 14906
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5460 14521 5488 14878
rect 5920 14872 5948 15558
rect 6104 15026 6132 15574
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 5736 14844 5948 14872
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5446 14512 5502 14521
rect 5446 14447 5502 14456
rect 5552 14464 5580 14758
rect 5736 14464 5764 14844
rect 6104 14804 6132 14962
rect 5828 14776 6132 14804
rect 5828 14600 5856 14776
rect 5886 14716 6182 14736
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6126 14716
rect 5964 14662 5966 14714
rect 6028 14662 6040 14714
rect 6102 14662 6104 14714
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6126 14662
rect 5886 14640 6182 14660
rect 5828 14572 6040 14600
rect 5908 14476 5960 14482
rect 5356 14408 5408 14414
rect 5354 14376 5356 14385
rect 5460 14396 5488 14447
rect 5552 14436 5672 14464
rect 5736 14436 5908 14464
rect 5408 14376 5410 14385
rect 5460 14368 5580 14396
rect 5354 14311 5410 14320
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5262 12880 5318 12889
rect 5262 12815 5318 12824
rect 5262 12336 5318 12345
rect 5262 12271 5264 12280
rect 5316 12271 5318 12280
rect 5264 12242 5316 12248
rect 5368 11626 5396 13466
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5460 11937 5488 12718
rect 5446 11928 5502 11937
rect 5446 11863 5502 11872
rect 5356 11620 5408 11626
rect 5408 11580 5488 11608
rect 5356 11562 5408 11568
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5276 9586 5304 9998
rect 5368 9994 5396 10950
rect 5460 10554 5488 11580
rect 5552 11082 5580 14368
rect 5644 12753 5672 14436
rect 5908 14418 5960 14424
rect 6012 14362 6040 14572
rect 6288 14532 6316 16730
rect 6380 16561 6408 17002
rect 6366 16552 6422 16561
rect 6366 16487 6422 16496
rect 6472 15745 6500 17156
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6552 16992 6604 16998
rect 6550 16960 6552 16969
rect 6604 16960 6606 16969
rect 6550 16895 6606 16904
rect 6458 15736 6514 15745
rect 6458 15671 6514 15680
rect 6564 15586 6592 16895
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6380 15558 6592 15586
rect 6380 14958 6408 15558
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 5828 14334 6040 14362
rect 6104 14504 6316 14532
rect 5630 12744 5686 12753
rect 5630 12679 5686 12688
rect 5724 12640 5776 12646
rect 5722 12608 5724 12617
rect 5776 12608 5778 12617
rect 5722 12543 5778 12552
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5460 10526 5580 10554
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5460 10198 5488 10406
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5368 9042 5396 9930
rect 5552 9704 5580 10526
rect 5543 9676 5580 9704
rect 5543 9636 5571 9676
rect 5460 9608 5571 9636
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5262 8120 5318 8129
rect 5262 8055 5318 8064
rect 5276 7886 5304 8055
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5276 7546 5304 7822
rect 5354 7576 5410 7585
rect 5264 7540 5316 7546
rect 5354 7511 5410 7520
rect 5264 7482 5316 7488
rect 5368 7274 5396 7511
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5092 6854 5212 6882
rect 4988 6792 5040 6798
rect 4894 6760 4950 6769
rect 4988 6734 5040 6740
rect 4894 6695 4950 6704
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4816 5556 4844 6190
rect 4908 5914 4936 6598
rect 5000 5914 5028 6734
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4896 5568 4948 5574
rect 4816 5528 4896 5556
rect 4896 5510 4948 5516
rect 4802 5400 4858 5409
rect 4802 5335 4804 5344
rect 4856 5335 4858 5344
rect 4804 5306 4856 5312
rect 4908 5166 4936 5510
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4540 4984 4752 5012
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4540 4604 4568 4984
rect 4816 4758 4844 5034
rect 5000 4826 5028 5646
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4448 4576 4568 4604
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 4448 3924 4476 4576
rect 4710 4448 4766 4457
rect 4710 4383 4766 4392
rect 4356 3896 4476 3924
rect 4250 3224 4306 3233
rect 4250 3159 4306 3168
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 3988 1630 4016 2314
rect 4160 2304 4212 2310
rect 4264 2292 4292 2994
rect 4356 2446 4384 3896
rect 4528 3528 4580 3534
rect 4526 3496 4528 3505
rect 4580 3496 4582 3505
rect 4436 3460 4488 3466
rect 4526 3431 4582 3440
rect 4436 3402 4488 3408
rect 4448 2922 4476 3402
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4632 2990 4660 3334
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 4212 2264 4292 2292
rect 4342 2272 4398 2281
rect 4160 2246 4212 2252
rect 4342 2207 4398 2216
rect 3976 1624 4028 1630
rect 3976 1566 4028 1572
rect 4356 480 4384 2207
rect 4448 1834 4476 2314
rect 4540 2310 4568 2926
rect 4618 2544 4674 2553
rect 4618 2479 4620 2488
rect 4672 2479 4674 2488
rect 4620 2450 4672 2456
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4436 1828 4488 1834
rect 4436 1770 4488 1776
rect 4724 480 4752 4383
rect 4802 4312 4858 4321
rect 4802 4247 4858 4256
rect 4986 4312 5042 4321
rect 4986 4247 5042 4256
rect 4816 2854 4844 4247
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4908 2650 4936 4014
rect 5000 3618 5028 4247
rect 5092 3738 5120 6854
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5262 6760 5318 6769
rect 5184 5098 5212 6734
rect 5262 6695 5318 6704
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5000 3590 5120 3618
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5000 1601 5028 3402
rect 5092 3194 5120 3590
rect 5184 3534 5212 4218
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5184 2446 5212 3470
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5276 2292 5304 6695
rect 5460 5846 5488 9608
rect 5644 8906 5672 11562
rect 5736 10849 5764 12378
rect 5722 10840 5778 10849
rect 5722 10775 5778 10784
rect 5828 10266 5856 14334
rect 6104 13841 6132 14504
rect 6380 13938 6408 14894
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6276 13864 6328 13870
rect 6090 13832 6146 13841
rect 6276 13806 6328 13812
rect 6090 13767 6146 13776
rect 5886 13628 6182 13648
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6126 13628
rect 5964 13574 5966 13626
rect 6028 13574 6040 13626
rect 6102 13574 6104 13626
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6126 13574
rect 5886 13552 6182 13572
rect 5886 12540 6182 12560
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6126 12540
rect 5964 12486 5966 12538
rect 6028 12486 6040 12538
rect 6102 12486 6104 12538
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6126 12486
rect 5886 12464 6182 12484
rect 5886 11452 6182 11472
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6126 11452
rect 5964 11398 5966 11450
rect 6028 11398 6040 11450
rect 6102 11398 6104 11450
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6126 11398
rect 5886 11376 6182 11396
rect 6288 10810 6316 13806
rect 6472 13802 6500 15438
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6564 14550 6592 15302
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6656 14006 6684 16526
rect 6748 14278 6776 17070
rect 6840 15314 6868 17190
rect 7380 17206 7432 17212
rect 7286 17167 7342 17176
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6932 15706 6960 16390
rect 7024 16250 7052 17070
rect 7300 16794 7328 17167
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7194 16688 7250 16697
rect 7194 16623 7196 16632
rect 7248 16623 7250 16632
rect 7196 16594 7248 16600
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7116 15910 7144 16186
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7104 15904 7156 15910
rect 7010 15872 7066 15881
rect 7104 15846 7156 15852
rect 7010 15807 7066 15816
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 7024 15434 7052 15807
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 6840 15286 6960 15314
rect 6826 15192 6882 15201
rect 6826 15127 6882 15136
rect 6840 14657 6868 15127
rect 6932 15065 6960 15286
rect 6918 15056 6974 15065
rect 6918 14991 6974 15000
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6826 14648 6882 14657
rect 6826 14583 6882 14592
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6460 13796 6512 13802
rect 6460 13738 6512 13744
rect 6380 13530 6408 13738
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6472 12442 6500 13738
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6368 12368 6420 12374
rect 6564 12322 6592 13874
rect 6840 13870 6868 14350
rect 6828 13864 6880 13870
rect 6826 13832 6828 13841
rect 6880 13832 6882 13841
rect 6826 13767 6882 13776
rect 6840 13326 6868 13767
rect 6932 13530 6960 14826
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 7024 13274 7052 14214
rect 7116 13530 7144 15438
rect 7208 14793 7236 16050
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7300 15337 7328 15846
rect 7286 15328 7342 15337
rect 7286 15263 7342 15272
rect 7392 15162 7420 17206
rect 7576 17066 7604 17478
rect 8116 17264 8168 17270
rect 8116 17206 8168 17212
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7472 16108 7524 16114
rect 7576 16096 7604 16730
rect 7524 16068 7604 16096
rect 7472 16050 7524 16056
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7484 15570 7512 15914
rect 7472 15564 7524 15570
rect 7472 15506 7524 15512
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7288 14816 7340 14822
rect 7194 14784 7250 14793
rect 7288 14758 7340 14764
rect 7194 14719 7250 14728
rect 7300 14618 7328 14758
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7392 13802 7420 15098
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7102 13424 7158 13433
rect 7102 13359 7104 13368
rect 7156 13359 7158 13368
rect 7104 13330 7156 13336
rect 6644 13184 6696 13190
rect 6642 13152 6644 13161
rect 6696 13152 6698 13161
rect 6642 13087 6698 13096
rect 6368 12310 6420 12316
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 5886 10364 6182 10384
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6126 10364
rect 5964 10310 5966 10362
rect 6028 10310 6040 10362
rect 6102 10310 6104 10362
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6126 10310
rect 5886 10288 6182 10308
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 6288 10198 6316 10746
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6276 9580 6328 9586
rect 5828 9540 6276 9568
rect 5828 9042 5856 9540
rect 6276 9522 6328 9528
rect 6274 9344 6330 9353
rect 5886 9276 6182 9296
rect 6274 9279 6330 9288
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6126 9276
rect 5964 9222 5966 9274
rect 6028 9222 6040 9274
rect 6102 9222 6104 9274
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6126 9222
rect 5886 9200 6182 9220
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 6288 8537 6316 9279
rect 6380 9217 6408 12310
rect 6472 12294 6592 12322
rect 6472 9761 6500 12294
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6564 11218 6592 12174
rect 6656 11694 6684 13087
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6564 10713 6592 10746
rect 6550 10704 6606 10713
rect 6550 10639 6606 10648
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6458 9752 6514 9761
rect 6564 9722 6592 10202
rect 6458 9687 6514 9696
rect 6552 9716 6604 9722
rect 6366 9208 6422 9217
rect 6366 9143 6422 9152
rect 6274 8528 6330 8537
rect 5644 8486 5856 8514
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5448 5840 5500 5846
rect 5552 5828 5580 8298
rect 5644 8129 5672 8486
rect 5828 8412 5856 8486
rect 6000 8492 6052 8498
rect 6274 8463 6330 8472
rect 6368 8492 6420 8498
rect 6000 8434 6052 8440
rect 6472 8480 6500 9687
rect 6552 9658 6604 9664
rect 6748 9518 6776 12242
rect 6840 11762 6868 13262
rect 7024 13246 7144 13274
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 12442 6960 12582
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6840 11150 6868 11698
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6840 10674 6868 11086
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 7024 9450 7052 12038
rect 7116 11558 7144 13246
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7208 12442 7236 13126
rect 7380 12776 7432 12782
rect 7300 12736 7380 12764
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7194 11792 7250 11801
rect 7194 11727 7250 11736
rect 7208 11626 7236 11727
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7300 9654 7328 12736
rect 7380 12718 7432 12724
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7392 11286 7420 12378
rect 7484 12186 7512 15370
rect 7576 15366 7604 15914
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7576 12345 7604 14962
rect 7668 12918 7696 17138
rect 7932 16992 7984 16998
rect 7932 16934 7984 16940
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7760 15609 7788 16050
rect 7746 15600 7802 15609
rect 7746 15535 7802 15544
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7746 15328 7802 15337
rect 7746 15263 7802 15272
rect 7760 14958 7788 15263
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7852 14482 7880 15438
rect 7944 15026 7972 16934
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 8036 15473 8064 15982
rect 8128 15502 8156 17206
rect 8220 16674 8248 18158
rect 8312 17746 8340 19520
rect 8680 19502 8715 19520
rect 8687 19394 8715 19502
rect 8687 19366 8800 19394
rect 8772 18222 8800 19366
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8668 17604 8720 17610
rect 8668 17546 8720 17552
rect 8352 17436 8648 17456
rect 8408 17434 8432 17436
rect 8488 17434 8512 17436
rect 8568 17434 8592 17436
rect 8430 17382 8432 17434
rect 8494 17382 8506 17434
rect 8568 17382 8570 17434
rect 8408 17380 8432 17382
rect 8488 17380 8512 17382
rect 8568 17380 8592 17382
rect 8352 17360 8648 17380
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 16794 8432 16934
rect 8680 16794 8708 17546
rect 8956 16794 8984 17682
rect 9048 17513 9076 19520
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9034 17504 9090 17513
rect 9034 17439 9090 17448
rect 9140 17134 9168 18362
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9128 17128 9180 17134
rect 9128 17070 9180 17076
rect 9218 17096 9274 17105
rect 9218 17031 9274 17040
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8944 16788 8996 16794
rect 9232 16776 9260 17031
rect 8944 16730 8996 16736
rect 9140 16748 9260 16776
rect 8220 16646 8708 16674
rect 8680 16640 8708 16646
rect 9036 16652 9088 16658
rect 8680 16612 8800 16640
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8576 16584 8628 16590
rect 8628 16544 8708 16572
rect 8576 16526 8628 16532
rect 8220 16454 8248 16526
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8352 16348 8648 16368
rect 8408 16346 8432 16348
rect 8488 16346 8512 16348
rect 8568 16346 8592 16348
rect 8430 16294 8432 16346
rect 8494 16294 8506 16346
rect 8568 16294 8570 16346
rect 8408 16292 8432 16294
rect 8488 16292 8512 16294
rect 8568 16292 8592 16294
rect 8206 16280 8262 16289
rect 8352 16272 8648 16292
rect 8206 16215 8262 16224
rect 8220 15722 8248 16215
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8312 15722 8340 15982
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8220 15694 8340 15722
rect 8116 15496 8168 15502
rect 8022 15464 8078 15473
rect 8116 15438 8168 15444
rect 8022 15399 8078 15408
rect 8116 15360 8168 15366
rect 8496 15348 8524 15846
rect 8680 15722 8708 16544
rect 8772 15881 8800 16612
rect 9036 16594 9088 16600
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8864 16250 8892 16390
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8758 15872 8814 15881
rect 8942 15872 8998 15881
rect 8814 15830 8892 15858
rect 8758 15807 8814 15816
rect 8680 15694 8800 15722
rect 8668 15564 8720 15570
rect 8220 15337 8524 15348
rect 8116 15302 8168 15308
rect 8206 15328 8524 15337
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 7840 14476 7892 14482
rect 7892 14436 7972 14464
rect 7840 14418 7892 14424
rect 7748 13796 7800 13802
rect 7748 13738 7800 13744
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7760 12764 7788 13738
rect 7944 13705 7972 14436
rect 7930 13696 7986 13705
rect 7930 13631 7986 13640
rect 7840 13524 7892 13530
rect 7892 13484 7972 13512
rect 7840 13466 7892 13472
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7852 13161 7880 13194
rect 7838 13152 7894 13161
rect 7838 13087 7894 13096
rect 7944 12850 7972 13484
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7668 12736 7788 12764
rect 7562 12336 7618 12345
rect 7562 12271 7618 12280
rect 7484 12158 7604 12186
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7484 10713 7512 12038
rect 7576 11393 7604 12158
rect 7668 11626 7696 12736
rect 7852 12424 7880 12786
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7944 12617 7972 12650
rect 7930 12608 7986 12617
rect 8036 12594 8064 14758
rect 8128 14006 8156 15302
rect 8262 15320 8524 15328
rect 8588 15524 8668 15552
rect 8588 15348 8616 15524
rect 8668 15506 8720 15512
rect 8588 15320 8708 15348
rect 8772 15337 8800 15694
rect 8864 15570 8892 15830
rect 8942 15807 8998 15816
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 8852 15428 8904 15434
rect 8852 15370 8904 15376
rect 8206 15263 8262 15272
rect 8352 15260 8648 15280
rect 8408 15258 8432 15260
rect 8488 15258 8512 15260
rect 8568 15258 8592 15260
rect 8430 15206 8432 15258
rect 8494 15206 8506 15258
rect 8568 15206 8570 15258
rect 8408 15204 8432 15206
rect 8488 15204 8512 15206
rect 8568 15204 8592 15206
rect 8206 15192 8262 15201
rect 8352 15184 8648 15204
rect 8206 15127 8262 15136
rect 8220 14804 8248 15127
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8680 14906 8708 15320
rect 8758 15328 8814 15337
rect 8758 15263 8814 15272
rect 8864 14940 8892 15370
rect 8956 15094 8984 15807
rect 8944 15088 8996 15094
rect 8944 15030 8996 15036
rect 8864 14912 8984 14940
rect 8496 14804 8524 14894
rect 8680 14878 8800 14906
rect 8220 14776 8524 14804
rect 8668 14816 8720 14822
rect 8574 14784 8630 14793
rect 8668 14758 8720 14764
rect 8574 14719 8630 14728
rect 8206 14512 8262 14521
rect 8206 14447 8208 14456
rect 8260 14447 8262 14456
rect 8208 14418 8260 14424
rect 8588 14346 8616 14719
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8220 14056 8248 14214
rect 8352 14172 8648 14192
rect 8408 14170 8432 14172
rect 8488 14170 8512 14172
rect 8568 14170 8592 14172
rect 8430 14118 8432 14170
rect 8494 14118 8506 14170
rect 8568 14118 8570 14170
rect 8408 14116 8432 14118
rect 8488 14116 8512 14118
rect 8568 14116 8592 14118
rect 8352 14096 8648 14116
rect 8220 14028 8340 14056
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 8128 13433 8156 13942
rect 8206 13696 8262 13705
rect 8206 13631 8262 13640
rect 8220 13530 8248 13631
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 8114 13424 8170 13433
rect 8312 13394 8340 14028
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8484 13932 8536 13938
rect 8484 13874 8536 13880
rect 8496 13841 8524 13874
rect 8482 13832 8538 13841
rect 8482 13767 8538 13776
rect 8588 13705 8616 13942
rect 8680 13841 8708 14758
rect 8666 13832 8722 13841
rect 8666 13767 8722 13776
rect 8574 13696 8630 13705
rect 8574 13631 8630 13640
rect 8114 13359 8170 13368
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8352 13084 8648 13104
rect 8408 13082 8432 13084
rect 8488 13082 8512 13084
rect 8568 13082 8592 13084
rect 8430 13030 8432 13082
rect 8494 13030 8506 13082
rect 8568 13030 8570 13082
rect 8408 13028 8432 13030
rect 8488 13028 8512 13030
rect 8568 13028 8592 13030
rect 8352 13008 8648 13028
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8392 12912 8444 12918
rect 8392 12854 8444 12860
rect 8208 12640 8260 12646
rect 8036 12566 8156 12594
rect 8208 12582 8260 12588
rect 7930 12543 7986 12552
rect 7852 12396 8064 12424
rect 7852 12238 7880 12396
rect 7930 12336 7986 12345
rect 7930 12271 7986 12280
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7748 12096 7800 12102
rect 7852 12073 7880 12174
rect 7748 12038 7800 12044
rect 7838 12064 7894 12073
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7562 11384 7618 11393
rect 7562 11319 7618 11328
rect 7470 10704 7526 10713
rect 7470 10639 7526 10648
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6828 9444 6880 9450
rect 6828 9386 6880 9392
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6420 8452 6500 8480
rect 6368 8434 6420 8440
rect 5908 8424 5960 8430
rect 5722 8392 5778 8401
rect 5828 8384 5908 8412
rect 5908 8366 5960 8372
rect 5722 8327 5778 8336
rect 5630 8120 5686 8129
rect 5630 8055 5686 8064
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5644 7546 5672 7890
rect 5736 7886 5764 8327
rect 6012 8276 6040 8434
rect 6184 8356 6236 8362
rect 6236 8316 6316 8344
rect 6184 8298 6236 8304
rect 5828 8248 6040 8276
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5828 7721 5856 8248
rect 5886 8188 6182 8208
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6126 8188
rect 5964 8134 5966 8186
rect 6028 8134 6040 8186
rect 6102 8134 6104 8186
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6126 8134
rect 5886 8112 6182 8132
rect 6288 8129 6316 8316
rect 6368 8288 6420 8294
rect 6656 8242 6684 9318
rect 6840 8906 6868 9386
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6932 8838 6960 9318
rect 7116 9042 7144 9522
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6828 8424 6880 8430
rect 6734 8392 6790 8401
rect 6828 8366 6880 8372
rect 6734 8327 6790 8336
rect 6368 8230 6420 8236
rect 6274 8120 6330 8129
rect 6380 8090 6408 8230
rect 6472 8214 6684 8242
rect 6274 8055 6330 8064
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6000 8016 6052 8022
rect 6052 7976 6316 8004
rect 6000 7958 6052 7964
rect 5814 7712 5870 7721
rect 5814 7647 5870 7656
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5908 7472 5960 7478
rect 5736 7432 5908 7460
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5644 7206 5672 7278
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5632 6724 5684 6730
rect 5736 6712 5764 7432
rect 5908 7414 5960 7420
rect 6288 7206 6316 7976
rect 6276 7200 6328 7206
rect 6472 7177 6500 8214
rect 6748 8106 6776 8327
rect 6564 8078 6776 8106
rect 6276 7142 6328 7148
rect 6458 7168 6514 7177
rect 5886 7100 6182 7120
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6126 7100
rect 5964 7046 5966 7098
rect 6028 7046 6040 7098
rect 6102 7046 6104 7098
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6126 7046
rect 5886 7024 6182 7044
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5684 6684 5764 6712
rect 5632 6666 5684 6672
rect 5828 6633 5856 6734
rect 5814 6624 5870 6633
rect 6288 6610 6316 7142
rect 6458 7103 6514 7112
rect 5814 6559 5870 6568
rect 6196 6582 6316 6610
rect 5908 6384 5960 6390
rect 5828 6344 5908 6372
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5736 6089 5764 6190
rect 5828 6118 5856 6344
rect 6196 6361 6224 6582
rect 6276 6384 6328 6390
rect 5908 6326 5960 6332
rect 6182 6352 6238 6361
rect 6276 6326 6328 6332
rect 6182 6287 6238 6296
rect 5816 6112 5868 6118
rect 5722 6080 5778 6089
rect 5816 6054 5868 6060
rect 5722 6015 5778 6024
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 6288 5846 6316 6326
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5953 6408 6054
rect 6366 5944 6422 5953
rect 6366 5879 6422 5888
rect 6276 5840 6328 5846
rect 5448 5782 5500 5788
rect 5543 5800 6132 5828
rect 5448 5704 5500 5710
rect 5354 5672 5410 5681
rect 5543 5692 5571 5800
rect 5500 5664 5571 5692
rect 5632 5704 5684 5710
rect 5448 5646 5500 5652
rect 5632 5646 5684 5652
rect 5722 5672 5778 5681
rect 5354 5607 5356 5616
rect 5408 5607 5410 5616
rect 5356 5578 5408 5584
rect 5354 5400 5410 5409
rect 5354 5335 5410 5344
rect 5368 5001 5396 5335
rect 5644 5114 5672 5646
rect 5722 5607 5778 5616
rect 5460 5086 5672 5114
rect 5354 4992 5410 5001
rect 5354 4927 5410 4936
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5368 4690 5396 4762
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5368 4010 5396 4490
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5368 3505 5396 3538
rect 5354 3496 5410 3505
rect 5354 3431 5410 3440
rect 5354 3224 5410 3233
rect 5354 3159 5410 3168
rect 5368 2854 5396 3159
rect 5460 3058 5488 5086
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5552 4282 5580 4966
rect 5644 4826 5672 4966
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5644 4282 5672 4626
rect 5736 4570 5764 5607
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 5816 5092 5868 5098
rect 6012 5080 6040 5510
rect 6104 5370 6132 5800
rect 6276 5782 6328 5788
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6012 5052 6316 5080
rect 5816 5034 5868 5040
rect 5828 4690 5856 5034
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 6288 4690 6316 5052
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 5736 4542 5948 4570
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5552 3058 5580 4082
rect 5736 3738 5764 4422
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5724 3528 5776 3534
rect 5644 3488 5724 3516
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5446 2816 5502 2825
rect 5446 2751 5502 2760
rect 5354 2408 5410 2417
rect 5460 2378 5488 2751
rect 5644 2689 5672 3488
rect 5724 3470 5776 3476
rect 5828 3210 5856 4422
rect 5920 4010 5948 4542
rect 6274 4040 6330 4049
rect 5908 4004 5960 4010
rect 6274 3975 6330 3984
rect 5908 3946 5960 3952
rect 5886 3836 6182 3856
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 5736 3182 5856 3210
rect 5736 2990 5764 3182
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5630 2680 5686 2689
rect 5828 2650 5856 3062
rect 5920 2990 5948 3606
rect 6104 3398 6132 3606
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6196 3210 6224 3538
rect 6288 3398 6316 3975
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6196 3182 6316 3210
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 5630 2615 5686 2624
rect 5816 2644 5868 2650
rect 5644 2514 5672 2615
rect 6288 2632 6316 3182
rect 6380 3058 6408 5879
rect 6472 5574 6500 6122
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 5816 2586 5868 2592
rect 6196 2604 6316 2632
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5354 2343 5410 2352
rect 5448 2372 5500 2378
rect 5184 2264 5304 2292
rect 4986 1592 5042 1601
rect 4986 1527 5042 1536
rect 5184 480 5212 2264
rect 5368 1494 5396 2343
rect 5448 2314 5500 2320
rect 6000 1896 6052 1902
rect 6000 1838 6052 1844
rect 5356 1488 5408 1494
rect 5356 1430 5408 1436
rect 5538 1184 5594 1193
rect 5538 1119 5594 1128
rect 5552 480 5580 1119
rect 6012 480 6040 1838
rect 6196 1057 6224 2604
rect 6472 2446 6500 5034
rect 6564 4128 6592 8078
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6748 7721 6776 7958
rect 6734 7712 6790 7721
rect 6734 7647 6790 7656
rect 6642 7440 6698 7449
rect 6642 7375 6698 7384
rect 6656 7342 6684 7375
rect 6840 7342 6868 8366
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 8090 6960 8230
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6835 7336 6887 7342
rect 6835 7278 6887 7284
rect 6736 6996 6788 7002
rect 6736 6938 6788 6944
rect 6642 6488 6698 6497
rect 6642 6423 6698 6432
rect 6656 5137 6684 6423
rect 6748 5642 6776 6938
rect 6840 6254 6868 7278
rect 6932 6866 6960 7890
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6932 6633 6960 6666
rect 6918 6624 6974 6633
rect 6918 6559 6974 6568
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 7024 6118 7052 8978
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 6662 7144 8774
rect 7208 8362 7236 8842
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7208 7002 7236 8298
rect 7300 7585 7328 9386
rect 7392 7857 7420 10202
rect 7470 10024 7526 10033
rect 7470 9959 7526 9968
rect 7378 7848 7434 7857
rect 7378 7783 7434 7792
rect 7286 7576 7342 7585
rect 7286 7511 7342 7520
rect 7484 7460 7512 9959
rect 7576 8537 7604 11319
rect 7562 8528 7618 8537
rect 7562 8463 7618 8472
rect 7668 7585 7696 11562
rect 7760 10266 7788 12038
rect 7838 11999 7894 12008
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7852 10198 7880 11834
rect 7944 10742 7972 12271
rect 8036 12170 8064 12396
rect 8024 12164 8076 12170
rect 8024 12106 8076 12112
rect 8128 11778 8156 12566
rect 8220 12374 8248 12582
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8312 12238 8340 12854
rect 8404 12782 8432 12854
rect 8392 12776 8444 12782
rect 8772 12764 8800 14878
rect 8852 14816 8904 14822
rect 8956 14793 8984 14912
rect 8852 14758 8904 14764
rect 8942 14784 8998 14793
rect 8864 14249 8892 14758
rect 8942 14719 8998 14728
rect 8942 14376 8998 14385
rect 8942 14311 8998 14320
rect 8956 14278 8984 14311
rect 8944 14272 8996 14278
rect 8850 14240 8906 14249
rect 8944 14214 8996 14220
rect 8850 14175 8906 14184
rect 8942 13968 8998 13977
rect 8942 13903 8998 13912
rect 8850 13696 8906 13705
rect 8850 13631 8906 13640
rect 8864 13326 8892 13631
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8956 12832 8984 13903
rect 9048 12850 9076 16594
rect 9140 16114 9168 16748
rect 9218 16688 9274 16697
rect 9218 16623 9220 16632
rect 9272 16623 9274 16632
rect 9220 16594 9272 16600
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 9140 15722 9168 15914
rect 9232 15881 9260 15982
rect 9218 15872 9274 15881
rect 9218 15807 9274 15816
rect 9140 15694 9260 15722
rect 9232 15434 9260 15694
rect 9324 15688 9352 16526
rect 9416 15881 9444 17750
rect 9508 16561 9536 19520
rect 9876 18170 9904 19520
rect 9680 18148 9732 18154
rect 9876 18142 10180 18170
rect 9680 18090 9732 18096
rect 9586 17368 9642 17377
rect 9586 17303 9642 17312
rect 9600 16998 9628 17303
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9494 16552 9550 16561
rect 9494 16487 9550 16496
rect 9586 16280 9642 16289
rect 9692 16266 9720 18090
rect 9954 17368 10010 17377
rect 9954 17303 10010 17312
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9784 16697 9812 16934
rect 9770 16688 9826 16697
rect 9770 16623 9826 16632
rect 9692 16250 9812 16266
rect 9692 16244 9824 16250
rect 9692 16238 9772 16244
rect 9586 16215 9642 16224
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9402 15872 9458 15881
rect 9402 15807 9458 15816
rect 9324 15660 9444 15688
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9128 15360 9180 15366
rect 9126 15328 9128 15337
rect 9180 15328 9182 15337
rect 9126 15263 9182 15272
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9126 14512 9182 14521
rect 9126 14447 9182 14456
rect 9140 12986 9168 14447
rect 9232 13161 9260 14962
rect 9324 14482 9352 15506
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9416 14074 9444 15660
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9324 13802 9352 14010
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9218 13152 9274 13161
rect 9218 13087 9274 13096
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 8392 12718 8444 12724
rect 8496 12736 8800 12764
rect 8864 12804 8984 12832
rect 9036 12844 9088 12850
rect 8496 12442 8524 12736
rect 8666 12472 8722 12481
rect 8484 12436 8536 12442
rect 8864 12442 8892 12804
rect 9036 12786 9088 12792
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 8666 12407 8722 12416
rect 8852 12436 8904 12442
rect 8484 12378 8536 12384
rect 8680 12374 8708 12407
rect 8852 12378 8904 12384
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8588 12186 8616 12242
rect 8772 12186 8800 12242
rect 8588 12158 8800 12186
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11937 8248 12038
rect 8352 11996 8648 12016
rect 8408 11994 8432 11996
rect 8488 11994 8512 11996
rect 8568 11994 8592 11996
rect 8430 11942 8432 11994
rect 8494 11942 8506 11994
rect 8568 11942 8570 11994
rect 8408 11940 8432 11942
rect 8488 11940 8512 11942
rect 8568 11940 8592 11942
rect 8206 11928 8262 11937
rect 8352 11920 8648 11940
rect 8206 11863 8262 11872
rect 8128 11750 8524 11778
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 11286 8248 11494
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8312 11132 8340 11630
rect 8496 11626 8524 11750
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8220 11104 8340 11132
rect 8760 11144 8812 11150
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 8036 10606 8064 11018
rect 8114 10840 8170 10849
rect 8114 10775 8170 10784
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 8128 10198 8156 10775
rect 8220 10606 8248 11104
rect 8760 11086 8812 11092
rect 8352 10908 8648 10928
rect 8408 10906 8432 10908
rect 8488 10906 8512 10908
rect 8568 10906 8592 10908
rect 8430 10854 8432 10906
rect 8494 10854 8506 10906
rect 8568 10854 8570 10906
rect 8408 10852 8432 10854
rect 8488 10852 8512 10854
rect 8568 10852 8592 10854
rect 8352 10832 8648 10852
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 7840 10192 7892 10198
rect 7840 10134 7892 10140
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8114 10024 8170 10033
rect 8114 9959 8170 9968
rect 7746 9752 7802 9761
rect 7746 9687 7802 9696
rect 7760 9586 7788 9687
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7932 8832 7984 8838
rect 8036 8809 8064 9590
rect 7932 8774 7984 8780
rect 8022 8800 8078 8809
rect 7840 8628 7892 8634
rect 7760 8588 7840 8616
rect 7760 8090 7788 8588
rect 7840 8570 7892 8576
rect 7944 8378 7972 8774
rect 8022 8735 8078 8744
rect 8022 8528 8078 8537
rect 8022 8463 8024 8472
rect 8076 8463 8078 8472
rect 8024 8434 8076 8440
rect 7852 8350 7972 8378
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7654 7576 7710 7585
rect 7564 7540 7616 7546
rect 7654 7511 7710 7520
rect 7564 7482 7616 7488
rect 7300 7432 7512 7460
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7300 6338 7328 7432
rect 7576 7274 7604 7482
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7392 7177 7420 7210
rect 7378 7168 7434 7177
rect 7562 7168 7618 7177
rect 7378 7103 7434 7112
rect 7484 7126 7562 7154
rect 7208 6310 7328 6338
rect 7012 6112 7064 6118
rect 6826 6080 6882 6089
rect 7012 6054 7064 6060
rect 6826 6015 6882 6024
rect 6840 5760 6868 6015
rect 6840 5732 6875 5760
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6847 5386 6875 5732
rect 7024 5692 7052 6054
rect 7208 5760 7236 6310
rect 7380 6248 7432 6254
rect 6840 5358 6875 5386
rect 6932 5664 7052 5692
rect 7096 5732 7236 5760
rect 7300 6208 7380 6236
rect 6642 5128 6698 5137
rect 6642 5063 6698 5072
rect 6736 4752 6788 4758
rect 6736 4694 6788 4700
rect 6564 4100 6684 4128
rect 6550 4040 6606 4049
rect 6550 3975 6552 3984
rect 6604 3975 6606 3984
rect 6552 3946 6604 3952
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6564 3194 6592 3470
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 6276 2304 6328 2310
rect 6656 2292 6684 4100
rect 6748 3913 6776 4694
rect 6840 4457 6868 5358
rect 6826 4448 6882 4457
rect 6826 4383 6882 4392
rect 6932 4146 6960 5664
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7024 5098 7052 5510
rect 7096 5386 7124 5732
rect 7096 5358 7144 5386
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 7024 4457 7052 4626
rect 7010 4448 7066 4457
rect 7010 4383 7066 4392
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6734 3904 6790 3913
rect 6734 3839 6790 3848
rect 6748 3466 6776 3839
rect 6736 3460 6788 3466
rect 6736 3402 6788 3408
rect 6734 3360 6790 3369
rect 6734 3295 6790 3304
rect 6748 2825 6776 3295
rect 6840 3194 6868 3946
rect 6932 3534 6960 4082
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6920 3528 6972 3534
rect 7024 3516 7052 3878
rect 7116 3584 7144 5358
rect 7300 5216 7328 6208
rect 7380 6190 7432 6196
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7392 5234 7420 5646
rect 7208 5188 7328 5216
rect 7380 5228 7432 5234
rect 7208 5098 7236 5188
rect 7380 5170 7432 5176
rect 7286 5128 7342 5137
rect 7196 5092 7248 5098
rect 7286 5063 7342 5072
rect 7380 5092 7432 5098
rect 7196 5034 7248 5040
rect 7194 4992 7250 5001
rect 7194 4927 7250 4936
rect 7208 3738 7236 4927
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7116 3556 7236 3584
rect 7024 3488 7144 3516
rect 6920 3470 6972 3476
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7024 2854 7052 2926
rect 6920 2848 6972 2854
rect 6734 2816 6790 2825
rect 6920 2790 6972 2796
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 6734 2751 6790 2760
rect 6826 2680 6882 2689
rect 6826 2615 6882 2624
rect 6276 2246 6328 2252
rect 6380 2264 6684 2292
rect 6288 1698 6316 2246
rect 6276 1692 6328 1698
rect 6276 1634 6328 1640
rect 6182 1048 6238 1057
rect 6182 983 6238 992
rect 6380 480 6408 2264
rect 6840 480 6868 2615
rect 6932 2496 6960 2790
rect 7012 2508 7064 2514
rect 6932 2468 7012 2496
rect 7012 2450 7064 2456
rect 7116 1290 7144 3488
rect 7104 1284 7156 1290
rect 7104 1226 7156 1232
rect 7208 480 7236 3556
rect 7300 3058 7328 5063
rect 7380 5034 7432 5040
rect 7392 3534 7420 5034
rect 7484 4196 7512 7126
rect 7562 7103 7618 7112
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7576 6254 7604 6938
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 6254 7696 6734
rect 7760 6338 7788 7890
rect 7852 7546 7880 8350
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7944 7857 7972 8230
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 7930 7848 7986 7857
rect 8036 7818 8064 7890
rect 7930 7783 7986 7792
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7932 7200 7984 7206
rect 8128 7177 8156 9959
rect 8220 8616 8248 10202
rect 8312 10130 8340 10542
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8772 10044 8800 11086
rect 8864 10266 8892 12378
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8852 10056 8904 10062
rect 8772 10016 8852 10044
rect 8852 9998 8904 10004
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8352 9820 8648 9840
rect 8408 9818 8432 9820
rect 8488 9818 8512 9820
rect 8568 9818 8592 9820
rect 8430 9766 8432 9818
rect 8494 9766 8506 9818
rect 8568 9766 8570 9818
rect 8408 9764 8432 9766
rect 8488 9764 8512 9766
rect 8568 9764 8592 9766
rect 8352 9744 8648 9764
rect 8404 9540 8616 9568
rect 8404 9450 8432 9540
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8588 8906 8616 9540
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8668 8832 8720 8838
rect 8772 8809 8800 8978
rect 8668 8774 8720 8780
rect 8758 8800 8814 8809
rect 8352 8732 8648 8752
rect 8408 8730 8432 8732
rect 8488 8730 8512 8732
rect 8568 8730 8592 8732
rect 8430 8678 8432 8730
rect 8494 8678 8506 8730
rect 8568 8678 8570 8730
rect 8408 8676 8432 8678
rect 8488 8676 8512 8678
rect 8568 8676 8592 8678
rect 8352 8656 8648 8676
rect 8220 8588 8340 8616
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8220 8090 8248 8298
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8312 7970 8340 8588
rect 8680 8498 8708 8774
rect 8758 8735 8814 8744
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8404 8090 8432 8434
rect 8864 8378 8892 9862
rect 8680 8350 8892 8378
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8680 8022 8708 8350
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8220 7942 8340 7970
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 7932 7142 7984 7148
rect 8114 7168 8170 7177
rect 7944 6848 7972 7142
rect 8114 7103 8170 7112
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8128 6905 8156 6938
rect 7935 6820 7972 6848
rect 8114 6896 8170 6905
rect 8114 6831 8170 6840
rect 7935 6644 7963 6820
rect 8220 6780 8248 7942
rect 8772 7868 8800 8230
rect 8852 7880 8904 7886
rect 8772 7840 8852 7868
rect 8852 7822 8904 7828
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8352 7644 8648 7664
rect 8408 7642 8432 7644
rect 8488 7642 8512 7644
rect 8568 7642 8592 7644
rect 8430 7590 8432 7642
rect 8494 7590 8506 7642
rect 8568 7590 8570 7642
rect 8408 7588 8432 7590
rect 8488 7588 8512 7590
rect 8568 7588 8592 7590
rect 8352 7568 8648 7588
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8128 6752 8248 6780
rect 7935 6616 7972 6644
rect 7944 6458 7972 6616
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7760 6310 7972 6338
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7668 5710 7696 6190
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7760 5953 7788 6122
rect 7746 5944 7802 5953
rect 7746 5879 7802 5888
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7576 4622 7604 5306
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7668 4321 7696 5306
rect 7654 4312 7710 4321
rect 7654 4247 7710 4256
rect 7484 4168 7696 4196
rect 7562 4040 7618 4049
rect 7472 4004 7524 4010
rect 7562 3975 7618 3984
rect 7472 3946 7524 3952
rect 7484 3670 7512 3946
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7392 1902 7420 3062
rect 7484 2553 7512 3606
rect 7576 3058 7604 3975
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7470 2544 7526 2553
rect 7470 2479 7526 2488
rect 7576 2417 7604 2994
rect 7562 2408 7618 2417
rect 7562 2343 7618 2352
rect 7380 1896 7432 1902
rect 7380 1838 7432 1844
rect 7668 480 7696 4168
rect 7760 3942 7788 5714
rect 7852 5012 7880 6190
rect 7944 5166 7972 6310
rect 8128 6168 8156 6752
rect 8312 6644 8340 7414
rect 8680 7392 8708 7686
rect 8588 7364 8708 7392
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8404 7002 8432 7278
rect 8392 6996 8444 7002
rect 8588 6984 8616 7364
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8680 7177 8708 7210
rect 8666 7168 8722 7177
rect 8666 7103 8722 7112
rect 8588 6956 8715 6984
rect 8392 6938 8444 6944
rect 8687 6798 8715 6956
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8220 6616 8340 6644
rect 8220 6236 8248 6616
rect 8772 6610 8800 7686
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8680 6582 8800 6610
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8352 6480 8648 6500
rect 8392 6384 8444 6390
rect 8576 6384 8628 6390
rect 8392 6326 8444 6332
rect 8496 6344 8576 6372
rect 8220 6208 8340 6236
rect 8128 6140 8248 6168
rect 8220 5760 8248 6140
rect 8128 5732 8248 5760
rect 8128 5692 8156 5732
rect 8312 5692 8340 6208
rect 8036 5664 8156 5692
rect 8220 5664 8340 5692
rect 8036 5216 8064 5664
rect 8220 5624 8248 5664
rect 8128 5596 8248 5624
rect 8128 5284 8156 5596
rect 8404 5556 8432 6326
rect 8496 6118 8524 6344
rect 8576 6326 8628 6332
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8588 5953 8616 6054
rect 8574 5944 8630 5953
rect 8574 5879 8630 5888
rect 8680 5658 8708 6582
rect 8758 6488 8814 6497
rect 8758 6423 8814 6432
rect 8680 5630 8715 5658
rect 8220 5528 8432 5556
rect 8220 5352 8248 5528
rect 8687 5522 8715 5630
rect 8680 5494 8715 5522
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8352 5392 8648 5412
rect 8220 5324 8432 5352
rect 8128 5256 8248 5284
rect 8036 5188 8156 5216
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 7852 4984 7972 5012
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7852 4486 7880 4626
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7852 4282 7880 4422
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 7852 1358 7880 3538
rect 7944 3126 7972 4984
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 8036 3738 8064 4490
rect 8128 4010 8156 5188
rect 8220 4214 8248 5256
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8312 4690 8340 5034
rect 8404 4826 8432 5324
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8588 4826 8616 5102
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8680 4554 8708 5494
rect 8772 5030 8800 6423
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8772 4457 8800 4558
rect 8758 4448 8814 4457
rect 8352 4380 8648 4400
rect 8758 4383 8814 4392
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 8758 4312 8814 4321
rect 8680 4270 8758 4298
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8298 4176 8354 4185
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8116 3664 8168 3670
rect 8036 3612 8116 3618
rect 8036 3606 8168 3612
rect 8036 3590 8156 3606
rect 8036 3194 8064 3590
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8128 3233 8156 3470
rect 8114 3224 8170 3233
rect 8024 3188 8076 3194
rect 8114 3159 8170 3168
rect 8024 3130 8076 3136
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 8022 2680 8078 2689
rect 8022 2615 8078 2624
rect 7930 2272 7986 2281
rect 7930 2207 7986 2216
rect 7944 1698 7972 2207
rect 7932 1692 7984 1698
rect 7932 1634 7984 1640
rect 7840 1352 7892 1358
rect 7840 1294 7892 1300
rect 8036 480 8064 2615
rect 8220 2514 8248 4150
rect 8298 4111 8354 4120
rect 8574 4176 8630 4185
rect 8574 4111 8576 4120
rect 8312 3942 8340 4111
rect 8628 4111 8630 4120
rect 8576 4082 8628 4088
rect 8484 4072 8536 4078
rect 8482 4040 8484 4049
rect 8536 4040 8538 4049
rect 8482 3975 8538 3984
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8680 3652 8708 4270
rect 8758 4247 8814 4256
rect 8864 4128 8892 6666
rect 8588 3624 8708 3652
rect 8772 4100 8892 4128
rect 8588 3466 8616 3624
rect 8772 3584 8800 4100
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 8680 3556 8800 3584
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8352 3216 8648 3236
rect 8680 2990 8708 3556
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8576 2644 8628 2650
rect 8772 2632 8800 3402
rect 8628 2604 8800 2632
rect 8576 2586 8628 2592
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 8484 1896 8536 1902
rect 8484 1838 8536 1844
rect 8496 480 8524 1838
rect 8680 1426 8708 2604
rect 8864 2553 8892 3946
rect 8956 2990 8984 12650
rect 9220 12640 9272 12646
rect 9034 12608 9090 12617
rect 9220 12582 9272 12588
rect 9034 12543 9090 12552
rect 9048 9926 9076 12543
rect 9232 12374 9260 12582
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9220 12368 9272 12374
rect 9220 12310 9272 12316
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 10266 9168 12038
rect 9324 10266 9352 12378
rect 9416 11286 9444 14010
rect 9508 13530 9536 16050
rect 9600 15910 9628 16215
rect 9772 16186 9824 16192
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9692 16017 9720 16118
rect 9678 16008 9734 16017
rect 9678 15943 9734 15952
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9784 15706 9812 15846
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9600 14113 9628 15098
rect 9692 14346 9720 15370
rect 9876 15094 9904 17002
rect 9864 15088 9916 15094
rect 9864 15030 9916 15036
rect 9862 14784 9918 14793
rect 9862 14719 9918 14728
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9586 14104 9642 14113
rect 9586 14039 9642 14048
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9508 11082 9536 13466
rect 9600 13394 9628 13738
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9692 13258 9720 13806
rect 9784 13394 9812 14350
rect 9876 14278 9904 14719
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9968 14090 9996 17303
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 10060 16969 10088 17002
rect 10046 16960 10102 16969
rect 10046 16895 10102 16904
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 10060 15722 10088 16594
rect 10152 16590 10180 18142
rect 10336 17542 10364 19520
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10244 16969 10272 17138
rect 10230 16960 10286 16969
rect 10230 16895 10286 16904
rect 10336 16810 10364 17478
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10244 16782 10364 16810
rect 10140 16584 10192 16590
rect 10138 16552 10140 16561
rect 10192 16552 10194 16561
rect 10138 16487 10194 16496
rect 10138 16416 10194 16425
rect 10138 16351 10194 16360
rect 10152 15910 10180 16351
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10244 15722 10272 16782
rect 10428 16658 10456 16934
rect 10520 16726 10548 17070
rect 10612 16998 10640 18022
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10508 16720 10560 16726
rect 10508 16662 10560 16668
rect 10704 16674 10732 19520
rect 11072 18154 11100 19520
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 10796 17338 10824 17478
rect 11256 17338 11284 17478
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 10817 16892 11113 16912
rect 10873 16890 10897 16892
rect 10953 16890 10977 16892
rect 11033 16890 11057 16892
rect 10895 16838 10897 16890
rect 10959 16838 10971 16890
rect 11033 16838 11035 16890
rect 10873 16836 10897 16838
rect 10953 16836 10977 16838
rect 11033 16836 11057 16838
rect 10817 16816 11113 16836
rect 10416 16652 10468 16658
rect 10704 16646 10824 16674
rect 10416 16594 10468 16600
rect 10796 15892 10824 16646
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10980 16250 11008 16526
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10980 16114 11008 16186
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10520 15864 10824 15892
rect 10414 15736 10470 15745
rect 10060 15694 10180 15722
rect 10244 15694 10364 15722
rect 10152 15484 10180 15694
rect 10152 15456 10272 15484
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 10060 15094 10088 15370
rect 10138 15328 10194 15337
rect 10138 15263 10194 15272
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 10152 14822 10180 15263
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 10060 14113 10088 14282
rect 10152 14249 10180 14350
rect 10138 14240 10194 14249
rect 10138 14175 10194 14184
rect 9876 14062 9996 14090
rect 10046 14104 10102 14113
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9770 13016 9826 13025
rect 9588 12980 9640 12986
rect 9770 12951 9826 12960
rect 9588 12922 9640 12928
rect 9600 12782 9628 12922
rect 9784 12918 9812 12951
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9692 12209 9720 12718
rect 9772 12640 9824 12646
rect 9770 12608 9772 12617
rect 9824 12608 9826 12617
rect 9770 12543 9826 12552
rect 9770 12472 9826 12481
rect 9770 12407 9826 12416
rect 9784 12306 9812 12407
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9678 12200 9734 12209
rect 9678 12135 9734 12144
rect 9876 11914 9904 14062
rect 10046 14039 10102 14048
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9968 13870 9996 13942
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9968 12986 9996 13670
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9968 12073 9996 12582
rect 10060 12442 10088 13806
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 9954 12064 10010 12073
rect 9954 11999 10010 12008
rect 9876 11886 9996 11914
rect 9864 11824 9916 11830
rect 9862 11792 9864 11801
rect 9916 11792 9918 11801
rect 9862 11727 9918 11736
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9692 10674 9720 11086
rect 9770 10840 9826 10849
rect 9770 10775 9826 10784
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9034 9752 9090 9761
rect 9034 9687 9090 9696
rect 9048 9654 9076 9687
rect 9036 9648 9088 9654
rect 9036 9590 9088 9596
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9048 8974 9076 9454
rect 9126 9208 9182 9217
rect 9232 9178 9260 9862
rect 9126 9143 9182 9152
rect 9220 9172 9272 9178
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9048 8838 9076 8910
rect 9140 8838 9168 9143
rect 9220 9114 9272 9120
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9232 8514 9260 8842
rect 9140 8486 9260 8514
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 7750 9076 8230
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9140 7274 9168 8486
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9232 7585 9260 8366
rect 9218 7576 9274 7585
rect 9218 7511 9274 7520
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 9128 7268 9180 7274
rect 9128 7210 9180 7216
rect 9048 5574 9076 7210
rect 9324 6984 9352 9998
rect 9402 9888 9458 9897
rect 9402 9823 9458 9832
rect 9416 9450 9444 9823
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9416 7342 9444 8978
rect 9508 8906 9536 10202
rect 9692 10062 9720 10610
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9518 9720 9998
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9600 9178 9628 9454
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 9217 9720 9318
rect 9678 9208 9734 9217
rect 9588 9172 9640 9178
rect 9678 9143 9734 9152
rect 9588 9114 9640 9120
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9494 8800 9550 8809
rect 9494 8735 9550 8744
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9232 6956 9352 6984
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9140 6304 9168 6802
rect 9232 6497 9260 6956
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9218 6488 9274 6497
rect 9218 6423 9274 6432
rect 9140 6276 9260 6304
rect 9126 6216 9182 6225
rect 9126 6151 9182 6160
rect 9140 5681 9168 6151
rect 9232 6118 9260 6276
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9126 5672 9182 5681
rect 9126 5607 9182 5616
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9048 5098 9076 5510
rect 9232 5370 9260 5714
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9126 5264 9182 5273
rect 9126 5199 9182 5208
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 9140 4826 9168 5199
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 9048 4457 9076 4694
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9034 4448 9090 4457
rect 9034 4383 9090 4392
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9048 3738 9076 4082
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 9048 2650 9076 3402
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 8850 2544 8906 2553
rect 8850 2479 8906 2488
rect 8758 2136 8814 2145
rect 8758 2071 8814 2080
rect 8772 1902 8800 2071
rect 8760 1896 8812 1902
rect 8760 1838 8812 1844
rect 8956 1601 8984 2586
rect 9140 2446 9168 4218
rect 9232 3194 9260 4626
rect 9324 3738 9352 6666
rect 9416 6254 9444 6802
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9402 5944 9458 5953
rect 9402 5879 9458 5888
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9310 3632 9366 3641
rect 9310 3567 9366 3576
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9324 2689 9352 3567
rect 9416 3058 9444 5879
rect 9508 5234 9536 8735
rect 9692 8430 9720 8910
rect 9784 8498 9812 10775
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9680 8424 9732 8430
rect 9600 8384 9680 8412
rect 9600 7954 9628 8384
rect 9680 8366 9732 8372
rect 9678 8120 9734 8129
rect 9678 8055 9734 8064
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9586 7712 9642 7721
rect 9586 7647 9642 7656
rect 9600 7546 9628 7647
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9600 5778 9628 7210
rect 9692 6730 9720 8055
rect 9770 7712 9826 7721
rect 9770 7647 9826 7656
rect 9784 7041 9812 7647
rect 9770 7032 9826 7041
rect 9770 6967 9826 6976
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9508 4622 9536 5170
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9508 4185 9536 4558
rect 9494 4176 9550 4185
rect 9494 4111 9550 4120
rect 9600 4060 9628 5510
rect 9692 5370 9720 6054
rect 9784 5846 9812 6734
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9680 5364 9732 5370
rect 9732 5324 9812 5352
rect 9680 5306 9732 5312
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9692 4457 9720 4966
rect 9678 4448 9734 4457
rect 9678 4383 9734 4392
rect 9678 4312 9734 4321
rect 9678 4247 9734 4256
rect 9508 4032 9628 4060
rect 9508 3602 9536 4032
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9692 3534 9720 4247
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9310 2680 9366 2689
rect 9310 2615 9366 2624
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 8942 1592 8998 1601
rect 8942 1527 8998 1536
rect 8668 1420 8720 1426
rect 8668 1362 8720 1368
rect 9312 1352 9364 1358
rect 9416 1329 9444 2314
rect 9600 1698 9628 3062
rect 9784 3058 9812 5324
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9876 2904 9904 11562
rect 9968 11121 9996 11886
rect 9954 11112 10010 11121
rect 9954 11047 10010 11056
rect 10060 10554 10088 12242
rect 10152 10674 10180 13942
rect 10244 12306 10272 15456
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10336 11880 10364 15694
rect 10414 15671 10416 15680
rect 10468 15671 10470 15680
rect 10416 15642 10468 15648
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 15337 10456 15438
rect 10414 15328 10470 15337
rect 10414 15263 10470 15272
rect 10520 14634 10548 15864
rect 10817 15804 11113 15824
rect 10873 15802 10897 15804
rect 10953 15802 10977 15804
rect 11033 15802 11057 15804
rect 10895 15750 10897 15802
rect 10959 15750 10971 15802
rect 11033 15750 11035 15802
rect 10873 15748 10897 15750
rect 10953 15748 10977 15750
rect 11033 15748 11057 15750
rect 10817 15728 11113 15748
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10598 15464 10654 15473
rect 10598 15399 10654 15408
rect 10244 11852 10364 11880
rect 10428 14606 10548 14634
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10060 10526 10180 10554
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10060 9722 10088 10406
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10046 9616 10102 9625
rect 10046 9551 10048 9560
rect 10100 9551 10102 9560
rect 10048 9522 10100 9528
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9968 8838 9996 9318
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 10046 8800 10102 8809
rect 10046 8735 10102 8744
rect 10060 8566 10088 8735
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9968 7546 9996 8434
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9968 6644 9996 7346
rect 10060 6798 10088 7686
rect 10152 7290 10180 10526
rect 10244 8537 10272 11852
rect 10322 11792 10378 11801
rect 10322 11727 10378 11736
rect 10230 8528 10286 8537
rect 10230 8463 10286 8472
rect 10336 7954 10364 11727
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10152 7262 10364 7290
rect 10140 7200 10192 7206
rect 10232 7200 10284 7206
rect 10140 7142 10192 7148
rect 10230 7168 10232 7177
rect 10284 7168 10286 7177
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9968 6616 10088 6644
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9968 4758 9996 6190
rect 9956 4752 10008 4758
rect 9956 4694 10008 4700
rect 10060 4434 10088 6616
rect 10152 5234 10180 7142
rect 10230 7103 10286 7112
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 10244 6458 10272 6870
rect 10336 6780 10364 7262
rect 10428 7002 10456 14606
rect 10508 14544 10560 14550
rect 10508 14486 10560 14492
rect 10520 14074 10548 14486
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10520 13394 10548 13466
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10612 12866 10640 15399
rect 10704 15162 10732 15642
rect 10968 15632 11020 15638
rect 10968 15574 11020 15580
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10782 15328 10838 15337
rect 10782 15263 10838 15272
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10796 14804 10824 15263
rect 10888 14958 10916 15438
rect 10980 15434 11008 15574
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 11072 15473 11100 15506
rect 11058 15464 11114 15473
rect 10968 15428 11020 15434
rect 11058 15399 11114 15408
rect 10968 15370 11020 15376
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10704 14776 10824 14804
rect 10704 13870 10732 14776
rect 10817 14716 11113 14736
rect 10873 14714 10897 14716
rect 10953 14714 10977 14716
rect 11033 14714 11057 14716
rect 10895 14662 10897 14714
rect 10959 14662 10971 14714
rect 11033 14662 11035 14714
rect 10873 14660 10897 14662
rect 10953 14660 10977 14662
rect 11033 14660 11057 14662
rect 10817 14640 11113 14660
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11072 14385 11100 14418
rect 11058 14376 11114 14385
rect 11058 14311 11114 14320
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10704 13025 10732 13670
rect 10817 13628 11113 13648
rect 10873 13626 10897 13628
rect 10953 13626 10977 13628
rect 11033 13626 11057 13628
rect 10895 13574 10897 13626
rect 10959 13574 10971 13626
rect 11033 13574 11035 13626
rect 10873 13572 10897 13574
rect 10953 13572 10977 13574
rect 11033 13572 11057 13574
rect 10817 13552 11113 13572
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 10690 13016 10746 13025
rect 11072 12986 11100 13194
rect 10690 12951 10746 12960
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10520 12838 10640 12866
rect 10874 12880 10930 12889
rect 10520 11898 10548 12838
rect 10874 12815 10876 12824
rect 10928 12815 10930 12824
rect 10876 12786 10928 12792
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10612 12481 10640 12718
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10598 12472 10654 12481
rect 10704 12442 10732 12650
rect 10817 12540 11113 12560
rect 10873 12538 10897 12540
rect 10953 12538 10977 12540
rect 11033 12538 11057 12540
rect 10895 12486 10897 12538
rect 10959 12486 10971 12538
rect 11033 12486 11035 12538
rect 10873 12484 10897 12486
rect 10953 12484 10977 12486
rect 11033 12484 11057 12486
rect 10817 12464 11113 12484
rect 10598 12407 10654 12416
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10968 12368 11020 12374
rect 10796 12328 10968 12356
rect 10598 12200 10654 12209
rect 10598 12135 10654 12144
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10506 11792 10562 11801
rect 10506 11727 10562 11736
rect 10520 11529 10548 11727
rect 10506 11520 10562 11529
rect 10506 11455 10562 11464
rect 10506 11384 10562 11393
rect 10506 11319 10562 11328
rect 10520 11286 10548 11319
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10506 10432 10562 10441
rect 10506 10367 10562 10376
rect 10520 10266 10548 10367
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10336 6752 10456 6780
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10324 6384 10376 6390
rect 10324 6326 10376 6332
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10244 5953 10272 6190
rect 10230 5944 10286 5953
rect 10230 5879 10286 5888
rect 10336 5710 10364 6326
rect 10324 5704 10376 5710
rect 10230 5672 10286 5681
rect 10324 5646 10376 5652
rect 10230 5607 10286 5616
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10152 4865 10180 5170
rect 10138 4856 10194 4865
rect 10244 4826 10272 5607
rect 10322 5536 10378 5545
rect 10322 5471 10378 5480
rect 10138 4791 10194 4800
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 9948 4406 10088 4434
rect 9948 4196 9976 4406
rect 10048 4208 10100 4214
rect 9948 4168 9996 4196
rect 9968 4060 9996 4168
rect 10152 4196 10180 4558
rect 10100 4168 10180 4196
rect 10048 4150 10100 4156
rect 10336 4146 10364 5471
rect 10428 5273 10456 6752
rect 10520 5370 10548 10066
rect 10612 9761 10640 12135
rect 10796 11626 10824 12328
rect 10968 12310 11020 12316
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10888 11694 10916 11834
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10817 11452 11113 11472
rect 10873 11450 10897 11452
rect 10953 11450 10977 11452
rect 11033 11450 11057 11452
rect 10895 11398 10897 11450
rect 10959 11398 10971 11450
rect 11033 11398 11035 11450
rect 10873 11396 10897 11398
rect 10953 11396 10977 11398
rect 11033 11396 11057 11398
rect 10817 11376 11113 11396
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10704 9897 10732 11086
rect 10796 11082 10824 11222
rect 11164 11098 11192 16390
rect 11256 15910 11284 16594
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11244 15904 11296 15910
rect 11242 15872 11244 15881
rect 11296 15872 11298 15881
rect 11242 15807 11298 15816
rect 11348 13938 11376 16186
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 11440 15638 11468 15982
rect 11532 15745 11560 19520
rect 11702 17232 11758 17241
rect 11702 17167 11758 17176
rect 11610 16688 11666 16697
rect 11716 16658 11744 17167
rect 11610 16623 11612 16632
rect 11664 16623 11666 16632
rect 11704 16652 11756 16658
rect 11612 16594 11664 16600
rect 11704 16594 11756 16600
rect 11794 16552 11850 16561
rect 11612 16516 11664 16522
rect 11794 16487 11850 16496
rect 11612 16458 11664 16464
rect 11518 15736 11574 15745
rect 11518 15671 11574 15680
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11348 12209 11376 12242
rect 11334 12200 11390 12209
rect 11334 12135 11390 12144
rect 11440 11626 11468 15574
rect 11518 15192 11574 15201
rect 11518 15127 11574 15136
rect 11532 14822 11560 15127
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11624 14482 11652 16458
rect 11702 16144 11758 16153
rect 11702 16079 11758 16088
rect 11716 16046 11744 16079
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11808 15552 11836 16487
rect 11900 16454 11928 19520
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12072 17264 12124 17270
rect 12072 17206 12124 17212
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11900 15609 11928 16118
rect 11716 15524 11836 15552
rect 11886 15600 11942 15609
rect 11886 15535 11942 15544
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11518 14240 11574 14249
rect 11518 14175 11574 14184
rect 11532 13394 11560 14175
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11624 13841 11652 13874
rect 11610 13832 11666 13841
rect 11610 13767 11666 13776
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11532 12850 11560 13126
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11334 11520 11390 11529
rect 11532 11506 11560 12582
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11334 11455 11390 11464
rect 11440 11478 11560 11506
rect 11348 11354 11376 11455
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 10784 11076 10836 11082
rect 11164 11070 11376 11098
rect 10784 11018 10836 11024
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 10817 10364 11113 10384
rect 10873 10362 10897 10364
rect 10953 10362 10977 10364
rect 11033 10362 11057 10364
rect 10895 10310 10897 10362
rect 10959 10310 10971 10362
rect 11033 10310 11035 10362
rect 10873 10308 10897 10310
rect 10953 10308 10977 10310
rect 11033 10308 11057 10310
rect 10817 10288 11113 10308
rect 11164 9994 11192 10474
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 10690 9888 10746 9897
rect 10690 9823 10746 9832
rect 10598 9752 10654 9761
rect 10796 9738 10824 9930
rect 11256 9897 11284 10746
rect 11242 9888 11298 9897
rect 11242 9823 11298 9832
rect 10598 9687 10654 9696
rect 10704 9710 10824 9738
rect 11152 9716 11204 9722
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10612 9217 10640 9386
rect 10598 9208 10654 9217
rect 10598 9143 10654 9152
rect 10704 8809 10732 9710
rect 11152 9658 11204 9664
rect 10817 9276 11113 9296
rect 10873 9274 10897 9276
rect 10953 9274 10977 9276
rect 11033 9274 11057 9276
rect 10895 9222 10897 9274
rect 10959 9222 10971 9274
rect 11033 9222 11035 9274
rect 10873 9220 10897 9222
rect 10953 9220 10977 9222
rect 11033 9220 11057 9222
rect 10817 9200 11113 9220
rect 10690 8800 10746 8809
rect 10690 8735 10746 8744
rect 11164 8650 11192 9658
rect 11256 8838 11284 9823
rect 11348 8838 11376 11070
rect 11440 8974 11468 11478
rect 11518 11384 11574 11393
rect 11518 11319 11520 11328
rect 11572 11319 11574 11328
rect 11520 11290 11572 11296
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11532 10674 11560 11154
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11624 10606 11652 11698
rect 11716 11354 11744 15524
rect 11888 15496 11940 15502
rect 11808 15456 11888 15484
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11716 11121 11744 11290
rect 11808 11150 11836 15456
rect 11888 15438 11940 15444
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11900 14414 11928 14962
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11900 13705 11928 13806
rect 11886 13696 11942 13705
rect 11886 13631 11942 13640
rect 11900 12306 11928 13631
rect 11992 13569 12020 17138
rect 12084 15638 12112 17206
rect 12176 16454 12204 17614
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12360 15858 12388 19520
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12544 16794 12572 17750
rect 12636 17338 12664 17818
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12728 16289 12756 19520
rect 13096 18170 13124 19520
rect 12912 18142 13124 18170
rect 12808 17944 12860 17950
rect 12808 17886 12860 17892
rect 12820 16794 12848 17886
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12912 16674 12940 18142
rect 12992 18012 13044 18018
rect 12992 17954 13044 17960
rect 13004 17202 13032 17954
rect 13556 17678 13584 19520
rect 13726 17912 13782 17921
rect 13726 17847 13782 17856
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13282 17436 13578 17456
rect 13338 17434 13362 17436
rect 13418 17434 13442 17436
rect 13498 17434 13522 17436
rect 13360 17382 13362 17434
rect 13424 17382 13436 17434
rect 13498 17382 13500 17434
rect 13338 17380 13362 17382
rect 13418 17380 13442 17382
rect 13498 17380 13522 17382
rect 13082 17368 13138 17377
rect 13282 17360 13578 17380
rect 13082 17303 13138 17312
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12820 16646 12940 16674
rect 13096 16658 13124 17303
rect 13740 17202 13768 17847
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13084 16652 13136 16658
rect 12714 16280 12770 16289
rect 12714 16215 12770 16224
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12176 15830 12388 15858
rect 12072 15632 12124 15638
rect 12072 15574 12124 15580
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 12084 15201 12112 15302
rect 12070 15192 12126 15201
rect 12070 15127 12126 15136
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 11978 13560 12034 13569
rect 11978 13495 11980 13504
rect 12032 13495 12034 13504
rect 11980 13466 12032 13472
rect 11992 13435 12020 13466
rect 11978 13152 12034 13161
rect 11978 13087 12034 13096
rect 11992 12628 12020 13087
rect 12084 12782 12112 14894
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 11992 12600 12112 12628
rect 11978 12472 12034 12481
rect 11978 12407 12034 12416
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11992 11506 12020 12407
rect 11900 11478 12020 11506
rect 11796 11144 11848 11150
rect 11702 11112 11758 11121
rect 11796 11086 11848 11092
rect 11900 11098 11928 11478
rect 12084 11150 12112 12600
rect 12176 12481 12204 15830
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12268 14521 12296 15642
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 12360 14618 12388 15370
rect 12452 15337 12480 15506
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12438 15328 12494 15337
rect 12438 15263 12494 15272
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14793 12480 14894
rect 12438 14784 12494 14793
rect 12438 14719 12494 14728
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12254 14512 12310 14521
rect 12254 14447 12310 14456
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12360 13938 12388 14350
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12256 13796 12308 13802
rect 12256 13738 12308 13744
rect 12268 13530 12296 13738
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12360 13326 12388 13874
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12452 12782 12480 13670
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12162 12472 12218 12481
rect 12162 12407 12218 12416
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12072 11144 12124 11150
rect 11702 11047 11758 11056
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11520 10464 11572 10470
rect 11518 10432 11520 10441
rect 11572 10432 11574 10441
rect 11518 10367 11574 10376
rect 11610 10296 11666 10305
rect 11610 10231 11612 10240
rect 11664 10231 11666 10240
rect 11612 10202 11664 10208
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11532 9450 11560 10066
rect 11716 10062 11744 10746
rect 11808 10742 11836 11086
rect 11900 11070 12020 11098
rect 12072 11086 12124 11092
rect 11796 10736 11848 10742
rect 11848 10696 11928 10724
rect 11796 10678 11848 10684
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11610 9752 11666 9761
rect 11610 9687 11612 9696
rect 11664 9687 11666 9696
rect 11612 9658 11664 9664
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11520 9444 11572 9450
rect 11520 9386 11572 9392
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11164 8622 11284 8650
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10612 7206 10640 8298
rect 10704 7732 10732 8298
rect 10817 8188 11113 8208
rect 10873 8186 10897 8188
rect 10953 8186 10977 8188
rect 11033 8186 11057 8188
rect 10895 8134 10897 8186
rect 10959 8134 10971 8186
rect 11033 8134 11035 8186
rect 10873 8132 10897 8134
rect 10953 8132 10977 8134
rect 11033 8132 11057 8134
rect 10817 8112 11113 8132
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10784 7744 10836 7750
rect 10704 7704 10784 7732
rect 10784 7686 10836 7692
rect 10796 7410 10824 7686
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10784 7268 10836 7274
rect 10704 7228 10784 7256
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10612 6798 10640 6938
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10612 5386 10640 6734
rect 10704 5846 10732 7228
rect 10888 7256 10916 7890
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11150 7848 11206 7857
rect 10980 7478 11008 7822
rect 11150 7783 11206 7792
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 11058 7440 11114 7449
rect 11058 7375 11114 7384
rect 11072 7274 11100 7375
rect 10836 7228 10916 7256
rect 11060 7268 11112 7274
rect 10784 7210 10836 7216
rect 11060 7210 11112 7216
rect 10817 7100 11113 7120
rect 10873 7098 10897 7100
rect 10953 7098 10977 7100
rect 11033 7098 11057 7100
rect 10895 7046 10897 7098
rect 10959 7046 10971 7098
rect 11033 7046 11035 7098
rect 10873 7044 10897 7046
rect 10953 7044 10977 7046
rect 11033 7044 11057 7046
rect 10817 7024 11113 7044
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 11072 6497 11100 6870
rect 11058 6488 11114 6497
rect 11058 6423 11114 6432
rect 11060 6316 11112 6322
rect 11164 6304 11192 7783
rect 11112 6276 11192 6304
rect 11060 6258 11112 6264
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 11256 5794 11284 8622
rect 11348 7342 11376 8774
rect 11440 8362 11468 8910
rect 11532 8498 11560 9386
rect 11624 8566 11652 9454
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11426 7712 11482 7721
rect 11426 7647 11482 7656
rect 11440 7449 11468 7647
rect 11426 7440 11482 7449
rect 11426 7375 11482 7384
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11348 6089 11376 7142
rect 11334 6080 11390 6089
rect 11334 6015 11390 6024
rect 11334 5944 11390 5953
rect 11334 5879 11336 5888
rect 11388 5879 11390 5888
rect 11336 5850 11388 5856
rect 10704 5545 10732 5782
rect 11256 5766 11376 5794
rect 10966 5672 11022 5681
rect 10966 5607 11022 5616
rect 11242 5672 11298 5681
rect 11242 5607 11298 5616
rect 10690 5536 10746 5545
rect 10690 5471 10746 5480
rect 10508 5364 10560 5370
rect 10612 5358 10732 5386
rect 10508 5306 10560 5312
rect 10414 5264 10470 5273
rect 10414 5199 10470 5208
rect 10428 5166 10456 5199
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10414 4992 10470 5001
rect 10414 4927 10470 4936
rect 10428 4298 10456 4927
rect 10600 4752 10652 4758
rect 10600 4694 10652 4700
rect 10428 4270 10548 4298
rect 10414 4176 10470 4185
rect 10324 4140 10376 4146
rect 10414 4111 10416 4120
rect 10324 4082 10376 4088
rect 10468 4111 10470 4120
rect 10416 4082 10468 4088
rect 9968 4032 10088 4060
rect 9954 3768 10010 3777
rect 9954 3703 10010 3712
rect 9968 3602 9996 3703
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 10060 3194 10088 4032
rect 10138 3904 10194 3913
rect 10138 3839 10194 3848
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 9692 2876 9904 2904
rect 9936 2916 9988 2922
rect 9692 2038 9720 2876
rect 9988 2864 9996 2904
rect 9936 2858 9996 2864
rect 9968 2836 9996 2858
rect 10060 2836 10088 2926
rect 9968 2808 10088 2836
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 9968 2310 9996 2518
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 9680 2032 9732 2038
rect 9680 1974 9732 1980
rect 10152 1902 10180 3839
rect 10336 3670 10364 4082
rect 10520 4078 10548 4270
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10416 3936 10468 3942
rect 10468 3896 10548 3924
rect 10416 3878 10468 3884
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10140 1896 10192 1902
rect 10140 1838 10192 1844
rect 9588 1692 9640 1698
rect 9588 1634 9640 1640
rect 9312 1294 9364 1300
rect 9402 1320 9458 1329
rect 8852 1216 8904 1222
rect 8852 1158 8904 1164
rect 8864 480 8892 1158
rect 9324 480 9352 1294
rect 9402 1255 9458 1264
rect 10244 1222 10272 3606
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10336 3194 10364 3470
rect 10428 3398 10456 3674
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10520 3058 10548 3896
rect 10612 3602 10640 4694
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10704 3534 10732 5358
rect 10980 5098 11008 5607
rect 11256 5574 11284 5607
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10817 4848 11113 4868
rect 11242 4856 11298 4865
rect 11164 4814 11242 4842
rect 11164 4740 11192 4814
rect 11242 4791 11298 4800
rect 10888 4712 11192 4740
rect 11244 4752 11296 4758
rect 10888 4554 10916 4712
rect 11244 4694 11296 4700
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10876 4208 10928 4214
rect 10874 4176 10876 4185
rect 10928 4176 10930 4185
rect 10980 4146 11008 4490
rect 11058 4312 11114 4321
rect 11058 4247 11060 4256
rect 11112 4247 11114 4256
rect 11060 4218 11112 4224
rect 10874 4111 10930 4120
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11072 4010 11100 4082
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10796 3194 10824 3470
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10508 2848 10560 2854
rect 10414 2816 10470 2825
rect 10600 2848 10652 2854
rect 10508 2790 10560 2796
rect 10598 2816 10600 2825
rect 10652 2816 10654 2825
rect 10414 2751 10470 2760
rect 10322 2680 10378 2689
rect 10322 2615 10378 2624
rect 10336 2446 10364 2615
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10336 1766 10364 2382
rect 10428 1766 10456 2751
rect 10324 1760 10376 1766
rect 10324 1702 10376 1708
rect 10416 1760 10468 1766
rect 10416 1702 10468 1708
rect 10232 1216 10284 1222
rect 9678 1184 9734 1193
rect 10232 1158 10284 1164
rect 9678 1119 9734 1128
rect 9692 480 9720 1119
rect 10138 1048 10194 1057
rect 10138 983 10194 992
rect 10152 480 10180 983
rect 10520 480 10548 2790
rect 10598 2751 10654 2760
rect 10704 2446 10732 2994
rect 10980 2922 11008 3538
rect 11072 3058 11100 3606
rect 11164 3194 11192 4558
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10817 2672 11113 2692
rect 11164 2650 11192 2858
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 11072 2310 11100 2518
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11256 1834 11284 4694
rect 11348 4078 11376 5766
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11348 3194 11376 4014
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11440 2990 11468 7142
rect 11532 5710 11560 7822
rect 11624 7342 11652 8230
rect 11716 7698 11744 9998
rect 11808 8090 11836 10542
rect 11900 9722 11928 10696
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11992 9382 12020 11070
rect 12176 10266 12204 12310
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12164 9920 12216 9926
rect 12162 9888 12164 9897
rect 12216 9888 12218 9897
rect 12162 9823 12218 9832
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11900 9110 11928 9318
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11886 8664 11942 8673
rect 11886 8599 11888 8608
rect 11940 8599 11942 8608
rect 11888 8570 11940 8576
rect 12176 8294 12204 9658
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 11886 8120 11942 8129
rect 11796 8084 11848 8090
rect 11886 8055 11942 8064
rect 11796 8026 11848 8032
rect 11716 7670 11836 7698
rect 11702 7576 11758 7585
rect 11702 7511 11758 7520
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11532 5166 11560 5510
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4321 11560 4966
rect 11624 4672 11652 6802
rect 11716 6798 11744 7511
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11716 5778 11744 6258
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11704 5568 11756 5574
rect 11808 5545 11836 7670
rect 11704 5510 11756 5516
rect 11794 5536 11850 5545
rect 11716 5030 11744 5510
rect 11794 5471 11850 5480
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11900 4706 11928 8055
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11992 7857 12020 7890
rect 12072 7880 12124 7886
rect 11978 7848 12034 7857
rect 12072 7822 12124 7828
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 11978 7783 12034 7792
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11992 7410 12020 7482
rect 12084 7410 12112 7822
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11978 7304 12034 7313
rect 11978 7239 12034 7248
rect 12072 7268 12124 7274
rect 11992 7206 12020 7239
rect 12072 7210 12124 7216
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11992 5846 12020 6598
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11992 4978 12020 5646
rect 12084 5284 12112 7210
rect 12176 7002 12204 7822
rect 12268 7177 12296 12038
rect 12360 8430 12388 12718
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12452 11218 12480 11630
rect 12544 11354 12572 15438
rect 12728 14793 12756 16050
rect 12820 15910 12848 16646
rect 13084 16594 13136 16600
rect 13082 16144 13138 16153
rect 12992 16108 13044 16114
rect 13082 16079 13138 16088
rect 12992 16050 13044 16056
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15570 12848 15846
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12714 14784 12770 14793
rect 12714 14719 12770 14728
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12622 14104 12678 14113
rect 12622 14039 12678 14048
rect 12636 13546 12664 14039
rect 12728 14006 12756 14418
rect 12716 14000 12768 14006
rect 12912 13977 12940 15982
rect 12716 13942 12768 13948
rect 12898 13968 12954 13977
rect 12898 13903 12954 13912
rect 12636 13518 12848 13546
rect 12624 13456 12676 13462
rect 12676 13416 12756 13444
rect 12624 13398 12676 13404
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12636 12345 12664 12854
rect 12622 12336 12678 12345
rect 12622 12271 12678 12280
rect 12624 12232 12676 12238
rect 12622 12200 12624 12209
rect 12676 12200 12678 12209
rect 12622 12135 12678 12144
rect 12728 11898 12756 13416
rect 12820 12968 12848 13518
rect 13004 12986 13032 16050
rect 13096 15094 13124 16079
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 13084 14952 13136 14958
rect 13082 14920 13084 14929
rect 13136 14920 13138 14929
rect 13082 14855 13138 14864
rect 13188 14550 13216 17070
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13282 16348 13578 16368
rect 13338 16346 13362 16348
rect 13418 16346 13442 16348
rect 13498 16346 13522 16348
rect 13360 16294 13362 16346
rect 13424 16294 13436 16346
rect 13498 16294 13500 16346
rect 13338 16292 13362 16294
rect 13418 16292 13442 16294
rect 13498 16292 13522 16294
rect 13282 16272 13578 16292
rect 13450 16008 13506 16017
rect 13450 15943 13506 15952
rect 13464 15706 13492 15943
rect 13648 15910 13676 17002
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13282 15260 13578 15280
rect 13338 15258 13362 15260
rect 13418 15258 13442 15260
rect 13498 15258 13522 15260
rect 13360 15206 13362 15258
rect 13424 15206 13436 15258
rect 13498 15206 13500 15258
rect 13338 15204 13362 15206
rect 13418 15204 13442 15206
rect 13498 15204 13522 15206
rect 13282 15184 13578 15204
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 13176 14544 13228 14550
rect 13176 14486 13228 14492
rect 13542 14512 13598 14521
rect 13096 12986 13124 14486
rect 13542 14447 13544 14456
rect 13596 14447 13598 14456
rect 13544 14418 13596 14424
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 12992 12980 13044 12986
rect 12820 12940 12940 12968
rect 12806 12472 12862 12481
rect 12806 12407 12862 12416
rect 12820 12306 12848 12407
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12912 12238 12940 12940
rect 12992 12922 13044 12928
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12820 11937 12848 12106
rect 12806 11928 12862 11937
rect 12716 11892 12768 11898
rect 12806 11863 12862 11872
rect 12716 11834 12768 11840
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10266 12480 10406
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12452 9994 12480 10066
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 12636 9518 12664 11562
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12440 9444 12492 9450
rect 12440 9386 12492 9392
rect 12452 8634 12480 9386
rect 12728 8974 12756 11562
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12348 8424 12400 8430
rect 12400 8384 12480 8412
rect 12348 8366 12400 8372
rect 12348 8288 12400 8294
rect 12348 8230 12400 8236
rect 12254 7168 12310 7177
rect 12254 7103 12310 7112
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12162 6896 12218 6905
rect 12162 6831 12164 6840
rect 12216 6831 12218 6840
rect 12164 6802 12216 6808
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12176 5710 12204 6326
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12268 5302 12296 6666
rect 12360 6322 12388 8230
rect 12452 7993 12480 8384
rect 12438 7984 12494 7993
rect 12438 7919 12494 7928
rect 12544 7834 12572 8910
rect 12716 8560 12768 8566
rect 12622 8528 12678 8537
rect 12716 8502 12768 8508
rect 12622 8463 12678 8472
rect 12452 7806 12572 7834
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12360 5778 12388 6258
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12346 5672 12402 5681
rect 12346 5607 12348 5616
rect 12400 5607 12402 5616
rect 12348 5578 12400 5584
rect 12452 5370 12480 7806
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12544 5545 12572 7686
rect 12636 7002 12664 8463
rect 12728 7041 12756 8502
rect 12714 7032 12770 7041
rect 12624 6996 12676 7002
rect 12714 6967 12770 6976
rect 12624 6938 12676 6944
rect 12716 6928 12768 6934
rect 12622 6896 12678 6905
rect 12716 6870 12768 6876
rect 12622 6831 12678 6840
rect 12636 6798 12664 6831
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12728 6633 12756 6870
rect 12820 6662 12848 11290
rect 12912 10810 12940 12174
rect 13004 11937 13032 12922
rect 13188 12832 13216 14214
rect 13282 14172 13578 14192
rect 13338 14170 13362 14172
rect 13418 14170 13442 14172
rect 13498 14170 13522 14172
rect 13360 14118 13362 14170
rect 13424 14118 13436 14170
rect 13498 14118 13500 14170
rect 13338 14116 13362 14118
rect 13418 14116 13442 14118
rect 13498 14116 13522 14118
rect 13282 14096 13578 14116
rect 13360 14000 13412 14006
rect 13360 13942 13412 13948
rect 13268 13864 13320 13870
rect 13266 13832 13268 13841
rect 13320 13832 13322 13841
rect 13266 13767 13322 13776
rect 13266 13696 13322 13705
rect 13266 13631 13322 13640
rect 13280 13394 13308 13631
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13372 13297 13400 13942
rect 13648 13870 13676 15846
rect 13820 15088 13872 15094
rect 13818 15056 13820 15065
rect 13872 15056 13874 15065
rect 13818 14991 13874 15000
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13832 14074 13860 14350
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13726 13968 13782 13977
rect 13726 13903 13782 13912
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13358 13288 13414 13297
rect 13358 13223 13414 13232
rect 13648 13172 13676 13806
rect 13740 13326 13768 13903
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 13462 13860 13670
rect 13924 13530 13952 19520
rect 14384 17796 14412 19520
rect 14384 17768 14596 17796
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14186 17096 14242 17105
rect 14186 17031 14242 17040
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 13912 13524 13964 13530
rect 14016 13512 14044 16526
rect 14200 15706 14228 17031
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14108 15042 14136 15506
rect 14108 15014 14228 15042
rect 14016 13484 14136 13512
rect 13912 13466 13964 13472
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 14002 13424 14058 13433
rect 14002 13359 14058 13368
rect 14016 13326 14044 13359
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13820 13252 13872 13258
rect 13820 13194 13872 13200
rect 13648 13144 13768 13172
rect 13282 13084 13578 13104
rect 13338 13082 13362 13084
rect 13418 13082 13442 13084
rect 13498 13082 13522 13084
rect 13360 13030 13362 13082
rect 13424 13030 13436 13082
rect 13498 13030 13500 13082
rect 13338 13028 13362 13030
rect 13418 13028 13442 13030
rect 13498 13028 13522 13030
rect 13282 13008 13578 13028
rect 13188 12804 13308 12832
rect 13174 12744 13230 12753
rect 13174 12679 13230 12688
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 12990 11928 13046 11937
rect 12990 11863 13046 11872
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 13004 11354 13032 11562
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13096 11218 13124 12582
rect 13188 11286 13216 12679
rect 13280 12374 13308 12804
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 13282 11996 13578 12016
rect 13338 11994 13362 11996
rect 13418 11994 13442 11996
rect 13498 11994 13522 11996
rect 13360 11942 13362 11994
rect 13424 11942 13436 11994
rect 13498 11942 13500 11994
rect 13338 11940 13362 11942
rect 13418 11940 13442 11942
rect 13498 11940 13522 11942
rect 13282 11920 13578 11940
rect 13648 11880 13676 12650
rect 13556 11852 13676 11880
rect 13452 11552 13504 11558
rect 13556 11540 13584 11852
rect 13504 11512 13584 11540
rect 13636 11552 13688 11558
rect 13452 11494 13504 11500
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 13556 11218 13584 11512
rect 13634 11520 13636 11529
rect 13688 11520 13690 11529
rect 13634 11455 13690 11464
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12912 7954 12940 10406
rect 13004 9586 13032 10610
rect 13096 10470 13124 11154
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13280 10996 13308 11086
rect 13188 10968 13308 10996
rect 13188 10792 13216 10968
rect 13282 10908 13578 10928
rect 13338 10906 13362 10908
rect 13418 10906 13442 10908
rect 13498 10906 13522 10908
rect 13360 10854 13362 10906
rect 13424 10854 13436 10906
rect 13498 10854 13500 10906
rect 13338 10852 13362 10854
rect 13418 10852 13442 10854
rect 13498 10852 13522 10854
rect 13282 10832 13578 10852
rect 13636 10804 13688 10810
rect 13188 10764 13308 10792
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13096 9722 13124 10066
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12912 6866 12940 7890
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 13004 6730 13032 9318
rect 13188 9110 13216 10610
rect 13280 10538 13308 10764
rect 13636 10746 13688 10752
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13464 10010 13492 10678
rect 13648 10130 13676 10746
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13464 9982 13676 10010
rect 13282 9820 13578 9840
rect 13338 9818 13362 9820
rect 13418 9818 13442 9820
rect 13498 9818 13522 9820
rect 13360 9766 13362 9818
rect 13424 9766 13436 9818
rect 13498 9766 13500 9818
rect 13338 9764 13362 9766
rect 13418 9764 13442 9766
rect 13498 9764 13522 9766
rect 13282 9744 13578 9764
rect 13648 9654 13676 9982
rect 13740 9897 13768 13144
rect 13832 12850 13860 13194
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13818 11656 13874 11665
rect 14108 11642 14136 13484
rect 13818 11591 13874 11600
rect 14016 11614 14136 11642
rect 13832 10266 13860 11591
rect 13910 11112 13966 11121
rect 14016 11082 14044 11614
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 11354 14136 11494
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 13910 11047 13966 11056
rect 14004 11076 14056 11082
rect 13924 10962 13952 11047
rect 14004 11018 14056 11024
rect 13924 10934 14044 10962
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13924 10538 13952 10746
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13818 10160 13874 10169
rect 13818 10095 13820 10104
rect 13872 10095 13874 10104
rect 13820 10066 13872 10072
rect 13924 10010 13952 10474
rect 13832 9982 13952 10010
rect 13726 9888 13782 9897
rect 13726 9823 13782 9832
rect 13832 9738 13860 9982
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13740 9710 13860 9738
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13634 9480 13690 9489
rect 13280 9217 13308 9454
rect 13634 9415 13690 9424
rect 13648 9382 13676 9415
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13266 9208 13322 9217
rect 13266 9143 13322 9152
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13634 9072 13690 9081
rect 13634 9007 13690 9016
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13358 8936 13414 8945
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13096 8430 13124 8842
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 12808 6656 12860 6662
rect 12714 6624 12770 6633
rect 12808 6598 12860 6604
rect 12714 6559 12770 6568
rect 13096 6440 13124 7414
rect 12912 6412 13124 6440
rect 12806 6352 12862 6361
rect 12806 6287 12862 6296
rect 12820 6254 12848 6287
rect 12624 6248 12676 6254
rect 12808 6248 12860 6254
rect 12676 6208 12756 6236
rect 12624 6190 12676 6196
rect 12624 6112 12676 6118
rect 12728 6100 12756 6208
rect 12808 6190 12860 6196
rect 12728 6072 12848 6100
rect 12624 6054 12676 6060
rect 12636 5914 12664 6054
rect 12714 5944 12770 5953
rect 12624 5908 12676 5914
rect 12714 5879 12770 5888
rect 12624 5850 12676 5856
rect 12728 5760 12756 5879
rect 12636 5732 12756 5760
rect 12530 5536 12586 5545
rect 12530 5471 12586 5480
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12164 5296 12216 5302
rect 12084 5256 12164 5284
rect 12164 5238 12216 5244
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 11992 4950 12112 4978
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11992 4729 12020 4762
rect 11704 4684 11756 4690
rect 11624 4644 11704 4672
rect 11518 4312 11574 4321
rect 11518 4247 11574 4256
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11532 4010 11560 4150
rect 11520 4004 11572 4010
rect 11520 3946 11572 3952
rect 11624 3670 11652 4644
rect 11704 4626 11756 4632
rect 11808 4678 11928 4706
rect 11978 4720 12034 4729
rect 11702 4312 11758 4321
rect 11702 4247 11758 4256
rect 11716 3913 11744 4247
rect 11702 3904 11758 3913
rect 11702 3839 11758 3848
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11808 3584 11836 4678
rect 11978 4655 12034 4664
rect 12084 4622 12112 4950
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11900 4282 11928 4490
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11992 4026 12020 4218
rect 12176 4146 12204 5238
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12268 4826 12296 5102
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12348 4752 12400 4758
rect 12346 4720 12348 4729
rect 12400 4720 12402 4729
rect 12346 4655 12402 4664
rect 12440 4616 12492 4622
rect 12438 4584 12440 4593
rect 12492 4584 12494 4593
rect 12438 4519 12494 4528
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12268 4214 12296 4422
rect 12256 4208 12308 4214
rect 12544 4185 12572 5306
rect 12636 5234 12664 5732
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12636 4622 12664 4762
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12622 4312 12678 4321
rect 12622 4247 12678 4256
rect 12256 4150 12308 4156
rect 12530 4176 12586 4185
rect 12164 4140 12216 4146
rect 12636 4146 12664 4247
rect 12530 4111 12586 4120
rect 12624 4140 12676 4146
rect 12164 4082 12216 4088
rect 12624 4082 12676 4088
rect 12532 4072 12584 4078
rect 11900 4010 12020 4026
rect 11888 4004 12020 4010
rect 11940 3998 12020 4004
rect 12070 4040 12126 4049
rect 12532 4014 12584 4020
rect 12070 3975 12126 3984
rect 11888 3946 11940 3952
rect 11716 3556 11836 3584
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11624 3398 11652 3470
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11428 2848 11480 2854
rect 11624 2825 11652 2926
rect 11428 2790 11480 2796
rect 11610 2816 11666 2825
rect 11440 2514 11468 2790
rect 11610 2751 11666 2760
rect 11518 2544 11574 2553
rect 11428 2508 11480 2514
rect 11518 2479 11574 2488
rect 11428 2450 11480 2456
rect 11334 2272 11390 2281
rect 11334 2207 11390 2216
rect 11244 1828 11296 1834
rect 11244 1770 11296 1776
rect 10968 1284 11020 1290
rect 10968 1226 11020 1232
rect 10980 480 11008 1226
rect 11348 480 11376 2207
rect 11532 1873 11560 2479
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11624 2106 11652 2382
rect 11716 2310 11744 3556
rect 11900 3482 11928 3946
rect 12084 3942 12112 3975
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12544 3670 12572 4014
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11808 3454 11928 3482
rect 11808 2922 11836 3454
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 11794 2816 11850 2825
rect 11794 2751 11850 2760
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11612 2100 11664 2106
rect 11612 2042 11664 2048
rect 11518 1864 11574 1873
rect 11518 1799 11574 1808
rect 11808 480 11836 2751
rect 11900 1630 11928 3334
rect 11992 3233 12020 3538
rect 12162 3496 12218 3505
rect 12162 3431 12218 3440
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 11978 3224 12034 3233
rect 11978 3159 12034 3168
rect 11992 2938 12020 3159
rect 12084 3058 12112 3334
rect 12176 3097 12204 3431
rect 12162 3088 12218 3097
rect 12072 3052 12124 3058
rect 12162 3023 12218 3032
rect 12072 2994 12124 3000
rect 11992 2910 12112 2938
rect 12084 2514 12112 2910
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 12176 2689 12204 2858
rect 12162 2680 12218 2689
rect 12162 2615 12218 2624
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 11992 1970 12020 2450
rect 12164 2100 12216 2106
rect 12164 2042 12216 2048
rect 11980 1964 12032 1970
rect 11980 1906 12032 1912
rect 11888 1624 11940 1630
rect 11888 1566 11940 1572
rect 12176 480 12204 2042
rect 12360 1970 12388 3606
rect 12636 3534 12664 4082
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12452 3058 12480 3470
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 2650 12480 2790
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12544 2417 12572 2994
rect 12636 2990 12664 3470
rect 12728 3194 12756 5578
rect 12820 5545 12848 6072
rect 12806 5536 12862 5545
rect 12806 5471 12862 5480
rect 12912 4826 12940 6412
rect 12990 6352 13046 6361
rect 12990 6287 13046 6296
rect 13084 6316 13136 6322
rect 13004 5778 13032 6287
rect 13084 6258 13136 6264
rect 13096 6186 13124 6258
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 12992 5568 13044 5574
rect 12990 5536 12992 5545
rect 13044 5536 13046 5545
rect 12990 5471 13046 5480
rect 13096 5166 13124 5578
rect 13188 5352 13216 8910
rect 13358 8871 13360 8880
rect 13412 8871 13414 8880
rect 13360 8842 13412 8848
rect 13282 8732 13578 8752
rect 13338 8730 13362 8732
rect 13418 8730 13442 8732
rect 13498 8730 13522 8732
rect 13360 8678 13362 8730
rect 13424 8678 13436 8730
rect 13498 8678 13500 8730
rect 13338 8676 13362 8678
rect 13418 8676 13442 8678
rect 13498 8676 13522 8678
rect 13282 8656 13578 8676
rect 13648 8634 13676 9007
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13740 7954 13768 9710
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13832 8498 13860 8910
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13282 7644 13578 7664
rect 13338 7642 13362 7644
rect 13418 7642 13442 7644
rect 13498 7642 13522 7644
rect 13360 7590 13362 7642
rect 13424 7590 13436 7642
rect 13498 7590 13500 7642
rect 13338 7588 13362 7590
rect 13418 7588 13442 7590
rect 13498 7588 13522 7590
rect 13282 7568 13578 7588
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13648 6458 13676 6802
rect 13728 6792 13780 6798
rect 13726 6760 13728 6769
rect 13780 6760 13782 6769
rect 13726 6695 13782 6704
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13280 5710 13308 6326
rect 13544 6112 13596 6118
rect 13728 6112 13780 6118
rect 13544 6054 13596 6060
rect 13634 6080 13690 6089
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13556 5642 13584 6054
rect 13728 6054 13780 6060
rect 13634 6015 13690 6024
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13648 5352 13676 6015
rect 13188 5324 13308 5352
rect 13174 5264 13230 5273
rect 13174 5199 13230 5208
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12806 4720 12862 4729
rect 12862 4678 13124 4706
rect 12806 4655 12862 4664
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12820 4026 12848 4150
rect 12912 4146 12940 4558
rect 12990 4176 13046 4185
rect 12900 4140 12952 4146
rect 12990 4111 13046 4120
rect 12900 4082 12952 4088
rect 12820 3998 12940 4026
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12820 3738 12848 3878
rect 12912 3754 12940 3998
rect 13004 3942 13032 4111
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 12808 3732 12860 3738
rect 12912 3726 13032 3754
rect 13096 3738 13124 4678
rect 12808 3674 12860 3680
rect 12900 3664 12952 3670
rect 12898 3632 12900 3641
rect 12952 3632 12954 3641
rect 13004 3618 13032 3726
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13004 3590 13124 3618
rect 12898 3567 12954 3576
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12806 3360 12862 3369
rect 12806 3295 12862 3304
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12622 2680 12678 2689
rect 12622 2615 12624 2624
rect 12676 2615 12678 2624
rect 12624 2586 12676 2592
rect 12530 2408 12586 2417
rect 12530 2343 12586 2352
rect 12820 2281 12848 3295
rect 13004 3058 13032 3470
rect 13096 3369 13124 3590
rect 13082 3360 13138 3369
rect 13082 3295 13138 3304
rect 13082 3224 13138 3233
rect 13082 3159 13138 3168
rect 13096 3058 13124 3159
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 13096 2650 13124 2994
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 12806 2272 12862 2281
rect 12806 2207 12862 2216
rect 12348 1964 12400 1970
rect 12348 1906 12400 1912
rect 12624 1420 12676 1426
rect 12624 1362 12676 1368
rect 12636 480 12664 1362
rect 12912 1193 12940 2382
rect 13188 2258 13216 5199
rect 13280 5001 13308 5324
rect 13556 5324 13676 5352
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13266 4992 13322 5001
rect 13266 4927 13322 4936
rect 13372 4865 13400 5170
rect 13450 4992 13506 5001
rect 13450 4927 13506 4936
rect 13358 4856 13414 4865
rect 13358 4791 13414 4800
rect 13464 4758 13492 4927
rect 13556 4842 13584 5324
rect 13634 5128 13690 5137
rect 13634 5063 13690 5072
rect 13648 5030 13676 5063
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13556 4814 13676 4842
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13282 4380 13578 4400
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13266 4040 13322 4049
rect 13266 3975 13322 3984
rect 13280 3942 13308 3975
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13556 3534 13584 4082
rect 13648 4010 13676 4814
rect 13740 4729 13768 6054
rect 13832 5370 13860 8298
rect 13924 7274 13952 9862
rect 14016 9518 14044 10934
rect 14108 10810 14136 11154
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 9178 14044 9318
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 14016 8090 14044 8230
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 13910 7032 13966 7041
rect 13910 6967 13966 6976
rect 13924 6798 13952 6967
rect 14016 6905 14044 7142
rect 14002 6896 14058 6905
rect 14108 6866 14136 10542
rect 14200 9625 14228 15014
rect 14292 12306 14320 16390
rect 14476 14890 14504 17614
rect 14568 16454 14596 17768
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14476 13988 14504 14826
rect 14384 13960 14504 13988
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14278 11248 14334 11257
rect 14278 11183 14280 11192
rect 14332 11183 14334 11192
rect 14280 11154 14332 11160
rect 14384 10606 14412 13960
rect 14462 12472 14518 12481
rect 14462 12407 14518 12416
rect 14476 11778 14504 12407
rect 14660 11937 14688 15982
rect 14646 11928 14702 11937
rect 14646 11863 14702 11872
rect 14476 11750 14596 11778
rect 14752 11762 14780 19520
rect 15120 16561 15148 19520
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15106 16552 15162 16561
rect 15106 16487 15162 16496
rect 15212 15314 15240 17546
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15120 15286 15240 15314
rect 14924 14544 14976 14550
rect 14924 14486 14976 14492
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14476 10146 14504 11630
rect 14568 10606 14596 11750
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14740 11620 14792 11626
rect 14740 11562 14792 11568
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14292 10118 14504 10146
rect 14186 9616 14242 9625
rect 14186 9551 14242 9560
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14200 7818 14228 8774
rect 14292 7886 14320 10118
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14188 7812 14240 7818
rect 14188 7754 14240 7760
rect 14200 7410 14228 7754
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14002 6831 14058 6840
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 13912 6792 13964 6798
rect 14200 6746 14228 6938
rect 13912 6734 13964 6740
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 14108 6718 14228 6746
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13818 5264 13874 5273
rect 13924 5234 13952 6122
rect 14016 5302 14044 6666
rect 14108 5370 14136 6718
rect 14292 6390 14320 7822
rect 14384 7546 14412 9998
rect 14476 8498 14504 9998
rect 14568 9217 14596 10542
rect 14554 9208 14610 9217
rect 14554 9143 14610 9152
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14370 7440 14426 7449
rect 14370 7375 14426 7384
rect 14384 7206 14412 7375
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 14186 5944 14242 5953
rect 14186 5879 14242 5888
rect 14370 5944 14426 5953
rect 14370 5879 14426 5888
rect 14200 5778 14228 5879
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14278 5672 14334 5681
rect 14278 5607 14334 5616
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 13818 5199 13874 5208
rect 13912 5228 13964 5234
rect 13832 5166 13860 5199
rect 13912 5170 13964 5176
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13726 4720 13782 4729
rect 13726 4655 13782 4664
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13634 3768 13690 3777
rect 13634 3703 13636 3712
rect 13688 3703 13690 3712
rect 13636 3674 13688 3680
rect 13544 3528 13596 3534
rect 13740 3482 13768 4150
rect 13544 3470 13596 3476
rect 13648 3454 13768 3482
rect 13832 3466 13860 4966
rect 13820 3460 13872 3466
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13280 2446 13308 2586
rect 13648 2582 13676 3454
rect 13820 3402 13872 3408
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 2961 13768 3334
rect 13818 3224 13874 3233
rect 13818 3159 13874 3168
rect 13726 2952 13782 2961
rect 13832 2922 13860 3159
rect 13924 3058 13952 5034
rect 14016 4264 14044 5238
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14108 4690 14136 5170
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 14016 4236 14136 4264
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14108 2938 14136 4236
rect 14200 3097 14228 4966
rect 14292 3602 14320 5607
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 14186 3088 14242 3097
rect 14186 3023 14242 3032
rect 13726 2887 13782 2896
rect 13820 2916 13872 2922
rect 14016 2910 14136 2938
rect 13872 2876 13952 2904
rect 13820 2858 13872 2864
rect 13726 2816 13782 2825
rect 13726 2751 13782 2760
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13004 2230 13216 2258
rect 12898 1184 12954 1193
rect 12898 1119 12954 1128
rect 13004 480 13032 2230
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 13740 1986 13768 2751
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13832 2553 13860 2586
rect 13818 2544 13874 2553
rect 13818 2479 13874 2488
rect 13818 2272 13874 2281
rect 13818 2207 13874 2216
rect 13464 1958 13768 1986
rect 13464 480 13492 1958
rect 13832 480 13860 2207
rect 13924 2106 13952 2876
rect 14016 2854 14044 2910
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 14002 2680 14058 2689
rect 14002 2615 14058 2624
rect 14016 2514 14044 2615
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 13912 2100 13964 2106
rect 13912 2042 13964 2048
rect 14108 2009 14136 2790
rect 14292 2666 14320 3402
rect 14384 3058 14412 5879
rect 14476 4690 14504 8230
rect 14568 5914 14596 8910
rect 14660 6118 14688 11086
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14660 5817 14688 5850
rect 14646 5808 14702 5817
rect 14646 5743 14702 5752
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14568 3505 14596 5306
rect 14554 3496 14610 3505
rect 14554 3431 14610 3440
rect 14568 3058 14596 3431
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14556 2916 14608 2922
rect 14608 2876 14688 2904
rect 14556 2858 14608 2864
rect 14200 2638 14320 2666
rect 14094 2000 14150 2009
rect 14094 1935 14150 1944
rect 14200 1902 14228 2638
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14188 1896 14240 1902
rect 14188 1838 14240 1844
rect 14292 1737 14320 2450
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 14476 2038 14504 2382
rect 14464 2032 14516 2038
rect 14464 1974 14516 1980
rect 14278 1728 14334 1737
rect 14278 1663 14334 1672
rect 14278 1592 14334 1601
rect 14278 1527 14334 1536
rect 14292 480 14320 1527
rect 14660 480 14688 2876
rect 14752 2378 14780 11562
rect 14844 7342 14872 13466
rect 14936 10742 14964 14486
rect 15120 12481 15148 15286
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15106 12472 15162 12481
rect 15212 12442 15240 14894
rect 15106 12407 15162 12416
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 15028 10577 15056 11494
rect 15014 10568 15070 10577
rect 15014 10503 15070 10512
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15028 10033 15056 10406
rect 15014 10024 15070 10033
rect 15014 9959 15070 9968
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14844 2650 14872 6054
rect 14936 5846 14964 9454
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15016 8560 15068 8566
rect 15016 8502 15068 8508
rect 15028 8401 15056 8502
rect 15014 8392 15070 8401
rect 15014 8327 15070 8336
rect 15120 8265 15148 9114
rect 15106 8256 15162 8265
rect 15106 8191 15162 8200
rect 15014 6216 15070 6225
rect 15014 6151 15070 6160
rect 15028 6118 15056 6151
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 14924 5840 14976 5846
rect 14924 5782 14976 5788
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 14832 2508 14884 2514
rect 14832 2450 14884 2456
rect 14740 2372 14792 2378
rect 14740 2314 14792 2320
rect 14844 1494 14872 2450
rect 14936 1766 14964 4422
rect 15016 3936 15068 3942
rect 15014 3904 15016 3913
rect 15068 3904 15070 3913
rect 15014 3839 15070 3848
rect 15120 3754 15148 8191
rect 15028 3726 15148 3754
rect 15028 2825 15056 3726
rect 15212 2922 15240 12378
rect 15304 6254 15332 15438
rect 15580 13938 15608 19520
rect 15948 17610 15976 19520
rect 15936 17604 15988 17610
rect 15936 17546 15988 17552
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 16408 13802 16436 19520
rect 16776 16114 16804 19520
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15488 10713 15516 11698
rect 16408 11694 16436 13738
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 15474 10704 15530 10713
rect 15474 10639 15530 10648
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15304 4282 15332 6190
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 15108 2848 15160 2854
rect 15014 2816 15070 2825
rect 15108 2790 15160 2796
rect 15014 2751 15070 2760
rect 15120 2582 15148 2790
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 15396 1970 15424 9590
rect 15488 8430 15516 10639
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15488 4010 15516 8366
rect 15566 7304 15622 7313
rect 15566 7239 15622 7248
rect 15476 4004 15528 4010
rect 15476 3946 15528 3952
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15384 1964 15436 1970
rect 15384 1906 15436 1912
rect 14924 1760 14976 1766
rect 14924 1702 14976 1708
rect 14832 1488 14884 1494
rect 14832 1430 14884 1436
rect 15106 1456 15162 1465
rect 15106 1391 15162 1400
rect 15120 480 15148 1391
rect 15488 480 15516 2246
rect 15580 2009 15608 7239
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 15566 2000 15622 2009
rect 15566 1935 15622 1944
rect 15936 1964 15988 1970
rect 15936 1906 15988 1912
rect 15948 480 15976 1906
rect 16316 480 16344 3062
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16776 480 16804 2790
rect 1122 439 1178 448
rect 1398 0 1454 480
rect 1858 0 1914 480
rect 2226 0 2282 480
rect 2686 0 2742 480
rect 3054 0 3110 480
rect 3514 0 3570 480
rect 3882 0 3938 480
rect 4342 0 4398 480
rect 4710 0 4766 480
rect 5170 0 5226 480
rect 5538 0 5594 480
rect 5998 0 6054 480
rect 6366 0 6422 480
rect 6826 0 6882 480
rect 7194 0 7250 480
rect 7654 0 7710 480
rect 8022 0 8078 480
rect 8482 0 8538 480
rect 8850 0 8906 480
rect 9310 0 9366 480
rect 9678 0 9734 480
rect 10138 0 10194 480
rect 10506 0 10562 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12622 0 12678 480
rect 12990 0 13046 480
rect 13450 0 13506 480
rect 13818 0 13874 480
rect 14278 0 14334 480
rect 14646 0 14702 480
rect 15106 0 15162 480
rect 15474 0 15530 480
rect 15934 0 15990 480
rect 16302 0 16358 480
rect 16762 0 16818 480
<< via2 >>
rect 938 15952 994 16008
rect 2134 16632 2190 16688
rect 1858 15680 1914 15736
rect 1490 12552 1546 12608
rect 1214 9832 1270 9888
rect 938 7928 994 7984
rect 754 7112 810 7168
rect 846 5208 902 5264
rect 1858 11872 1914 11928
rect 1766 11192 1822 11248
rect 1766 11056 1822 11112
rect 1398 7928 1454 7984
rect 1398 5752 1454 5808
rect 1398 5072 1454 5128
rect 2870 19488 2926 19544
rect 2778 17584 2834 17640
rect 2962 17584 3018 17640
rect 3421 17434 3477 17436
rect 3501 17434 3557 17436
rect 3581 17434 3637 17436
rect 3661 17434 3717 17436
rect 3421 17382 3447 17434
rect 3447 17382 3477 17434
rect 3501 17382 3511 17434
rect 3511 17382 3557 17434
rect 3581 17382 3627 17434
rect 3627 17382 3637 17434
rect 3661 17382 3691 17434
rect 3691 17382 3717 17434
rect 3421 17380 3477 17382
rect 3501 17380 3557 17382
rect 3581 17380 3637 17382
rect 3661 17380 3717 17382
rect 2686 15680 2742 15736
rect 2594 15408 2650 15464
rect 2778 15000 2834 15056
rect 2410 13252 2466 13288
rect 2410 13232 2412 13252
rect 2412 13232 2464 13252
rect 2464 13232 2466 13252
rect 2134 12416 2190 12472
rect 1950 8472 2006 8528
rect 1858 7248 1914 7304
rect 1674 4800 1730 4856
rect 1674 3984 1730 4040
rect 1674 3304 1730 3360
rect 1858 4120 1914 4176
rect 2318 11620 2374 11656
rect 2318 11600 2320 11620
rect 2320 11600 2372 11620
rect 2372 11600 2374 11620
rect 2870 13912 2926 13968
rect 2686 11736 2742 11792
rect 2502 11056 2558 11112
rect 2502 10956 2504 10976
rect 2504 10956 2556 10976
rect 2556 10956 2558 10976
rect 2502 10920 2558 10956
rect 2502 10668 2558 10704
rect 2502 10648 2504 10668
rect 2504 10648 2556 10668
rect 2556 10648 2558 10668
rect 2502 9832 2558 9888
rect 2226 9424 2282 9480
rect 2134 7792 2190 7848
rect 1858 3848 1914 3904
rect 2226 6840 2282 6896
rect 2410 6024 2466 6080
rect 1306 2488 1362 2544
rect 1122 448 1178 504
rect 1858 1944 1914 2000
rect 3054 14728 3110 14784
rect 3054 12688 3110 12744
rect 2962 12416 3018 12472
rect 2870 9968 2926 10024
rect 2686 9560 2742 9616
rect 2778 9016 2834 9072
rect 2686 8880 2742 8936
rect 2594 7520 2650 7576
rect 2502 5208 2558 5264
rect 2778 5616 2834 5672
rect 3054 8064 3110 8120
rect 3054 7404 3110 7440
rect 3054 7384 3056 7404
rect 3056 7384 3108 7404
rect 3108 7384 3110 7404
rect 3054 6432 3110 6488
rect 2870 4548 2926 4584
rect 2870 4528 2872 4548
rect 2872 4528 2924 4548
rect 2924 4528 2926 4548
rect 2870 4256 2926 4312
rect 2686 2896 2742 2952
rect 2226 1264 2282 1320
rect 3421 16346 3477 16348
rect 3501 16346 3557 16348
rect 3581 16346 3637 16348
rect 3661 16346 3717 16348
rect 3421 16294 3447 16346
rect 3447 16294 3477 16346
rect 3501 16294 3511 16346
rect 3511 16294 3557 16346
rect 3581 16294 3627 16346
rect 3627 16294 3637 16346
rect 3661 16294 3691 16346
rect 3691 16294 3717 16346
rect 3421 16292 3477 16294
rect 3501 16292 3557 16294
rect 3581 16292 3637 16294
rect 3661 16292 3717 16294
rect 4066 18536 4122 18592
rect 3974 16632 4030 16688
rect 3790 15816 3846 15872
rect 3421 15258 3477 15260
rect 3501 15258 3557 15260
rect 3581 15258 3637 15260
rect 3661 15258 3717 15260
rect 3421 15206 3447 15258
rect 3447 15206 3477 15258
rect 3501 15206 3511 15258
rect 3511 15206 3557 15258
rect 3581 15206 3627 15258
rect 3627 15206 3637 15258
rect 3661 15206 3691 15258
rect 3691 15206 3717 15258
rect 3421 15204 3477 15206
rect 3501 15204 3557 15206
rect 3581 15204 3637 15206
rect 3661 15204 3717 15206
rect 4066 16088 4122 16144
rect 4158 15564 4214 15600
rect 4158 15544 4160 15564
rect 4160 15544 4212 15564
rect 4212 15544 4214 15564
rect 3882 15136 3938 15192
rect 3421 14170 3477 14172
rect 3501 14170 3557 14172
rect 3581 14170 3637 14172
rect 3661 14170 3717 14172
rect 3421 14118 3447 14170
rect 3447 14118 3477 14170
rect 3501 14118 3511 14170
rect 3511 14118 3557 14170
rect 3581 14118 3627 14170
rect 3627 14118 3637 14170
rect 3661 14118 3691 14170
rect 3691 14118 3717 14170
rect 3421 14116 3477 14118
rect 3501 14116 3557 14118
rect 3581 14116 3637 14118
rect 3661 14116 3717 14118
rect 3421 13082 3477 13084
rect 3501 13082 3557 13084
rect 3581 13082 3637 13084
rect 3661 13082 3717 13084
rect 3421 13030 3447 13082
rect 3447 13030 3477 13082
rect 3501 13030 3511 13082
rect 3511 13030 3557 13082
rect 3581 13030 3627 13082
rect 3627 13030 3637 13082
rect 3661 13030 3691 13082
rect 3691 13030 3717 13082
rect 3421 13028 3477 13030
rect 3501 13028 3557 13030
rect 3581 13028 3637 13030
rect 3661 13028 3717 13030
rect 3330 12824 3386 12880
rect 3238 12688 3294 12744
rect 3330 12280 3386 12336
rect 3238 7540 3294 7576
rect 3238 7520 3240 7540
rect 3240 7520 3292 7540
rect 3292 7520 3294 7540
rect 3422 12144 3478 12200
rect 3421 11994 3477 11996
rect 3501 11994 3557 11996
rect 3581 11994 3637 11996
rect 3661 11994 3717 11996
rect 3421 11942 3447 11994
rect 3447 11942 3477 11994
rect 3501 11942 3511 11994
rect 3511 11942 3557 11994
rect 3581 11942 3627 11994
rect 3627 11942 3637 11994
rect 3661 11942 3691 11994
rect 3691 11942 3717 11994
rect 3421 11940 3477 11942
rect 3501 11940 3557 11942
rect 3581 11940 3637 11942
rect 3661 11940 3717 11942
rect 3421 10906 3477 10908
rect 3501 10906 3557 10908
rect 3581 10906 3637 10908
rect 3661 10906 3717 10908
rect 3421 10854 3447 10906
rect 3447 10854 3477 10906
rect 3501 10854 3511 10906
rect 3511 10854 3557 10906
rect 3581 10854 3627 10906
rect 3627 10854 3637 10906
rect 3661 10854 3691 10906
rect 3691 10854 3717 10906
rect 3421 10852 3477 10854
rect 3501 10852 3557 10854
rect 3581 10852 3637 10854
rect 3661 10852 3717 10854
rect 3422 9988 3478 10024
rect 3422 9968 3424 9988
rect 3424 9968 3476 9988
rect 3476 9968 3478 9988
rect 3421 9818 3477 9820
rect 3501 9818 3557 9820
rect 3581 9818 3637 9820
rect 3661 9818 3717 9820
rect 3421 9766 3447 9818
rect 3447 9766 3477 9818
rect 3501 9766 3511 9818
rect 3511 9766 3557 9818
rect 3581 9766 3627 9818
rect 3627 9766 3637 9818
rect 3661 9766 3691 9818
rect 3691 9766 3717 9818
rect 3421 9764 3477 9766
rect 3501 9764 3557 9766
rect 3581 9764 3637 9766
rect 3661 9764 3717 9766
rect 3514 9152 3570 9208
rect 3421 8730 3477 8732
rect 3501 8730 3557 8732
rect 3581 8730 3637 8732
rect 3661 8730 3717 8732
rect 3421 8678 3447 8730
rect 3447 8678 3477 8730
rect 3501 8678 3511 8730
rect 3511 8678 3557 8730
rect 3581 8678 3627 8730
rect 3627 8678 3637 8730
rect 3661 8678 3691 8730
rect 3691 8678 3717 8730
rect 3421 8676 3477 8678
rect 3501 8676 3557 8678
rect 3581 8676 3637 8678
rect 3661 8676 3717 8678
rect 3421 7642 3477 7644
rect 3501 7642 3557 7644
rect 3581 7642 3637 7644
rect 3661 7642 3717 7644
rect 3421 7590 3447 7642
rect 3447 7590 3477 7642
rect 3501 7590 3511 7642
rect 3511 7590 3557 7642
rect 3581 7590 3627 7642
rect 3627 7590 3637 7642
rect 3661 7590 3691 7642
rect 3691 7590 3717 7642
rect 3421 7588 3477 7590
rect 3501 7588 3557 7590
rect 3581 7588 3637 7590
rect 3661 7588 3717 7590
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 3790 6296 3846 6352
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 3514 5108 3516 5128
rect 3516 5108 3568 5128
rect 3568 5108 3570 5128
rect 3514 5072 3570 5108
rect 3238 3712 3294 3768
rect 3238 3440 3294 3496
rect 3054 2760 3110 2816
rect 2778 1400 2834 1456
rect 3146 2644 3202 2680
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 3514 4120 3570 4176
rect 3514 3576 3570 3632
rect 3698 4120 3754 4176
rect 3422 3440 3478 3496
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 3514 3032 3570 3088
rect 3422 2760 3478 2816
rect 3146 2624 3148 2644
rect 3148 2624 3200 2644
rect 3200 2624 3202 2644
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 3882 3168 3938 3224
rect 3514 1672 3570 1728
rect 4802 16496 4858 16552
rect 4526 16224 4582 16280
rect 5814 17720 5870 17776
rect 4066 13776 4122 13832
rect 4250 13812 4252 13832
rect 4252 13812 4304 13832
rect 4304 13812 4306 13832
rect 4250 13776 4306 13812
rect 4066 13504 4122 13560
rect 4158 12980 4214 13016
rect 4158 12960 4160 12980
rect 4160 12960 4212 12980
rect 4212 12960 4214 12980
rect 4434 14728 4490 14784
rect 4618 15272 4674 15328
rect 4802 15680 4858 15736
rect 4986 15816 5042 15872
rect 4894 15408 4950 15464
rect 4986 15272 5042 15328
rect 5078 15136 5134 15192
rect 4618 12416 4674 12472
rect 4618 12144 4674 12200
rect 4894 14728 4950 14784
rect 4802 12144 4858 12200
rect 4802 12008 4858 12064
rect 4618 10104 4674 10160
rect 4618 9560 4674 9616
rect 4618 9016 4674 9072
rect 4158 4256 4214 4312
rect 4158 4004 4214 4040
rect 4158 3984 4160 4004
rect 4160 3984 4212 4004
rect 4212 3984 4214 4004
rect 3974 2760 4030 2816
rect 4434 6196 4436 6216
rect 4436 6196 4488 6216
rect 4488 6196 4490 6216
rect 4434 6160 4490 6196
rect 4894 10512 4950 10568
rect 5078 12824 5134 12880
rect 4986 9560 5042 9616
rect 5078 8608 5134 8664
rect 4986 8472 5042 8528
rect 4894 8372 4896 8392
rect 4896 8372 4948 8392
rect 4948 8372 4950 8392
rect 4894 8336 4950 8372
rect 4802 7520 4858 7576
rect 4894 7404 4950 7440
rect 4894 7384 4896 7404
rect 4896 7384 4948 7404
rect 4948 7384 4950 7404
rect 5886 16890 5942 16892
rect 5966 16890 6022 16892
rect 6046 16890 6102 16892
rect 6126 16890 6182 16892
rect 5886 16838 5912 16890
rect 5912 16838 5942 16890
rect 5966 16838 5976 16890
rect 5976 16838 6022 16890
rect 6046 16838 6092 16890
rect 6092 16838 6102 16890
rect 6126 16838 6156 16890
rect 6156 16838 6182 16890
rect 5886 16836 5942 16838
rect 5966 16836 6022 16838
rect 6046 16836 6102 16838
rect 6126 16836 6182 16838
rect 5886 15802 5942 15804
rect 5966 15802 6022 15804
rect 6046 15802 6102 15804
rect 6126 15802 6182 15804
rect 5886 15750 5912 15802
rect 5912 15750 5942 15802
rect 5966 15750 5976 15802
rect 5976 15750 6022 15802
rect 6046 15750 6092 15802
rect 6092 15750 6102 15802
rect 6126 15750 6156 15802
rect 6156 15750 6182 15802
rect 5886 15748 5942 15750
rect 5966 15748 6022 15750
rect 6046 15748 6102 15750
rect 6126 15748 6182 15750
rect 5446 14456 5502 14512
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 6126 14714 6182 14716
rect 5886 14662 5912 14714
rect 5912 14662 5942 14714
rect 5966 14662 5976 14714
rect 5976 14662 6022 14714
rect 6046 14662 6092 14714
rect 6092 14662 6102 14714
rect 6126 14662 6156 14714
rect 6156 14662 6182 14714
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 6126 14660 6182 14662
rect 5354 14356 5356 14376
rect 5356 14356 5408 14376
rect 5408 14356 5410 14376
rect 5354 14320 5410 14356
rect 5262 12824 5318 12880
rect 5262 12300 5318 12336
rect 5262 12280 5264 12300
rect 5264 12280 5316 12300
rect 5316 12280 5318 12300
rect 5446 11872 5502 11928
rect 6366 16496 6422 16552
rect 6550 16940 6552 16960
rect 6552 16940 6604 16960
rect 6604 16940 6606 16960
rect 6550 16904 6606 16940
rect 6458 15680 6514 15736
rect 5630 12688 5686 12744
rect 5722 12588 5724 12608
rect 5724 12588 5776 12608
rect 5776 12588 5778 12608
rect 5722 12552 5778 12588
rect 5262 8064 5318 8120
rect 5354 7520 5410 7576
rect 4894 6704 4950 6760
rect 4802 5364 4858 5400
rect 4802 5344 4804 5364
rect 4804 5344 4856 5364
rect 4856 5344 4858 5364
rect 4710 4392 4766 4448
rect 4250 3168 4306 3224
rect 4526 3476 4528 3496
rect 4528 3476 4580 3496
rect 4580 3476 4582 3496
rect 4526 3440 4582 3476
rect 4342 2216 4398 2272
rect 4618 2508 4674 2544
rect 4618 2488 4620 2508
rect 4620 2488 4672 2508
rect 4672 2488 4674 2508
rect 4802 4256 4858 4312
rect 4986 4256 5042 4312
rect 5262 6704 5318 6760
rect 5722 10784 5778 10840
rect 6090 13776 6146 13832
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 6126 13626 6182 13628
rect 5886 13574 5912 13626
rect 5912 13574 5942 13626
rect 5966 13574 5976 13626
rect 5976 13574 6022 13626
rect 6046 13574 6092 13626
rect 6092 13574 6102 13626
rect 6126 13574 6156 13626
rect 6156 13574 6182 13626
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 6126 13572 6182 13574
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 6126 12538 6182 12540
rect 5886 12486 5912 12538
rect 5912 12486 5942 12538
rect 5966 12486 5976 12538
rect 5976 12486 6022 12538
rect 6046 12486 6092 12538
rect 6092 12486 6102 12538
rect 6126 12486 6156 12538
rect 6156 12486 6182 12538
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 6126 12484 6182 12486
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 6126 11450 6182 11452
rect 5886 11398 5912 11450
rect 5912 11398 5942 11450
rect 5966 11398 5976 11450
rect 5976 11398 6022 11450
rect 6046 11398 6092 11450
rect 6092 11398 6102 11450
rect 6126 11398 6156 11450
rect 6156 11398 6182 11450
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 6126 11396 6182 11398
rect 7286 17176 7342 17232
rect 7194 16652 7250 16688
rect 7194 16632 7196 16652
rect 7196 16632 7248 16652
rect 7248 16632 7250 16652
rect 7010 15816 7066 15872
rect 6826 15136 6882 15192
rect 6918 15000 6974 15056
rect 6826 14592 6882 14648
rect 6826 13812 6828 13832
rect 6828 13812 6880 13832
rect 6880 13812 6882 13832
rect 6826 13776 6882 13812
rect 7286 15272 7342 15328
rect 7194 14728 7250 14784
rect 7102 13388 7158 13424
rect 7102 13368 7104 13388
rect 7104 13368 7156 13388
rect 7156 13368 7158 13388
rect 6642 13132 6644 13152
rect 6644 13132 6696 13152
rect 6696 13132 6698 13152
rect 6642 13096 6698 13132
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 6126 10362 6182 10364
rect 5886 10310 5912 10362
rect 5912 10310 5942 10362
rect 5966 10310 5976 10362
rect 5976 10310 6022 10362
rect 6046 10310 6092 10362
rect 6092 10310 6102 10362
rect 6126 10310 6156 10362
rect 6156 10310 6182 10362
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 6126 10308 6182 10310
rect 6274 9288 6330 9344
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 6126 9274 6182 9276
rect 5886 9222 5912 9274
rect 5912 9222 5942 9274
rect 5966 9222 5976 9274
rect 5976 9222 6022 9274
rect 6046 9222 6092 9274
rect 6092 9222 6102 9274
rect 6126 9222 6156 9274
rect 6156 9222 6182 9274
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 6126 9220 6182 9222
rect 6550 10648 6606 10704
rect 6458 9696 6514 9752
rect 6366 9152 6422 9208
rect 6274 8472 6330 8528
rect 7194 11736 7250 11792
rect 7746 15544 7802 15600
rect 7746 15272 7802 15328
rect 8352 17434 8408 17436
rect 8432 17434 8488 17436
rect 8512 17434 8568 17436
rect 8592 17434 8648 17436
rect 8352 17382 8378 17434
rect 8378 17382 8408 17434
rect 8432 17382 8442 17434
rect 8442 17382 8488 17434
rect 8512 17382 8558 17434
rect 8558 17382 8568 17434
rect 8592 17382 8622 17434
rect 8622 17382 8648 17434
rect 8352 17380 8408 17382
rect 8432 17380 8488 17382
rect 8512 17380 8568 17382
rect 8592 17380 8648 17382
rect 9034 17448 9090 17504
rect 9218 17040 9274 17096
rect 8352 16346 8408 16348
rect 8432 16346 8488 16348
rect 8512 16346 8568 16348
rect 8592 16346 8648 16348
rect 8352 16294 8378 16346
rect 8378 16294 8408 16346
rect 8432 16294 8442 16346
rect 8442 16294 8488 16346
rect 8512 16294 8558 16346
rect 8558 16294 8568 16346
rect 8592 16294 8622 16346
rect 8622 16294 8648 16346
rect 8352 16292 8408 16294
rect 8432 16292 8488 16294
rect 8512 16292 8568 16294
rect 8592 16292 8648 16294
rect 8206 16224 8262 16280
rect 8022 15408 8078 15464
rect 8758 15816 8814 15872
rect 7930 13640 7986 13696
rect 7838 13096 7894 13152
rect 7562 12280 7618 12336
rect 7930 12552 7986 12608
rect 8206 15272 8262 15328
rect 8942 15816 8998 15872
rect 8352 15258 8408 15260
rect 8432 15258 8488 15260
rect 8512 15258 8568 15260
rect 8592 15258 8648 15260
rect 8352 15206 8378 15258
rect 8378 15206 8408 15258
rect 8432 15206 8442 15258
rect 8442 15206 8488 15258
rect 8512 15206 8558 15258
rect 8558 15206 8568 15258
rect 8592 15206 8622 15258
rect 8622 15206 8648 15258
rect 8352 15204 8408 15206
rect 8432 15204 8488 15206
rect 8512 15204 8568 15206
rect 8592 15204 8648 15206
rect 8206 15136 8262 15192
rect 8758 15272 8814 15328
rect 8574 14728 8630 14784
rect 8206 14476 8262 14512
rect 8206 14456 8208 14476
rect 8208 14456 8260 14476
rect 8260 14456 8262 14476
rect 8352 14170 8408 14172
rect 8432 14170 8488 14172
rect 8512 14170 8568 14172
rect 8592 14170 8648 14172
rect 8352 14118 8378 14170
rect 8378 14118 8408 14170
rect 8432 14118 8442 14170
rect 8442 14118 8488 14170
rect 8512 14118 8558 14170
rect 8558 14118 8568 14170
rect 8592 14118 8622 14170
rect 8622 14118 8648 14170
rect 8352 14116 8408 14118
rect 8432 14116 8488 14118
rect 8512 14116 8568 14118
rect 8592 14116 8648 14118
rect 8206 13640 8262 13696
rect 8114 13368 8170 13424
rect 8482 13776 8538 13832
rect 8666 13776 8722 13832
rect 8574 13640 8630 13696
rect 8352 13082 8408 13084
rect 8432 13082 8488 13084
rect 8512 13082 8568 13084
rect 8592 13082 8648 13084
rect 8352 13030 8378 13082
rect 8378 13030 8408 13082
rect 8432 13030 8442 13082
rect 8442 13030 8488 13082
rect 8512 13030 8558 13082
rect 8558 13030 8568 13082
rect 8592 13030 8622 13082
rect 8622 13030 8648 13082
rect 8352 13028 8408 13030
rect 8432 13028 8488 13030
rect 8512 13028 8568 13030
rect 8592 13028 8648 13030
rect 7930 12280 7986 12336
rect 7562 11328 7618 11384
rect 7470 10648 7526 10704
rect 5722 8336 5778 8392
rect 5630 8064 5686 8120
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 6126 8186 6182 8188
rect 5886 8134 5912 8186
rect 5912 8134 5942 8186
rect 5966 8134 5976 8186
rect 5976 8134 6022 8186
rect 6046 8134 6092 8186
rect 6092 8134 6102 8186
rect 6126 8134 6156 8186
rect 6156 8134 6182 8186
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 6126 8132 6182 8134
rect 6734 8336 6790 8392
rect 6274 8064 6330 8120
rect 5814 7656 5870 7712
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 6126 7098 6182 7100
rect 5886 7046 5912 7098
rect 5912 7046 5942 7098
rect 5966 7046 5976 7098
rect 5976 7046 6022 7098
rect 6046 7046 6092 7098
rect 6092 7046 6102 7098
rect 6126 7046 6156 7098
rect 6156 7046 6182 7098
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 6126 7044 6182 7046
rect 5814 6568 5870 6624
rect 6458 7112 6514 7168
rect 6182 6296 6238 6352
rect 5722 6024 5778 6080
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 6366 5888 6422 5944
rect 5354 5636 5410 5672
rect 5354 5616 5356 5636
rect 5356 5616 5408 5636
rect 5408 5616 5410 5636
rect 5354 5344 5410 5400
rect 5722 5616 5778 5672
rect 5354 4936 5410 4992
rect 5354 3440 5410 3496
rect 5354 3168 5410 3224
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 5446 2760 5502 2816
rect 5354 2352 5410 2408
rect 6274 3984 6330 4040
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 5630 2624 5686 2680
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 4986 1536 5042 1592
rect 5538 1128 5594 1184
rect 6734 7656 6790 7712
rect 6642 7384 6698 7440
rect 6642 6432 6698 6488
rect 6918 6568 6974 6624
rect 7470 9968 7526 10024
rect 7378 7792 7434 7848
rect 7286 7520 7342 7576
rect 7562 8472 7618 8528
rect 7838 12008 7894 12064
rect 8942 14728 8998 14784
rect 8942 14320 8998 14376
rect 8850 14184 8906 14240
rect 8942 13912 8998 13968
rect 8850 13640 8906 13696
rect 9218 16652 9274 16688
rect 9218 16632 9220 16652
rect 9220 16632 9272 16652
rect 9272 16632 9274 16652
rect 9218 15816 9274 15872
rect 9586 17312 9642 17368
rect 9494 16496 9550 16552
rect 9586 16224 9642 16280
rect 9954 17312 10010 17368
rect 9770 16632 9826 16688
rect 9402 15816 9458 15872
rect 9126 15308 9128 15328
rect 9128 15308 9180 15328
rect 9180 15308 9182 15328
rect 9126 15272 9182 15308
rect 9126 14456 9182 14512
rect 9218 13096 9274 13152
rect 8666 12416 8722 12472
rect 8352 11994 8408 11996
rect 8432 11994 8488 11996
rect 8512 11994 8568 11996
rect 8592 11994 8648 11996
rect 8352 11942 8378 11994
rect 8378 11942 8408 11994
rect 8432 11942 8442 11994
rect 8442 11942 8488 11994
rect 8512 11942 8558 11994
rect 8558 11942 8568 11994
rect 8592 11942 8622 11994
rect 8622 11942 8648 11994
rect 8352 11940 8408 11942
rect 8432 11940 8488 11942
rect 8512 11940 8568 11942
rect 8592 11940 8648 11942
rect 8206 11872 8262 11928
rect 8114 10784 8170 10840
rect 8352 10906 8408 10908
rect 8432 10906 8488 10908
rect 8512 10906 8568 10908
rect 8592 10906 8648 10908
rect 8352 10854 8378 10906
rect 8378 10854 8408 10906
rect 8432 10854 8442 10906
rect 8442 10854 8488 10906
rect 8512 10854 8558 10906
rect 8558 10854 8568 10906
rect 8592 10854 8622 10906
rect 8622 10854 8648 10906
rect 8352 10852 8408 10854
rect 8432 10852 8488 10854
rect 8512 10852 8568 10854
rect 8592 10852 8648 10854
rect 8114 9968 8170 10024
rect 7746 9696 7802 9752
rect 8022 8744 8078 8800
rect 8022 8492 8078 8528
rect 8022 8472 8024 8492
rect 8024 8472 8076 8492
rect 8076 8472 8078 8492
rect 7654 7520 7710 7576
rect 7378 7112 7434 7168
rect 6826 6024 6882 6080
rect 6642 5072 6698 5128
rect 6550 4004 6606 4040
rect 6550 3984 6552 4004
rect 6552 3984 6604 4004
rect 6604 3984 6606 4004
rect 6826 4392 6882 4448
rect 7010 4392 7066 4448
rect 6734 3848 6790 3904
rect 6734 3304 6790 3360
rect 7286 5072 7342 5128
rect 7194 4936 7250 4992
rect 6734 2760 6790 2816
rect 6826 2624 6882 2680
rect 6182 992 6238 1048
rect 7562 7112 7618 7168
rect 7930 7792 7986 7848
rect 8352 9818 8408 9820
rect 8432 9818 8488 9820
rect 8512 9818 8568 9820
rect 8592 9818 8648 9820
rect 8352 9766 8378 9818
rect 8378 9766 8408 9818
rect 8432 9766 8442 9818
rect 8442 9766 8488 9818
rect 8512 9766 8558 9818
rect 8558 9766 8568 9818
rect 8592 9766 8622 9818
rect 8622 9766 8648 9818
rect 8352 9764 8408 9766
rect 8432 9764 8488 9766
rect 8512 9764 8568 9766
rect 8592 9764 8648 9766
rect 8352 8730 8408 8732
rect 8432 8730 8488 8732
rect 8512 8730 8568 8732
rect 8592 8730 8648 8732
rect 8352 8678 8378 8730
rect 8378 8678 8408 8730
rect 8432 8678 8442 8730
rect 8442 8678 8488 8730
rect 8512 8678 8558 8730
rect 8558 8678 8568 8730
rect 8592 8678 8622 8730
rect 8622 8678 8648 8730
rect 8352 8676 8408 8678
rect 8432 8676 8488 8678
rect 8512 8676 8568 8678
rect 8592 8676 8648 8678
rect 8758 8744 8814 8800
rect 8114 7112 8170 7168
rect 8114 6840 8170 6896
rect 8352 7642 8408 7644
rect 8432 7642 8488 7644
rect 8512 7642 8568 7644
rect 8592 7642 8648 7644
rect 8352 7590 8378 7642
rect 8378 7590 8408 7642
rect 8432 7590 8442 7642
rect 8442 7590 8488 7642
rect 8512 7590 8558 7642
rect 8558 7590 8568 7642
rect 8592 7590 8622 7642
rect 8622 7590 8648 7642
rect 8352 7588 8408 7590
rect 8432 7588 8488 7590
rect 8512 7588 8568 7590
rect 8592 7588 8648 7590
rect 7746 5888 7802 5944
rect 7654 4256 7710 4312
rect 7562 3984 7618 4040
rect 7470 2488 7526 2544
rect 7562 2352 7618 2408
rect 8666 7112 8722 7168
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 8574 5888 8630 5944
rect 8758 6432 8814 6488
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 8758 4392 8814 4448
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 8114 3168 8170 3224
rect 8022 2624 8078 2680
rect 7930 2216 7986 2272
rect 8298 4120 8354 4176
rect 8574 4140 8630 4176
rect 8574 4120 8576 4140
rect 8576 4120 8628 4140
rect 8628 4120 8630 4140
rect 8482 4020 8484 4040
rect 8484 4020 8536 4040
rect 8536 4020 8538 4040
rect 8482 3984 8538 4020
rect 8758 4256 8814 4312
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 9034 12552 9090 12608
rect 9678 15952 9734 16008
rect 9862 14728 9918 14784
rect 9586 14048 9642 14104
rect 10046 16904 10102 16960
rect 10230 16904 10286 16960
rect 10138 16532 10140 16552
rect 10140 16532 10192 16552
rect 10192 16532 10194 16552
rect 10138 16496 10194 16532
rect 10138 16360 10194 16416
rect 10817 16890 10873 16892
rect 10897 16890 10953 16892
rect 10977 16890 11033 16892
rect 11057 16890 11113 16892
rect 10817 16838 10843 16890
rect 10843 16838 10873 16890
rect 10897 16838 10907 16890
rect 10907 16838 10953 16890
rect 10977 16838 11023 16890
rect 11023 16838 11033 16890
rect 11057 16838 11087 16890
rect 11087 16838 11113 16890
rect 10817 16836 10873 16838
rect 10897 16836 10953 16838
rect 10977 16836 11033 16838
rect 11057 16836 11113 16838
rect 10138 15272 10194 15328
rect 10138 14184 10194 14240
rect 9770 12960 9826 13016
rect 9770 12588 9772 12608
rect 9772 12588 9824 12608
rect 9824 12588 9826 12608
rect 9770 12552 9826 12588
rect 9770 12416 9826 12472
rect 9678 12144 9734 12200
rect 10046 14048 10102 14104
rect 9954 12008 10010 12064
rect 9862 11772 9864 11792
rect 9864 11772 9916 11792
rect 9916 11772 9918 11792
rect 9862 11736 9918 11772
rect 9770 10784 9826 10840
rect 9034 9696 9090 9752
rect 9126 9152 9182 9208
rect 9218 7520 9274 7576
rect 9402 9832 9458 9888
rect 9678 9152 9734 9208
rect 9494 8744 9550 8800
rect 9218 6432 9274 6488
rect 9126 6160 9182 6216
rect 9126 5616 9182 5672
rect 9126 5208 9182 5264
rect 9034 4392 9090 4448
rect 8850 2488 8906 2544
rect 8758 2080 8814 2136
rect 9402 5888 9458 5944
rect 9310 3576 9366 3632
rect 9678 8064 9734 8120
rect 9586 7656 9642 7712
rect 9770 7656 9826 7712
rect 9770 6976 9826 7032
rect 9494 4120 9550 4176
rect 9678 4392 9734 4448
rect 9678 4256 9734 4312
rect 9310 2624 9366 2680
rect 8942 1536 8998 1592
rect 9954 11056 10010 11112
rect 10414 15700 10470 15736
rect 10414 15680 10416 15700
rect 10416 15680 10468 15700
rect 10468 15680 10470 15700
rect 10414 15272 10470 15328
rect 10817 15802 10873 15804
rect 10897 15802 10953 15804
rect 10977 15802 11033 15804
rect 11057 15802 11113 15804
rect 10817 15750 10843 15802
rect 10843 15750 10873 15802
rect 10897 15750 10907 15802
rect 10907 15750 10953 15802
rect 10977 15750 11023 15802
rect 11023 15750 11033 15802
rect 11057 15750 11087 15802
rect 11087 15750 11113 15802
rect 10817 15748 10873 15750
rect 10897 15748 10953 15750
rect 10977 15748 11033 15750
rect 11057 15748 11113 15750
rect 10598 15408 10654 15464
rect 10046 9580 10102 9616
rect 10046 9560 10048 9580
rect 10048 9560 10100 9580
rect 10100 9560 10102 9580
rect 10046 8744 10102 8800
rect 10322 11736 10378 11792
rect 10230 8472 10286 8528
rect 10230 7148 10232 7168
rect 10232 7148 10284 7168
rect 10284 7148 10286 7168
rect 10230 7112 10286 7148
rect 10782 15272 10838 15328
rect 11058 15408 11114 15464
rect 10817 14714 10873 14716
rect 10897 14714 10953 14716
rect 10977 14714 11033 14716
rect 11057 14714 11113 14716
rect 10817 14662 10843 14714
rect 10843 14662 10873 14714
rect 10897 14662 10907 14714
rect 10907 14662 10953 14714
rect 10977 14662 11023 14714
rect 11023 14662 11033 14714
rect 11057 14662 11087 14714
rect 11087 14662 11113 14714
rect 10817 14660 10873 14662
rect 10897 14660 10953 14662
rect 10977 14660 11033 14662
rect 11057 14660 11113 14662
rect 11058 14320 11114 14376
rect 10817 13626 10873 13628
rect 10897 13626 10953 13628
rect 10977 13626 11033 13628
rect 11057 13626 11113 13628
rect 10817 13574 10843 13626
rect 10843 13574 10873 13626
rect 10897 13574 10907 13626
rect 10907 13574 10953 13626
rect 10977 13574 11023 13626
rect 11023 13574 11033 13626
rect 11057 13574 11087 13626
rect 11087 13574 11113 13626
rect 10817 13572 10873 13574
rect 10897 13572 10953 13574
rect 10977 13572 11033 13574
rect 11057 13572 11113 13574
rect 10690 12960 10746 13016
rect 10874 12844 10930 12880
rect 10874 12824 10876 12844
rect 10876 12824 10928 12844
rect 10928 12824 10930 12844
rect 10598 12416 10654 12472
rect 10817 12538 10873 12540
rect 10897 12538 10953 12540
rect 10977 12538 11033 12540
rect 11057 12538 11113 12540
rect 10817 12486 10843 12538
rect 10843 12486 10873 12538
rect 10897 12486 10907 12538
rect 10907 12486 10953 12538
rect 10977 12486 11023 12538
rect 11023 12486 11033 12538
rect 11057 12486 11087 12538
rect 11087 12486 11113 12538
rect 10817 12484 10873 12486
rect 10897 12484 10953 12486
rect 10977 12484 11033 12486
rect 11057 12484 11113 12486
rect 10598 12144 10654 12200
rect 10506 11736 10562 11792
rect 10506 11464 10562 11520
rect 10506 11328 10562 11384
rect 10506 10376 10562 10432
rect 10230 5888 10286 5944
rect 10230 5616 10286 5672
rect 10138 4800 10194 4856
rect 10322 5480 10378 5536
rect 10817 11450 10873 11452
rect 10897 11450 10953 11452
rect 10977 11450 11033 11452
rect 11057 11450 11113 11452
rect 10817 11398 10843 11450
rect 10843 11398 10873 11450
rect 10897 11398 10907 11450
rect 10907 11398 10953 11450
rect 10977 11398 11023 11450
rect 11023 11398 11033 11450
rect 11057 11398 11087 11450
rect 11087 11398 11113 11450
rect 10817 11396 10873 11398
rect 10897 11396 10953 11398
rect 10977 11396 11033 11398
rect 11057 11396 11113 11398
rect 11242 15852 11244 15872
rect 11244 15852 11296 15872
rect 11296 15852 11298 15872
rect 11242 15816 11298 15852
rect 11702 17176 11758 17232
rect 11610 16652 11666 16688
rect 11610 16632 11612 16652
rect 11612 16632 11664 16652
rect 11664 16632 11666 16652
rect 11794 16496 11850 16552
rect 11518 15680 11574 15736
rect 11334 12144 11390 12200
rect 11518 15136 11574 15192
rect 11702 16088 11758 16144
rect 11886 15544 11942 15600
rect 11518 14184 11574 14240
rect 11610 13776 11666 13832
rect 11334 11464 11390 11520
rect 10817 10362 10873 10364
rect 10897 10362 10953 10364
rect 10977 10362 11033 10364
rect 11057 10362 11113 10364
rect 10817 10310 10843 10362
rect 10843 10310 10873 10362
rect 10897 10310 10907 10362
rect 10907 10310 10953 10362
rect 10977 10310 11023 10362
rect 11023 10310 11033 10362
rect 11057 10310 11087 10362
rect 11087 10310 11113 10362
rect 10817 10308 10873 10310
rect 10897 10308 10953 10310
rect 10977 10308 11033 10310
rect 11057 10308 11113 10310
rect 10690 9832 10746 9888
rect 10598 9696 10654 9752
rect 11242 9832 11298 9888
rect 10598 9152 10654 9208
rect 10817 9274 10873 9276
rect 10897 9274 10953 9276
rect 10977 9274 11033 9276
rect 11057 9274 11113 9276
rect 10817 9222 10843 9274
rect 10843 9222 10873 9274
rect 10897 9222 10907 9274
rect 10907 9222 10953 9274
rect 10977 9222 11023 9274
rect 11023 9222 11033 9274
rect 11057 9222 11087 9274
rect 11087 9222 11113 9274
rect 10817 9220 10873 9222
rect 10897 9220 10953 9222
rect 10977 9220 11033 9222
rect 11057 9220 11113 9222
rect 10690 8744 10746 8800
rect 11518 11348 11574 11384
rect 11518 11328 11520 11348
rect 11520 11328 11572 11348
rect 11572 11328 11574 11348
rect 11886 13640 11942 13696
rect 13726 17856 13782 17912
rect 13282 17434 13338 17436
rect 13362 17434 13418 17436
rect 13442 17434 13498 17436
rect 13522 17434 13578 17436
rect 13282 17382 13308 17434
rect 13308 17382 13338 17434
rect 13362 17382 13372 17434
rect 13372 17382 13418 17434
rect 13442 17382 13488 17434
rect 13488 17382 13498 17434
rect 13522 17382 13552 17434
rect 13552 17382 13578 17434
rect 13282 17380 13338 17382
rect 13362 17380 13418 17382
rect 13442 17380 13498 17382
rect 13522 17380 13578 17382
rect 13082 17312 13138 17368
rect 12714 16224 12770 16280
rect 12070 15136 12126 15192
rect 11978 13524 12034 13560
rect 11978 13504 11980 13524
rect 11980 13504 12032 13524
rect 12032 13504 12034 13524
rect 11978 13096 12034 13152
rect 11978 12416 12034 12472
rect 11702 11056 11758 11112
rect 12438 15272 12494 15328
rect 12438 14728 12494 14784
rect 12254 14456 12310 14512
rect 12162 12416 12218 12472
rect 11518 10412 11520 10432
rect 11520 10412 11572 10432
rect 11572 10412 11574 10432
rect 11518 10376 11574 10412
rect 11610 10260 11666 10296
rect 11610 10240 11612 10260
rect 11612 10240 11664 10260
rect 11664 10240 11666 10260
rect 11610 9716 11666 9752
rect 11610 9696 11612 9716
rect 11612 9696 11664 9716
rect 11664 9696 11666 9716
rect 10817 8186 10873 8188
rect 10897 8186 10953 8188
rect 10977 8186 11033 8188
rect 11057 8186 11113 8188
rect 10817 8134 10843 8186
rect 10843 8134 10873 8186
rect 10897 8134 10907 8186
rect 10907 8134 10953 8186
rect 10977 8134 11023 8186
rect 11023 8134 11033 8186
rect 11057 8134 11087 8186
rect 11087 8134 11113 8186
rect 10817 8132 10873 8134
rect 10897 8132 10953 8134
rect 10977 8132 11033 8134
rect 11057 8132 11113 8134
rect 11150 7792 11206 7848
rect 11058 7384 11114 7440
rect 10817 7098 10873 7100
rect 10897 7098 10953 7100
rect 10977 7098 11033 7100
rect 11057 7098 11113 7100
rect 10817 7046 10843 7098
rect 10843 7046 10873 7098
rect 10897 7046 10907 7098
rect 10907 7046 10953 7098
rect 10977 7046 11023 7098
rect 11023 7046 11033 7098
rect 11057 7046 11087 7098
rect 11087 7046 11113 7098
rect 10817 7044 10873 7046
rect 10897 7044 10953 7046
rect 10977 7044 11033 7046
rect 11057 7044 11113 7046
rect 11058 6432 11114 6488
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 11426 7656 11482 7712
rect 11426 7384 11482 7440
rect 11334 6024 11390 6080
rect 11334 5908 11390 5944
rect 11334 5888 11336 5908
rect 11336 5888 11388 5908
rect 11388 5888 11390 5908
rect 10966 5616 11022 5672
rect 11242 5616 11298 5672
rect 10690 5480 10746 5536
rect 10414 5208 10470 5264
rect 10414 4936 10470 4992
rect 10414 4140 10470 4176
rect 10414 4120 10416 4140
rect 10416 4120 10468 4140
rect 10468 4120 10470 4140
rect 9954 3712 10010 3768
rect 10138 3848 10194 3904
rect 9402 1264 9458 1320
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 11242 4800 11298 4856
rect 10874 4156 10876 4176
rect 10876 4156 10928 4176
rect 10928 4156 10930 4176
rect 10874 4120 10930 4156
rect 11058 4276 11114 4312
rect 11058 4256 11060 4276
rect 11060 4256 11112 4276
rect 11112 4256 11114 4276
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 10414 2760 10470 2816
rect 10598 2796 10600 2816
rect 10600 2796 10652 2816
rect 10652 2796 10654 2816
rect 10322 2624 10378 2680
rect 9678 1128 9734 1184
rect 10138 992 10194 1048
rect 10598 2760 10654 2796
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 12162 9868 12164 9888
rect 12164 9868 12216 9888
rect 12216 9868 12218 9888
rect 12162 9832 12218 9868
rect 11886 8628 11942 8664
rect 11886 8608 11888 8628
rect 11888 8608 11940 8628
rect 11940 8608 11942 8628
rect 11886 8064 11942 8120
rect 11702 7520 11758 7576
rect 11794 5480 11850 5536
rect 11978 7792 12034 7848
rect 11978 7248 12034 7304
rect 13082 16088 13138 16144
rect 12714 14728 12770 14784
rect 12622 14048 12678 14104
rect 12898 13912 12954 13968
rect 12622 12280 12678 12336
rect 12622 12180 12624 12200
rect 12624 12180 12676 12200
rect 12676 12180 12678 12200
rect 12622 12144 12678 12180
rect 13082 14900 13084 14920
rect 13084 14900 13136 14920
rect 13136 14900 13138 14920
rect 13082 14864 13138 14900
rect 13282 16346 13338 16348
rect 13362 16346 13418 16348
rect 13442 16346 13498 16348
rect 13522 16346 13578 16348
rect 13282 16294 13308 16346
rect 13308 16294 13338 16346
rect 13362 16294 13372 16346
rect 13372 16294 13418 16346
rect 13442 16294 13488 16346
rect 13488 16294 13498 16346
rect 13522 16294 13552 16346
rect 13552 16294 13578 16346
rect 13282 16292 13338 16294
rect 13362 16292 13418 16294
rect 13442 16292 13498 16294
rect 13522 16292 13578 16294
rect 13450 15952 13506 16008
rect 13282 15258 13338 15260
rect 13362 15258 13418 15260
rect 13442 15258 13498 15260
rect 13522 15258 13578 15260
rect 13282 15206 13308 15258
rect 13308 15206 13338 15258
rect 13362 15206 13372 15258
rect 13372 15206 13418 15258
rect 13442 15206 13488 15258
rect 13488 15206 13498 15258
rect 13522 15206 13552 15258
rect 13552 15206 13578 15258
rect 13282 15204 13338 15206
rect 13362 15204 13418 15206
rect 13442 15204 13498 15206
rect 13522 15204 13578 15206
rect 13542 14476 13598 14512
rect 13542 14456 13544 14476
rect 13544 14456 13596 14476
rect 13596 14456 13598 14476
rect 12806 12416 12862 12472
rect 12806 11872 12862 11928
rect 12254 7112 12310 7168
rect 12162 6860 12218 6896
rect 12162 6840 12164 6860
rect 12164 6840 12216 6860
rect 12216 6840 12218 6860
rect 12438 7928 12494 7984
rect 12622 8472 12678 8528
rect 12346 5636 12402 5672
rect 12346 5616 12348 5636
rect 12348 5616 12400 5636
rect 12400 5616 12402 5636
rect 12714 6976 12770 7032
rect 12622 6840 12678 6896
rect 13282 14170 13338 14172
rect 13362 14170 13418 14172
rect 13442 14170 13498 14172
rect 13522 14170 13578 14172
rect 13282 14118 13308 14170
rect 13308 14118 13338 14170
rect 13362 14118 13372 14170
rect 13372 14118 13418 14170
rect 13442 14118 13488 14170
rect 13488 14118 13498 14170
rect 13522 14118 13552 14170
rect 13552 14118 13578 14170
rect 13282 14116 13338 14118
rect 13362 14116 13418 14118
rect 13442 14116 13498 14118
rect 13522 14116 13578 14118
rect 13266 13812 13268 13832
rect 13268 13812 13320 13832
rect 13320 13812 13322 13832
rect 13266 13776 13322 13812
rect 13266 13640 13322 13696
rect 13818 15036 13820 15056
rect 13820 15036 13872 15056
rect 13872 15036 13874 15056
rect 13818 15000 13874 15036
rect 13726 13912 13782 13968
rect 13358 13232 13414 13288
rect 14186 17040 14242 17096
rect 14002 13368 14058 13424
rect 13282 13082 13338 13084
rect 13362 13082 13418 13084
rect 13442 13082 13498 13084
rect 13522 13082 13578 13084
rect 13282 13030 13308 13082
rect 13308 13030 13338 13082
rect 13362 13030 13372 13082
rect 13372 13030 13418 13082
rect 13442 13030 13488 13082
rect 13488 13030 13498 13082
rect 13522 13030 13552 13082
rect 13552 13030 13578 13082
rect 13282 13028 13338 13030
rect 13362 13028 13418 13030
rect 13442 13028 13498 13030
rect 13522 13028 13578 13030
rect 13174 12688 13230 12744
rect 12990 11872 13046 11928
rect 13282 11994 13338 11996
rect 13362 11994 13418 11996
rect 13442 11994 13498 11996
rect 13522 11994 13578 11996
rect 13282 11942 13308 11994
rect 13308 11942 13338 11994
rect 13362 11942 13372 11994
rect 13372 11942 13418 11994
rect 13442 11942 13488 11994
rect 13488 11942 13498 11994
rect 13522 11942 13552 11994
rect 13552 11942 13578 11994
rect 13282 11940 13338 11942
rect 13362 11940 13418 11942
rect 13442 11940 13498 11942
rect 13522 11940 13578 11942
rect 13634 11500 13636 11520
rect 13636 11500 13688 11520
rect 13688 11500 13690 11520
rect 13634 11464 13690 11500
rect 13282 10906 13338 10908
rect 13362 10906 13418 10908
rect 13442 10906 13498 10908
rect 13522 10906 13578 10908
rect 13282 10854 13308 10906
rect 13308 10854 13338 10906
rect 13362 10854 13372 10906
rect 13372 10854 13418 10906
rect 13442 10854 13488 10906
rect 13488 10854 13498 10906
rect 13522 10854 13552 10906
rect 13552 10854 13578 10906
rect 13282 10852 13338 10854
rect 13362 10852 13418 10854
rect 13442 10852 13498 10854
rect 13522 10852 13578 10854
rect 13282 9818 13338 9820
rect 13362 9818 13418 9820
rect 13442 9818 13498 9820
rect 13522 9818 13578 9820
rect 13282 9766 13308 9818
rect 13308 9766 13338 9818
rect 13362 9766 13372 9818
rect 13372 9766 13418 9818
rect 13442 9766 13488 9818
rect 13488 9766 13498 9818
rect 13522 9766 13552 9818
rect 13552 9766 13578 9818
rect 13282 9764 13338 9766
rect 13362 9764 13418 9766
rect 13442 9764 13498 9766
rect 13522 9764 13578 9766
rect 13818 11600 13874 11656
rect 13910 11056 13966 11112
rect 13818 10124 13874 10160
rect 13818 10104 13820 10124
rect 13820 10104 13872 10124
rect 13872 10104 13874 10124
rect 13726 9832 13782 9888
rect 13634 9424 13690 9480
rect 13266 9152 13322 9208
rect 13634 9016 13690 9072
rect 12714 6568 12770 6624
rect 12806 6296 12862 6352
rect 12714 5888 12770 5944
rect 12530 5480 12586 5536
rect 11518 4256 11574 4312
rect 11702 4256 11758 4312
rect 11702 3848 11758 3904
rect 11978 4664 12034 4720
rect 12346 4700 12348 4720
rect 12348 4700 12400 4720
rect 12400 4700 12402 4720
rect 12346 4664 12402 4700
rect 12438 4564 12440 4584
rect 12440 4564 12492 4584
rect 12492 4564 12494 4584
rect 12438 4528 12494 4564
rect 12622 4256 12678 4312
rect 12530 4120 12586 4176
rect 12070 3984 12126 4040
rect 11610 2760 11666 2816
rect 11518 2488 11574 2544
rect 11334 2216 11390 2272
rect 11794 2760 11850 2816
rect 11518 1808 11574 1864
rect 12162 3440 12218 3496
rect 11978 3168 12034 3224
rect 12162 3032 12218 3088
rect 12162 2624 12218 2680
rect 12806 5480 12862 5536
rect 12990 6296 13046 6352
rect 12990 5516 12992 5536
rect 12992 5516 13044 5536
rect 13044 5516 13046 5536
rect 12990 5480 13046 5516
rect 13358 8900 13414 8936
rect 13358 8880 13360 8900
rect 13360 8880 13412 8900
rect 13412 8880 13414 8900
rect 13282 8730 13338 8732
rect 13362 8730 13418 8732
rect 13442 8730 13498 8732
rect 13522 8730 13578 8732
rect 13282 8678 13308 8730
rect 13308 8678 13338 8730
rect 13362 8678 13372 8730
rect 13372 8678 13418 8730
rect 13442 8678 13488 8730
rect 13488 8678 13498 8730
rect 13522 8678 13552 8730
rect 13552 8678 13578 8730
rect 13282 8676 13338 8678
rect 13362 8676 13418 8678
rect 13442 8676 13498 8678
rect 13522 8676 13578 8678
rect 13282 7642 13338 7644
rect 13362 7642 13418 7644
rect 13442 7642 13498 7644
rect 13522 7642 13578 7644
rect 13282 7590 13308 7642
rect 13308 7590 13338 7642
rect 13362 7590 13372 7642
rect 13372 7590 13418 7642
rect 13442 7590 13488 7642
rect 13488 7590 13498 7642
rect 13522 7590 13552 7642
rect 13552 7590 13578 7642
rect 13282 7588 13338 7590
rect 13362 7588 13418 7590
rect 13442 7588 13498 7590
rect 13522 7588 13578 7590
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 13726 6740 13728 6760
rect 13728 6740 13780 6760
rect 13780 6740 13782 6760
rect 13726 6704 13782 6740
rect 13634 6024 13690 6080
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 13174 5208 13230 5264
rect 12806 4664 12862 4720
rect 12990 4120 13046 4176
rect 12898 3612 12900 3632
rect 12900 3612 12952 3632
rect 12952 3612 12954 3632
rect 12898 3576 12954 3612
rect 12806 3304 12862 3360
rect 12622 2644 12678 2680
rect 12622 2624 12624 2644
rect 12624 2624 12676 2644
rect 12676 2624 12678 2644
rect 12530 2352 12586 2408
rect 13082 3304 13138 3360
rect 13082 3168 13138 3224
rect 12806 2216 12862 2272
rect 13266 4936 13322 4992
rect 13450 4936 13506 4992
rect 13358 4800 13414 4856
rect 13634 5072 13690 5128
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 13266 3984 13322 4040
rect 13910 6976 13966 7032
rect 14002 6840 14058 6896
rect 14278 11212 14334 11248
rect 14278 11192 14280 11212
rect 14280 11192 14332 11212
rect 14332 11192 14334 11212
rect 14462 12416 14518 12472
rect 14646 11872 14702 11928
rect 15106 16496 15162 16552
rect 14186 9560 14242 9616
rect 13818 5208 13874 5264
rect 14554 9152 14610 9208
rect 14370 7384 14426 7440
rect 14186 5888 14242 5944
rect 14370 5888 14426 5944
rect 14278 5616 14334 5672
rect 13726 4664 13782 4720
rect 13634 3732 13690 3768
rect 13634 3712 13636 3732
rect 13636 3712 13688 3732
rect 13688 3712 13690 3732
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 13818 3168 13874 3224
rect 13726 2896 13782 2952
rect 14186 3032 14242 3088
rect 13726 2760 13782 2816
rect 12898 1128 12954 1184
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
rect 13818 2488 13874 2544
rect 13818 2216 13874 2272
rect 14002 2624 14058 2680
rect 14646 5752 14702 5808
rect 14554 3440 14610 3496
rect 14094 1944 14150 2000
rect 14278 1672 14334 1728
rect 14278 1536 14334 1592
rect 15106 12416 15162 12472
rect 15014 10512 15070 10568
rect 15014 9968 15070 10024
rect 15014 8336 15070 8392
rect 15106 8200 15162 8256
rect 15014 6160 15070 6216
rect 15014 3884 15016 3904
rect 15016 3884 15068 3904
rect 15068 3884 15070 3904
rect 15014 3848 15070 3884
rect 15474 10648 15530 10704
rect 15014 2760 15070 2816
rect 15566 7248 15622 7304
rect 15106 1400 15162 1456
rect 15566 1944 15622 2000
<< metal3 >>
rect 0 19546 480 19576
rect 2865 19546 2931 19549
rect 0 19544 2931 19546
rect 0 19488 2870 19544
rect 2926 19488 2931 19544
rect 0 19486 2931 19488
rect 0 19456 480 19486
rect 2865 19483 2931 19486
rect 0 18594 480 18624
rect 4061 18594 4127 18597
rect 0 18592 4127 18594
rect 0 18536 4066 18592
rect 4122 18536 4127 18592
rect 0 18534 4127 18536
rect 0 18504 480 18534
rect 4061 18531 4127 18534
rect 13721 17914 13787 17917
rect 16520 17914 17000 17944
rect 13721 17912 17000 17914
rect 13721 17856 13726 17912
rect 13782 17856 17000 17912
rect 13721 17854 17000 17856
rect 13721 17851 13787 17854
rect 16520 17824 17000 17854
rect 5809 17778 5875 17781
rect 8886 17778 8892 17780
rect 5809 17776 8892 17778
rect 5809 17720 5814 17776
rect 5870 17720 8892 17776
rect 5809 17718 8892 17720
rect 5809 17715 5875 17718
rect 8886 17716 8892 17718
rect 8956 17716 8962 17780
rect 0 17642 480 17672
rect 2773 17642 2839 17645
rect 0 17640 2839 17642
rect 0 17584 2778 17640
rect 2834 17584 2839 17640
rect 0 17582 2839 17584
rect 0 17552 480 17582
rect 2773 17579 2839 17582
rect 2957 17642 3023 17645
rect 8150 17642 8156 17644
rect 2957 17640 8156 17642
rect 2957 17584 2962 17640
rect 3018 17584 8156 17640
rect 2957 17582 8156 17584
rect 2957 17579 3023 17582
rect 8150 17580 8156 17582
rect 8220 17580 8226 17644
rect 9029 17506 9095 17509
rect 10358 17506 10364 17508
rect 9029 17504 10364 17506
rect 9029 17448 9034 17504
rect 9090 17448 10364 17504
rect 9029 17446 10364 17448
rect 9029 17443 9095 17446
rect 10358 17444 10364 17446
rect 10428 17444 10434 17508
rect 3409 17440 3729 17441
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 17375 3729 17376
rect 8340 17440 8660 17441
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 17375 8660 17376
rect 13270 17440 13590 17441
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 13270 17375 13590 17376
rect 9581 17370 9647 17373
rect 9949 17370 10015 17373
rect 13077 17370 13143 17373
rect 9581 17368 13143 17370
rect 9581 17312 9586 17368
rect 9642 17312 9954 17368
rect 10010 17312 13082 17368
rect 13138 17312 13143 17368
rect 9581 17310 13143 17312
rect 9581 17307 9647 17310
rect 9949 17307 10015 17310
rect 13077 17307 13143 17310
rect 7281 17234 7347 17237
rect 7966 17234 7972 17236
rect 7281 17232 7972 17234
rect 7281 17176 7286 17232
rect 7342 17176 7972 17232
rect 7281 17174 7972 17176
rect 7281 17171 7347 17174
rect 7966 17172 7972 17174
rect 8036 17234 8042 17236
rect 11697 17234 11763 17237
rect 8036 17232 11763 17234
rect 8036 17176 11702 17232
rect 11758 17176 11763 17232
rect 8036 17174 11763 17176
rect 8036 17172 8042 17174
rect 11697 17171 11763 17174
rect 9213 17098 9279 17101
rect 14181 17098 14247 17101
rect 9213 17096 14247 17098
rect 9213 17040 9218 17096
rect 9274 17040 14186 17096
rect 14242 17040 14247 17096
rect 9213 17038 14247 17040
rect 9213 17035 9279 17038
rect 14181 17035 14247 17038
rect 6545 16962 6611 16965
rect 10041 16962 10107 16965
rect 6545 16960 10107 16962
rect 6545 16904 6550 16960
rect 6606 16904 10046 16960
rect 10102 16904 10107 16960
rect 6545 16902 10107 16904
rect 6545 16899 6611 16902
rect 10041 16899 10107 16902
rect 10225 16962 10291 16965
rect 10542 16962 10548 16964
rect 10225 16960 10548 16962
rect 10225 16904 10230 16960
rect 10286 16904 10548 16960
rect 10225 16902 10548 16904
rect 10225 16899 10291 16902
rect 10542 16900 10548 16902
rect 10612 16900 10618 16964
rect 5874 16896 6194 16897
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6194 16896
rect 5874 16831 6194 16832
rect 10805 16896 11125 16897
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 16831 11125 16832
rect 10174 16826 10180 16828
rect 6272 16766 10180 16826
rect 0 16690 480 16720
rect 2129 16690 2195 16693
rect 0 16688 2195 16690
rect 0 16632 2134 16688
rect 2190 16632 2195 16688
rect 0 16630 2195 16632
rect 0 16600 480 16630
rect 2129 16627 2195 16630
rect 3969 16690 4035 16693
rect 6272 16690 6332 16766
rect 10174 16764 10180 16766
rect 10244 16826 10250 16828
rect 10244 16766 10656 16826
rect 10244 16764 10250 16766
rect 3969 16688 6332 16690
rect 3969 16632 3974 16688
rect 4030 16632 6332 16688
rect 3969 16630 6332 16632
rect 7189 16690 7255 16693
rect 9213 16690 9279 16693
rect 7189 16688 9279 16690
rect 7189 16632 7194 16688
rect 7250 16632 9218 16688
rect 9274 16632 9279 16688
rect 7189 16630 9279 16632
rect 3969 16627 4035 16630
rect 7189 16627 7255 16630
rect 9213 16627 9279 16630
rect 9765 16692 9831 16693
rect 9765 16688 9812 16692
rect 9876 16690 9882 16692
rect 10596 16690 10656 16766
rect 11605 16690 11671 16693
rect 9765 16632 9770 16688
rect 9765 16628 9812 16632
rect 9876 16630 9922 16690
rect 10596 16688 11671 16690
rect 10596 16632 11610 16688
rect 11666 16632 11671 16688
rect 10596 16630 11671 16632
rect 9876 16628 9882 16630
rect 9765 16627 9831 16628
rect 11605 16627 11671 16630
rect 4797 16554 4863 16557
rect 6361 16554 6427 16557
rect 9489 16554 9555 16557
rect 4797 16552 9555 16554
rect 4797 16496 4802 16552
rect 4858 16496 6366 16552
rect 6422 16496 9494 16552
rect 9550 16496 9555 16552
rect 4797 16494 9555 16496
rect 4797 16491 4863 16494
rect 6361 16491 6427 16494
rect 9489 16491 9555 16494
rect 9622 16492 9628 16556
rect 9692 16554 9698 16556
rect 10133 16554 10199 16557
rect 11789 16554 11855 16557
rect 15101 16554 15167 16557
rect 9692 16552 10199 16554
rect 9692 16496 10138 16552
rect 10194 16496 10199 16552
rect 9692 16494 10199 16496
rect 9692 16492 9698 16494
rect 10133 16491 10199 16494
rect 10504 16552 15167 16554
rect 10504 16496 11794 16552
rect 11850 16496 15106 16552
rect 15162 16496 15167 16552
rect 10504 16494 15167 16496
rect 10133 16418 10199 16421
rect 10504 16418 10564 16494
rect 11789 16491 11855 16494
rect 15101 16491 15167 16494
rect 10133 16416 10564 16418
rect 10133 16360 10138 16416
rect 10194 16360 10564 16416
rect 10133 16358 10564 16360
rect 10133 16355 10199 16358
rect 3409 16352 3729 16353
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 16287 3729 16288
rect 8340 16352 8660 16353
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 16287 8660 16288
rect 13270 16352 13590 16353
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 16287 13590 16288
rect 4521 16282 4587 16285
rect 8201 16282 8267 16285
rect 4521 16280 8267 16282
rect 4521 16224 4526 16280
rect 4582 16224 8206 16280
rect 8262 16224 8267 16280
rect 4521 16222 8267 16224
rect 4521 16219 4587 16222
rect 8201 16219 8267 16222
rect 9070 16220 9076 16284
rect 9140 16282 9146 16284
rect 9581 16282 9647 16285
rect 9140 16280 9647 16282
rect 9140 16224 9586 16280
rect 9642 16224 9647 16280
rect 9140 16222 9647 16224
rect 9140 16220 9146 16222
rect 9581 16219 9647 16222
rect 9990 16220 9996 16284
rect 10060 16282 10066 16284
rect 12709 16282 12775 16285
rect 12934 16282 12940 16284
rect 10060 16222 11898 16282
rect 10060 16220 10066 16222
rect 4061 16146 4127 16149
rect 11697 16146 11763 16149
rect 4061 16144 11763 16146
rect 4061 16088 4066 16144
rect 4122 16088 11702 16144
rect 11758 16088 11763 16144
rect 4061 16086 11763 16088
rect 11838 16146 11898 16222
rect 12709 16280 12940 16282
rect 12709 16224 12714 16280
rect 12770 16224 12940 16280
rect 12709 16222 12940 16224
rect 12709 16219 12775 16222
rect 12934 16220 12940 16222
rect 13004 16220 13010 16284
rect 13077 16146 13143 16149
rect 11838 16144 13143 16146
rect 11838 16088 13082 16144
rect 13138 16088 13143 16144
rect 11838 16086 13143 16088
rect 4061 16083 4127 16086
rect 11697 16083 11763 16086
rect 13077 16083 13143 16086
rect 933 16010 999 16013
rect 9673 16010 9739 16013
rect 13445 16010 13511 16013
rect 933 16008 9739 16010
rect 933 15952 938 16008
rect 994 15952 9678 16008
rect 9734 15952 9739 16008
rect 933 15950 9739 15952
rect 933 15947 999 15950
rect 9673 15947 9739 15950
rect 10596 16008 13511 16010
rect 10596 15952 13450 16008
rect 13506 15952 13511 16008
rect 10596 15950 13511 15952
rect 3785 15874 3851 15877
rect 4981 15874 5047 15877
rect 3785 15872 5047 15874
rect 3785 15816 3790 15872
rect 3846 15816 4986 15872
rect 5042 15816 5047 15872
rect 3785 15814 5047 15816
rect 3785 15811 3851 15814
rect 4981 15811 5047 15814
rect 7005 15874 7071 15877
rect 8753 15874 8819 15877
rect 7005 15872 8819 15874
rect 7005 15816 7010 15872
rect 7066 15816 8758 15872
rect 8814 15816 8819 15872
rect 7005 15814 8819 15816
rect 7005 15811 7071 15814
rect 8753 15811 8819 15814
rect 8937 15874 9003 15877
rect 9213 15874 9279 15877
rect 8937 15872 9279 15874
rect 8937 15816 8942 15872
rect 8998 15816 9218 15872
rect 9274 15816 9279 15872
rect 8937 15814 9279 15816
rect 8937 15811 9003 15814
rect 9213 15811 9279 15814
rect 9397 15874 9463 15877
rect 10596 15874 10656 15950
rect 13445 15947 13511 15950
rect 9397 15872 10656 15874
rect 9397 15816 9402 15872
rect 9458 15816 10656 15872
rect 9397 15814 10656 15816
rect 11237 15874 11303 15877
rect 11646 15874 11652 15876
rect 11237 15872 11652 15874
rect 11237 15816 11242 15872
rect 11298 15816 11652 15872
rect 11237 15814 11652 15816
rect 9397 15811 9463 15814
rect 11237 15811 11303 15814
rect 11646 15812 11652 15814
rect 11716 15812 11722 15876
rect 5874 15808 6194 15809
rect 0 15738 480 15768
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6194 15808
rect 5874 15743 6194 15744
rect 10805 15808 11125 15809
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 15743 11125 15744
rect 1853 15738 1919 15741
rect 0 15736 1919 15738
rect 0 15680 1858 15736
rect 1914 15680 1919 15736
rect 0 15678 1919 15680
rect 0 15648 480 15678
rect 1853 15675 1919 15678
rect 2681 15738 2747 15741
rect 4797 15738 4863 15741
rect 2681 15736 4863 15738
rect 2681 15680 2686 15736
rect 2742 15680 4802 15736
rect 4858 15680 4863 15736
rect 2681 15678 4863 15680
rect 2681 15675 2747 15678
rect 4797 15675 4863 15678
rect 6453 15738 6519 15741
rect 10409 15738 10475 15741
rect 6453 15736 10475 15738
rect 6453 15680 6458 15736
rect 6514 15680 10414 15736
rect 10470 15680 10475 15736
rect 6453 15678 10475 15680
rect 6453 15675 6519 15678
rect 10409 15675 10475 15678
rect 11278 15676 11284 15740
rect 11348 15738 11354 15740
rect 11513 15738 11579 15741
rect 11348 15736 11579 15738
rect 11348 15680 11518 15736
rect 11574 15680 11579 15736
rect 11348 15678 11579 15680
rect 11348 15676 11354 15678
rect 11513 15675 11579 15678
rect 4153 15602 4219 15605
rect 7741 15604 7807 15605
rect 7741 15602 7788 15604
rect 4153 15600 7788 15602
rect 7852 15602 7858 15604
rect 4153 15544 4158 15600
rect 4214 15544 7746 15600
rect 4153 15542 7788 15544
rect 4153 15539 4219 15542
rect 7741 15540 7788 15542
rect 7852 15542 7934 15602
rect 7852 15540 7858 15542
rect 8150 15540 8156 15604
rect 8220 15602 8226 15604
rect 11881 15602 11947 15605
rect 8220 15600 11947 15602
rect 8220 15544 11886 15600
rect 11942 15544 11947 15600
rect 8220 15542 11947 15544
rect 8220 15540 8226 15542
rect 7741 15539 7807 15540
rect 11881 15539 11947 15542
rect 2589 15466 2655 15469
rect 3182 15466 3188 15468
rect 2589 15464 3188 15466
rect 2589 15408 2594 15464
rect 2650 15408 3188 15464
rect 2589 15406 3188 15408
rect 2589 15403 2655 15406
rect 3182 15404 3188 15406
rect 3252 15404 3258 15468
rect 4889 15466 4955 15469
rect 8017 15466 8083 15469
rect 4889 15464 9506 15466
rect 4889 15408 4894 15464
rect 4950 15408 8022 15464
rect 8078 15408 9506 15464
rect 4889 15406 9506 15408
rect 4889 15403 4955 15406
rect 8017 15403 8083 15406
rect 4613 15332 4679 15333
rect 4613 15328 4660 15332
rect 4724 15330 4730 15332
rect 4981 15330 5047 15333
rect 7281 15330 7347 15333
rect 7414 15330 7420 15332
rect 4613 15272 4618 15328
rect 4613 15268 4660 15272
rect 4724 15270 4770 15330
rect 4981 15328 7160 15330
rect 4981 15272 4986 15328
rect 5042 15272 7160 15328
rect 4981 15270 7160 15272
rect 4724 15268 4730 15270
rect 4613 15267 4679 15268
rect 4981 15267 5047 15270
rect 3409 15264 3729 15265
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 15199 3729 15200
rect 3877 15194 3943 15197
rect 5073 15194 5139 15197
rect 6821 15194 6887 15197
rect 3877 15192 4906 15194
rect 3877 15136 3882 15192
rect 3938 15136 4906 15192
rect 3877 15134 4906 15136
rect 3877 15131 3943 15134
rect 2773 15060 2839 15061
rect 2773 15056 2820 15060
rect 2884 15058 2890 15060
rect 2773 15000 2778 15056
rect 2773 14996 2820 15000
rect 2884 14998 2930 15058
rect 2884 14996 2890 14998
rect 2773 14995 2839 14996
rect 4846 14922 4906 15134
rect 5073 15192 6887 15194
rect 5073 15136 5078 15192
rect 5134 15136 6826 15192
rect 6882 15136 6887 15192
rect 5073 15134 6887 15136
rect 7100 15194 7160 15270
rect 7281 15328 7420 15330
rect 7281 15272 7286 15328
rect 7342 15272 7420 15328
rect 7281 15270 7420 15272
rect 7281 15267 7347 15270
rect 7414 15268 7420 15270
rect 7484 15268 7490 15332
rect 7741 15330 7807 15333
rect 8201 15330 8267 15333
rect 7741 15328 8267 15330
rect 7741 15272 7746 15328
rect 7802 15272 8206 15328
rect 8262 15272 8267 15328
rect 7741 15270 8267 15272
rect 7741 15267 7807 15270
rect 8201 15267 8267 15270
rect 8753 15330 8819 15333
rect 9121 15330 9187 15333
rect 9446 15332 9506 15406
rect 10358 15404 10364 15468
rect 10428 15466 10434 15468
rect 10593 15466 10659 15469
rect 11053 15466 11119 15469
rect 10428 15464 11119 15466
rect 10428 15408 10598 15464
rect 10654 15408 11058 15464
rect 11114 15408 11119 15464
rect 10428 15406 11119 15408
rect 10428 15404 10434 15406
rect 10593 15403 10659 15406
rect 11053 15403 11119 15406
rect 8753 15328 9187 15330
rect 8753 15272 8758 15328
rect 8814 15272 9126 15328
rect 9182 15272 9187 15328
rect 8753 15270 9187 15272
rect 8753 15267 8819 15270
rect 9121 15267 9187 15270
rect 9438 15268 9444 15332
rect 9508 15330 9514 15332
rect 10133 15330 10199 15333
rect 9508 15328 10199 15330
rect 9508 15272 10138 15328
rect 10194 15272 10199 15328
rect 9508 15270 10199 15272
rect 9508 15268 9514 15270
rect 10133 15267 10199 15270
rect 10409 15330 10475 15333
rect 10777 15330 10843 15333
rect 10409 15328 10843 15330
rect 10409 15272 10414 15328
rect 10470 15272 10782 15328
rect 10838 15272 10843 15328
rect 10409 15270 10843 15272
rect 10409 15267 10475 15270
rect 10777 15267 10843 15270
rect 12433 15330 12499 15333
rect 12750 15330 12756 15332
rect 12433 15328 12756 15330
rect 12433 15272 12438 15328
rect 12494 15272 12756 15328
rect 12433 15270 12756 15272
rect 12433 15267 12499 15270
rect 12750 15268 12756 15270
rect 12820 15268 12826 15332
rect 8340 15264 8660 15265
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 15199 8660 15200
rect 13270 15264 13590 15265
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 15199 13590 15200
rect 8201 15194 8267 15197
rect 7100 15192 8267 15194
rect 7100 15136 8206 15192
rect 8262 15136 8267 15192
rect 7100 15134 8267 15136
rect 5073 15131 5139 15134
rect 6821 15131 6887 15134
rect 8201 15131 8267 15134
rect 8886 15132 8892 15196
rect 8956 15194 8962 15196
rect 9990 15194 9996 15196
rect 8956 15134 9996 15194
rect 8956 15132 8962 15134
rect 9990 15132 9996 15134
rect 10060 15132 10066 15196
rect 10358 15132 10364 15196
rect 10428 15194 10434 15196
rect 11513 15194 11579 15197
rect 10428 15192 11579 15194
rect 10428 15136 11518 15192
rect 11574 15136 11579 15192
rect 10428 15134 11579 15136
rect 10428 15132 10434 15134
rect 11513 15131 11579 15134
rect 12065 15194 12131 15197
rect 12198 15194 12204 15196
rect 12065 15192 12204 15194
rect 12065 15136 12070 15192
rect 12126 15136 12204 15192
rect 12065 15134 12204 15136
rect 12065 15131 12131 15134
rect 12198 15132 12204 15134
rect 12268 15132 12274 15196
rect 6913 15058 6979 15061
rect 13813 15058 13879 15061
rect 6913 15056 13879 15058
rect 6913 15000 6918 15056
rect 6974 15000 13818 15056
rect 13874 15000 13879 15056
rect 6913 14998 13879 15000
rect 6913 14995 6979 14998
rect 13813 14995 13879 14998
rect 10358 14922 10364 14924
rect 4846 14862 10364 14922
rect 10358 14860 10364 14862
rect 10428 14860 10434 14924
rect 13077 14922 13143 14925
rect 10596 14920 13143 14922
rect 10596 14864 13082 14920
rect 13138 14864 13143 14920
rect 10596 14862 13143 14864
rect 0 14786 480 14816
rect 3049 14786 3115 14789
rect 0 14784 3115 14786
rect 0 14728 3054 14784
rect 3110 14728 3115 14784
rect 0 14726 3115 14728
rect 0 14696 480 14726
rect 3049 14723 3115 14726
rect 4429 14786 4495 14789
rect 4889 14786 4955 14789
rect 4429 14784 4955 14786
rect 4429 14728 4434 14784
rect 4490 14728 4894 14784
rect 4950 14728 4955 14784
rect 4429 14726 4955 14728
rect 4429 14723 4495 14726
rect 4889 14723 4955 14726
rect 7189 14786 7255 14789
rect 8569 14786 8635 14789
rect 7189 14784 8635 14786
rect 7189 14728 7194 14784
rect 7250 14728 8574 14784
rect 8630 14728 8635 14784
rect 7189 14726 8635 14728
rect 7189 14723 7255 14726
rect 8569 14723 8635 14726
rect 8937 14786 9003 14789
rect 9857 14786 9923 14789
rect 8937 14784 9923 14786
rect 8937 14728 8942 14784
rect 8998 14728 9862 14784
rect 9918 14728 9923 14784
rect 8937 14726 9923 14728
rect 8937 14723 9003 14726
rect 9857 14723 9923 14726
rect 5874 14720 6194 14721
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6194 14720
rect 5874 14655 6194 14656
rect 6821 14650 6887 14653
rect 9990 14650 9996 14652
rect 6821 14648 9996 14650
rect 6821 14592 6826 14648
rect 6882 14592 9996 14648
rect 6821 14590 9996 14592
rect 6821 14587 6887 14590
rect 9990 14588 9996 14590
rect 10060 14650 10066 14652
rect 10596 14650 10656 14862
rect 13077 14859 13143 14862
rect 12433 14786 12499 14789
rect 12709 14786 12775 14789
rect 13854 14786 13860 14788
rect 12433 14784 13860 14786
rect 12433 14728 12438 14784
rect 12494 14728 12714 14784
rect 12770 14728 13860 14784
rect 12433 14726 13860 14728
rect 12433 14723 12499 14726
rect 12709 14723 12775 14726
rect 13854 14724 13860 14726
rect 13924 14724 13930 14788
rect 10805 14720 11125 14721
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 14655 11125 14656
rect 10060 14590 10656 14650
rect 10060 14588 10066 14590
rect 5441 14514 5507 14517
rect 8201 14514 8267 14517
rect 5441 14512 8267 14514
rect 5441 14456 5446 14512
rect 5502 14456 8206 14512
rect 8262 14456 8267 14512
rect 5441 14454 8267 14456
rect 5441 14451 5507 14454
rect 8201 14451 8267 14454
rect 9121 14514 9187 14517
rect 12249 14514 12315 14517
rect 9121 14512 12315 14514
rect 9121 14456 9126 14512
rect 9182 14456 12254 14512
rect 12310 14456 12315 14512
rect 9121 14454 12315 14456
rect 9121 14451 9187 14454
rect 12249 14451 12315 14454
rect 12934 14452 12940 14516
rect 13004 14514 13010 14516
rect 13537 14514 13603 14517
rect 13004 14512 13603 14514
rect 13004 14456 13542 14512
rect 13598 14456 13603 14512
rect 13004 14454 13603 14456
rect 13004 14452 13010 14454
rect 13537 14451 13603 14454
rect 5349 14378 5415 14381
rect 8937 14378 9003 14381
rect 10358 14378 10364 14380
rect 5349 14376 9003 14378
rect 5349 14320 5354 14376
rect 5410 14320 8942 14376
rect 8998 14320 9003 14376
rect 5349 14318 9003 14320
rect 5349 14315 5415 14318
rect 8937 14315 9003 14318
rect 9400 14318 10364 14378
rect 8845 14242 8911 14245
rect 9400 14242 9460 14318
rect 10358 14316 10364 14318
rect 10428 14378 10434 14380
rect 11053 14378 11119 14381
rect 10428 14376 11119 14378
rect 10428 14320 11058 14376
rect 11114 14320 11119 14376
rect 10428 14318 11119 14320
rect 10428 14316 10434 14318
rect 11053 14315 11119 14318
rect 10133 14244 10199 14245
rect 10133 14242 10180 14244
rect 8845 14240 9460 14242
rect 8845 14184 8850 14240
rect 8906 14184 9460 14240
rect 8845 14182 9460 14184
rect 10088 14240 10180 14242
rect 10088 14184 10138 14240
rect 10088 14182 10180 14184
rect 8845 14179 8911 14182
rect 10133 14180 10180 14182
rect 10244 14180 10250 14244
rect 10542 14180 10548 14244
rect 10612 14242 10618 14244
rect 11513 14242 11579 14245
rect 10612 14240 11579 14242
rect 10612 14184 11518 14240
rect 11574 14184 11579 14240
rect 10612 14182 11579 14184
rect 10612 14180 10618 14182
rect 10133 14179 10242 14180
rect 11513 14179 11579 14182
rect 3409 14176 3729 14177
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 14111 3729 14112
rect 8340 14176 8660 14177
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 14111 8660 14112
rect 9581 14106 9647 14109
rect 10041 14106 10107 14109
rect 9581 14104 10107 14106
rect 9581 14048 9586 14104
rect 9642 14048 10046 14104
rect 10102 14048 10107 14104
rect 9581 14046 10107 14048
rect 10182 14106 10242 14179
rect 13270 14176 13590 14177
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 14111 13590 14112
rect 12617 14106 12683 14109
rect 10182 14104 12683 14106
rect 10182 14048 12622 14104
rect 12678 14048 12683 14104
rect 10182 14046 12683 14048
rect 9581 14043 9647 14046
rect 10041 14043 10107 14046
rect 12617 14043 12683 14046
rect 2865 13970 2931 13973
rect 8937 13970 9003 13973
rect 12893 13970 12959 13973
rect 2865 13968 12959 13970
rect 2865 13912 2870 13968
rect 2926 13912 8942 13968
rect 8998 13912 12898 13968
rect 12954 13912 12959 13968
rect 2865 13910 12959 13912
rect 2865 13907 2931 13910
rect 8937 13907 9003 13910
rect 12893 13907 12959 13910
rect 13721 13970 13787 13973
rect 16520 13970 17000 14000
rect 13721 13968 17000 13970
rect 13721 13912 13726 13968
rect 13782 13912 17000 13968
rect 13721 13910 17000 13912
rect 13721 13907 13787 13910
rect 16520 13880 17000 13910
rect 0 13834 480 13864
rect 4061 13834 4127 13837
rect 0 13832 4127 13834
rect 0 13776 4066 13832
rect 4122 13776 4127 13832
rect 0 13774 4127 13776
rect 0 13744 480 13774
rect 4061 13771 4127 13774
rect 4245 13834 4311 13837
rect 6085 13834 6151 13837
rect 4245 13832 6151 13834
rect 4245 13776 4250 13832
rect 4306 13776 6090 13832
rect 6146 13776 6151 13832
rect 4245 13774 6151 13776
rect 4245 13771 4311 13774
rect 6085 13771 6151 13774
rect 6821 13834 6887 13837
rect 8477 13834 8543 13837
rect 6821 13832 8543 13834
rect 6821 13776 6826 13832
rect 6882 13776 8482 13832
rect 8538 13776 8543 13832
rect 6821 13774 8543 13776
rect 6821 13771 6887 13774
rect 8477 13771 8543 13774
rect 8661 13834 8727 13837
rect 8886 13834 8892 13836
rect 8661 13832 8892 13834
rect 8661 13776 8666 13832
rect 8722 13776 8892 13832
rect 8661 13774 8892 13776
rect 8661 13771 8727 13774
rect 8886 13772 8892 13774
rect 8956 13772 8962 13836
rect 10174 13772 10180 13836
rect 10244 13834 10250 13836
rect 11605 13834 11671 13837
rect 10244 13832 11671 13834
rect 10244 13776 11610 13832
rect 11666 13776 11671 13832
rect 10244 13774 11671 13776
rect 10244 13772 10250 13774
rect 11605 13771 11671 13774
rect 12382 13772 12388 13836
rect 12452 13834 12458 13836
rect 13261 13834 13327 13837
rect 12452 13832 13327 13834
rect 12452 13776 13266 13832
rect 13322 13776 13327 13832
rect 12452 13774 13327 13776
rect 12452 13772 12458 13774
rect 13261 13771 13327 13774
rect 7925 13698 7991 13701
rect 8201 13698 8267 13701
rect 7925 13696 8267 13698
rect 7925 13640 7930 13696
rect 7986 13640 8206 13696
rect 8262 13640 8267 13696
rect 7925 13638 8267 13640
rect 7925 13635 7991 13638
rect 8201 13635 8267 13638
rect 8569 13698 8635 13701
rect 8845 13698 8911 13701
rect 8569 13696 8911 13698
rect 8569 13640 8574 13696
rect 8630 13640 8850 13696
rect 8906 13640 8911 13696
rect 8569 13638 8911 13640
rect 8569 13635 8635 13638
rect 8845 13635 8911 13638
rect 11881 13698 11947 13701
rect 13261 13698 13327 13701
rect 11881 13696 13327 13698
rect 11881 13640 11886 13696
rect 11942 13640 13266 13696
rect 13322 13640 13327 13696
rect 11881 13638 13327 13640
rect 11881 13635 11947 13638
rect 13261 13635 13327 13638
rect 5874 13632 6194 13633
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6194 13632
rect 5874 13567 6194 13568
rect 10805 13632 11125 13633
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 13567 11125 13568
rect 2814 13500 2820 13564
rect 2884 13562 2890 13564
rect 4061 13562 4127 13565
rect 2884 13560 5642 13562
rect 2884 13504 4066 13560
rect 4122 13504 5642 13560
rect 2884 13502 5642 13504
rect 2884 13500 2890 13502
rect 4061 13499 4127 13502
rect 5582 13426 5642 13502
rect 6318 13502 9874 13562
rect 6318 13426 6378 13502
rect 5582 13366 6378 13426
rect 7097 13426 7163 13429
rect 8109 13426 8175 13429
rect 7097 13424 8175 13426
rect 7097 13368 7102 13424
rect 7158 13368 8114 13424
rect 8170 13368 8175 13424
rect 7097 13366 8175 13368
rect 9814 13426 9874 13502
rect 11830 13500 11836 13564
rect 11900 13562 11906 13564
rect 11973 13562 12039 13565
rect 11900 13560 12039 13562
rect 11900 13504 11978 13560
rect 12034 13504 12039 13560
rect 11900 13502 12039 13504
rect 11900 13500 11906 13502
rect 11973 13499 12039 13502
rect 13997 13426 14063 13429
rect 9814 13424 14063 13426
rect 9814 13368 14002 13424
rect 14058 13368 14063 13424
rect 9814 13366 14063 13368
rect 7097 13363 7163 13366
rect 8109 13363 8175 13366
rect 13997 13363 14063 13366
rect 2405 13290 2471 13293
rect 13353 13290 13419 13293
rect 2405 13288 13419 13290
rect 2405 13232 2410 13288
rect 2466 13232 13358 13288
rect 13414 13232 13419 13288
rect 2405 13230 13419 13232
rect 2405 13227 2471 13230
rect 13353 13227 13419 13230
rect 6637 13154 6703 13157
rect 7833 13154 7899 13157
rect 6637 13152 7899 13154
rect 6637 13096 6642 13152
rect 6698 13096 7838 13152
rect 7894 13096 7899 13152
rect 6637 13094 7899 13096
rect 6637 13091 6703 13094
rect 7833 13091 7899 13094
rect 9213 13154 9279 13157
rect 11973 13154 12039 13157
rect 9213 13152 12039 13154
rect 9213 13096 9218 13152
rect 9274 13096 11978 13152
rect 12034 13096 12039 13152
rect 9213 13094 12039 13096
rect 9213 13091 9279 13094
rect 11973 13091 12039 13094
rect 3409 13088 3729 13089
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 13023 3729 13024
rect 8340 13088 8660 13089
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 13023 8660 13024
rect 13270 13088 13590 13089
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 13023 13590 13024
rect 4153 13018 4219 13021
rect 7966 13018 7972 13020
rect 4153 13016 7972 13018
rect 4153 12960 4158 13016
rect 4214 12960 7972 13016
rect 4153 12958 7972 12960
rect 4153 12955 4219 12958
rect 7966 12956 7972 12958
rect 8036 12956 8042 13020
rect 9765 13018 9831 13021
rect 10174 13018 10180 13020
rect 9765 13016 10180 13018
rect 9765 12960 9770 13016
rect 9826 12960 10180 13016
rect 9765 12958 10180 12960
rect 9765 12955 9831 12958
rect 10174 12956 10180 12958
rect 10244 12956 10250 13020
rect 10542 12956 10548 13020
rect 10612 13018 10618 13020
rect 10685 13018 10751 13021
rect 10612 13016 10751 13018
rect 10612 12960 10690 13016
rect 10746 12960 10751 13016
rect 10612 12958 10751 12960
rect 10612 12956 10618 12958
rect 10685 12955 10751 12958
rect 0 12882 480 12912
rect 3325 12882 3391 12885
rect 0 12880 3391 12882
rect 0 12824 3330 12880
rect 3386 12824 3391 12880
rect 0 12822 3391 12824
rect 0 12792 480 12822
rect 3325 12819 3391 12822
rect 5073 12882 5139 12885
rect 5257 12882 5323 12885
rect 10869 12882 10935 12885
rect 5073 12880 10935 12882
rect 5073 12824 5078 12880
rect 5134 12824 5262 12880
rect 5318 12824 10874 12880
rect 10930 12824 10935 12880
rect 5073 12822 10935 12824
rect 5073 12819 5139 12822
rect 5257 12819 5323 12822
rect 10869 12819 10935 12822
rect 3049 12746 3115 12749
rect 3233 12746 3299 12749
rect 3049 12744 3299 12746
rect 3049 12688 3054 12744
rect 3110 12688 3238 12744
rect 3294 12688 3299 12744
rect 3049 12686 3299 12688
rect 3049 12683 3115 12686
rect 3233 12683 3299 12686
rect 5625 12746 5691 12749
rect 13169 12746 13235 12749
rect 5625 12744 13235 12746
rect 5625 12688 5630 12744
rect 5686 12688 13174 12744
rect 13230 12688 13235 12744
rect 5625 12686 13235 12688
rect 5625 12683 5691 12686
rect 13169 12683 13235 12686
rect 1485 12610 1551 12613
rect 5717 12610 5783 12613
rect 1485 12608 5783 12610
rect 1485 12552 1490 12608
rect 1546 12552 5722 12608
rect 5778 12552 5783 12608
rect 1485 12550 5783 12552
rect 1485 12547 1551 12550
rect 5717 12547 5783 12550
rect 7925 12610 7991 12613
rect 9029 12610 9095 12613
rect 9622 12610 9628 12612
rect 7925 12608 9628 12610
rect 7925 12552 7930 12608
rect 7986 12552 9034 12608
rect 9090 12552 9628 12608
rect 7925 12550 9628 12552
rect 7925 12547 7991 12550
rect 9029 12547 9095 12550
rect 9622 12548 9628 12550
rect 9692 12548 9698 12612
rect 9765 12610 9831 12613
rect 10542 12610 10548 12612
rect 9765 12608 10548 12610
rect 9765 12552 9770 12608
rect 9826 12552 10548 12608
rect 9765 12550 10548 12552
rect 9765 12547 9831 12550
rect 10542 12548 10548 12550
rect 10612 12548 10618 12612
rect 5874 12544 6194 12545
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6194 12544
rect 5874 12479 6194 12480
rect 10805 12544 11125 12545
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 12479 11125 12480
rect 2129 12474 2195 12477
rect 2957 12474 3023 12477
rect 4613 12474 4679 12477
rect 2129 12472 4679 12474
rect 2129 12416 2134 12472
rect 2190 12416 2962 12472
rect 3018 12416 4618 12472
rect 4674 12416 4679 12472
rect 2129 12414 4679 12416
rect 2129 12411 2195 12414
rect 2957 12411 3023 12414
rect 4613 12411 4679 12414
rect 7782 12412 7788 12476
rect 7852 12474 7858 12476
rect 8661 12474 8727 12477
rect 7852 12472 8727 12474
rect 7852 12416 8666 12472
rect 8722 12416 8727 12472
rect 7852 12414 8727 12416
rect 7852 12412 7858 12414
rect 8661 12411 8727 12414
rect 9765 12474 9831 12477
rect 10593 12474 10659 12477
rect 9765 12472 10659 12474
rect 9765 12416 9770 12472
rect 9826 12416 10598 12472
rect 10654 12416 10659 12472
rect 9765 12414 10659 12416
rect 9765 12411 9831 12414
rect 10593 12411 10659 12414
rect 11973 12474 12039 12477
rect 12157 12474 12223 12477
rect 11973 12472 12223 12474
rect 11973 12416 11978 12472
rect 12034 12416 12162 12472
rect 12218 12416 12223 12472
rect 11973 12414 12223 12416
rect 11973 12411 12039 12414
rect 12157 12411 12223 12414
rect 12566 12412 12572 12476
rect 12636 12474 12642 12476
rect 12801 12474 12867 12477
rect 12636 12472 12867 12474
rect 12636 12416 12806 12472
rect 12862 12416 12867 12472
rect 12636 12414 12867 12416
rect 12636 12412 12642 12414
rect 12801 12411 12867 12414
rect 14457 12474 14523 12477
rect 15101 12474 15167 12477
rect 14457 12472 15167 12474
rect 14457 12416 14462 12472
rect 14518 12416 15106 12472
rect 15162 12416 15167 12472
rect 14457 12414 15167 12416
rect 14457 12411 14523 12414
rect 15101 12411 15167 12414
rect 3182 12276 3188 12340
rect 3252 12338 3258 12340
rect 3325 12338 3391 12341
rect 3252 12336 3391 12338
rect 3252 12280 3330 12336
rect 3386 12280 3391 12336
rect 3252 12278 3391 12280
rect 3252 12276 3258 12278
rect 3325 12275 3391 12278
rect 5257 12338 5323 12341
rect 7557 12338 7623 12341
rect 7925 12338 7991 12341
rect 12617 12338 12683 12341
rect 5257 12336 12683 12338
rect 5257 12280 5262 12336
rect 5318 12280 7562 12336
rect 7618 12280 7930 12336
rect 7986 12280 12622 12336
rect 12678 12280 12683 12336
rect 5257 12278 12683 12280
rect 5257 12275 5323 12278
rect 7557 12275 7623 12278
rect 7925 12275 7991 12278
rect 12617 12275 12683 12278
rect 3182 12140 3188 12204
rect 3252 12202 3258 12204
rect 3417 12202 3483 12205
rect 4613 12202 4679 12205
rect 3252 12200 4679 12202
rect 3252 12144 3422 12200
rect 3478 12144 4618 12200
rect 4674 12144 4679 12200
rect 3252 12142 4679 12144
rect 3252 12140 3258 12142
rect 3417 12139 3483 12142
rect 4613 12139 4679 12142
rect 4797 12202 4863 12205
rect 9673 12202 9739 12205
rect 10174 12202 10180 12204
rect 4797 12200 8816 12202
rect 4797 12144 4802 12200
rect 4858 12144 8816 12200
rect 4797 12142 8816 12144
rect 4797 12139 4863 12142
rect 4797 12066 4863 12069
rect 7833 12066 7899 12069
rect 4797 12064 7899 12066
rect 4797 12008 4802 12064
rect 4858 12008 7838 12064
rect 7894 12008 7899 12064
rect 4797 12006 7899 12008
rect 4797 12003 4863 12006
rect 7833 12003 7899 12006
rect 3409 12000 3729 12001
rect 0 11930 480 11960
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 11935 3729 11936
rect 8340 12000 8660 12001
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 11935 8660 11936
rect 1853 11930 1919 11933
rect 0 11928 1919 11930
rect 0 11872 1858 11928
rect 1914 11872 1919 11928
rect 0 11870 1919 11872
rect 0 11840 480 11870
rect 1853 11867 1919 11870
rect 4470 11868 4476 11932
rect 4540 11930 4546 11932
rect 5441 11930 5507 11933
rect 4540 11928 5507 11930
rect 4540 11872 5446 11928
rect 5502 11872 5507 11928
rect 4540 11870 5507 11872
rect 4540 11868 4546 11870
rect 5441 11867 5507 11870
rect 5574 11868 5580 11932
rect 5644 11930 5650 11932
rect 8201 11930 8267 11933
rect 5644 11928 8267 11930
rect 5644 11872 8206 11928
rect 8262 11872 8267 11928
rect 5644 11870 8267 11872
rect 8756 11930 8816 12142
rect 9673 12200 10180 12202
rect 9673 12144 9678 12200
rect 9734 12144 10180 12200
rect 9673 12142 10180 12144
rect 9673 12139 9739 12142
rect 10174 12140 10180 12142
rect 10244 12140 10250 12204
rect 10593 12202 10659 12205
rect 11329 12204 11395 12205
rect 11278 12202 11284 12204
rect 10593 12200 11284 12202
rect 11348 12202 11395 12204
rect 11348 12200 11440 12202
rect 10593 12144 10598 12200
rect 10654 12144 11284 12200
rect 11390 12144 11440 12200
rect 10593 12142 11284 12144
rect 10593 12139 10659 12142
rect 11278 12140 11284 12142
rect 11348 12142 11440 12144
rect 11348 12140 11395 12142
rect 12014 12140 12020 12204
rect 12084 12202 12090 12204
rect 12617 12202 12683 12205
rect 12084 12200 12683 12202
rect 12084 12144 12622 12200
rect 12678 12144 12683 12200
rect 12084 12142 12683 12144
rect 12084 12140 12090 12142
rect 11329 12139 11395 12140
rect 12617 12139 12683 12142
rect 9254 12004 9260 12068
rect 9324 12066 9330 12068
rect 9949 12066 10015 12069
rect 9324 12064 10015 12066
rect 9324 12008 9954 12064
rect 10010 12008 10015 12064
rect 9324 12006 10015 12008
rect 9324 12004 9330 12006
rect 9949 12003 10015 12006
rect 13270 12000 13590 12001
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 11935 13590 11936
rect 12801 11930 12867 11933
rect 8756 11928 12867 11930
rect 8756 11872 12806 11928
rect 12862 11872 12867 11928
rect 8756 11870 12867 11872
rect 5644 11868 5650 11870
rect 8201 11867 8267 11870
rect 12801 11867 12867 11870
rect 12985 11930 13051 11933
rect 13118 11930 13124 11932
rect 12985 11928 13124 11930
rect 12985 11872 12990 11928
rect 13046 11872 13124 11928
rect 12985 11870 13124 11872
rect 12985 11867 13051 11870
rect 13118 11868 13124 11870
rect 13188 11868 13194 11932
rect 14641 11930 14707 11933
rect 13678 11928 14707 11930
rect 13678 11872 14646 11928
rect 14702 11872 14707 11928
rect 13678 11870 14707 11872
rect 2681 11794 2747 11797
rect 6862 11794 6868 11796
rect 2681 11792 6868 11794
rect 2681 11736 2686 11792
rect 2742 11736 6868 11792
rect 2681 11734 6868 11736
rect 2681 11731 2747 11734
rect 6862 11732 6868 11734
rect 6932 11732 6938 11796
rect 7189 11794 7255 11797
rect 9857 11794 9923 11797
rect 7189 11792 9923 11794
rect 7189 11736 7194 11792
rect 7250 11736 9862 11792
rect 9918 11736 9923 11792
rect 7189 11734 9923 11736
rect 7189 11731 7255 11734
rect 9857 11731 9923 11734
rect 9990 11732 9996 11796
rect 10060 11794 10066 11796
rect 10317 11794 10383 11797
rect 10060 11792 10383 11794
rect 10060 11736 10322 11792
rect 10378 11736 10383 11792
rect 10060 11734 10383 11736
rect 10060 11732 10066 11734
rect 10317 11731 10383 11734
rect 10501 11794 10567 11797
rect 13678 11794 13738 11870
rect 14641 11867 14707 11870
rect 10501 11792 13738 11794
rect 10501 11736 10506 11792
rect 10562 11736 13738 11792
rect 10501 11734 13738 11736
rect 10501 11731 10567 11734
rect 2313 11658 2379 11661
rect 13813 11658 13879 11661
rect 2313 11656 13879 11658
rect 2313 11600 2318 11656
rect 2374 11600 13818 11656
rect 13874 11600 13879 11656
rect 2313 11598 13879 11600
rect 2313 11595 2379 11598
rect 13813 11595 13879 11598
rect 6862 11460 6868 11524
rect 6932 11522 6938 11524
rect 10501 11522 10567 11525
rect 6932 11520 10567 11522
rect 6932 11464 10506 11520
rect 10562 11464 10567 11520
rect 6932 11462 10567 11464
rect 6932 11460 6938 11462
rect 10501 11459 10567 11462
rect 11329 11522 11395 11525
rect 13629 11522 13695 11525
rect 11329 11520 13695 11522
rect 11329 11464 11334 11520
rect 11390 11464 13634 11520
rect 13690 11464 13695 11520
rect 11329 11462 13695 11464
rect 11329 11459 11395 11462
rect 13629 11459 13695 11462
rect 5874 11456 6194 11457
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6194 11456
rect 5874 11391 6194 11392
rect 10805 11456 11125 11457
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 11391 11125 11392
rect 7557 11386 7623 11389
rect 10501 11386 10567 11389
rect 7557 11384 10567 11386
rect 7557 11328 7562 11384
rect 7618 11328 10506 11384
rect 10562 11328 10567 11384
rect 7557 11326 10567 11328
rect 7557 11323 7623 11326
rect 10501 11323 10567 11326
rect 11278 11324 11284 11388
rect 11348 11386 11354 11388
rect 11513 11386 11579 11389
rect 11348 11384 11579 11386
rect 11348 11328 11518 11384
rect 11574 11328 11579 11384
rect 11348 11326 11579 11328
rect 11348 11324 11354 11326
rect 11513 11323 11579 11326
rect 1761 11250 1827 11253
rect 14273 11250 14339 11253
rect 1761 11248 14339 11250
rect 1761 11192 1766 11248
rect 1822 11192 14278 11248
rect 14334 11192 14339 11248
rect 1761 11190 14339 11192
rect 1761 11187 1827 11190
rect 14273 11187 14339 11190
rect 1761 11114 1827 11117
rect 2497 11114 2563 11117
rect 1761 11112 2563 11114
rect 1761 11056 1766 11112
rect 1822 11056 2502 11112
rect 2558 11056 2563 11112
rect 1761 11054 2563 11056
rect 1761 11051 1827 11054
rect 2497 11051 2563 11054
rect 9949 11116 10015 11117
rect 9949 11112 9996 11116
rect 10060 11114 10066 11116
rect 11697 11114 11763 11117
rect 13905 11114 13971 11117
rect 9949 11056 9954 11112
rect 9949 11052 9996 11056
rect 10060 11054 10106 11114
rect 11697 11112 13971 11114
rect 11697 11056 11702 11112
rect 11758 11056 13910 11112
rect 13966 11056 13971 11112
rect 11697 11054 13971 11056
rect 10060 11052 10066 11054
rect 9949 11051 10015 11052
rect 11697 11051 11763 11054
rect 13905 11051 13971 11054
rect 0 10978 480 11008
rect 2497 10978 2563 10981
rect 0 10976 2563 10978
rect 0 10920 2502 10976
rect 2558 10920 2563 10976
rect 0 10918 2563 10920
rect 0 10888 480 10918
rect 2497 10915 2563 10918
rect 3409 10912 3729 10913
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 10847 3729 10848
rect 8340 10912 8660 10913
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 10847 8660 10848
rect 13270 10912 13590 10913
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 10847 13590 10848
rect 5717 10842 5783 10845
rect 8109 10842 8175 10845
rect 5717 10840 8175 10842
rect 5717 10784 5722 10840
rect 5778 10784 8114 10840
rect 8170 10784 8175 10840
rect 5717 10782 8175 10784
rect 5717 10779 5783 10782
rect 8109 10779 8175 10782
rect 9438 10780 9444 10844
rect 9508 10842 9514 10844
rect 9765 10842 9831 10845
rect 9508 10840 9831 10842
rect 9508 10784 9770 10840
rect 9826 10784 9831 10840
rect 9508 10782 9831 10784
rect 9508 10780 9514 10782
rect 9765 10779 9831 10782
rect 2497 10706 2563 10709
rect 6545 10706 6611 10709
rect 2497 10704 6611 10706
rect 2497 10648 2502 10704
rect 2558 10648 6550 10704
rect 6606 10648 6611 10704
rect 2497 10646 6611 10648
rect 2497 10643 2563 10646
rect 6545 10643 6611 10646
rect 7465 10706 7531 10709
rect 15469 10706 15535 10709
rect 7465 10704 15535 10706
rect 7465 10648 7470 10704
rect 7526 10648 15474 10704
rect 15530 10648 15535 10704
rect 7465 10646 15535 10648
rect 7465 10643 7531 10646
rect 15469 10643 15535 10646
rect 4889 10570 4955 10573
rect 4889 10568 8034 10570
rect 4889 10512 4894 10568
rect 4950 10512 8034 10568
rect 4889 10510 8034 10512
rect 4889 10507 4955 10510
rect 7974 10434 8034 10510
rect 8150 10508 8156 10572
rect 8220 10570 8226 10572
rect 15009 10570 15075 10573
rect 8220 10568 15075 10570
rect 8220 10512 15014 10568
rect 15070 10512 15075 10568
rect 8220 10510 15075 10512
rect 8220 10508 8226 10510
rect 15009 10507 15075 10510
rect 10501 10434 10567 10437
rect 7974 10432 10567 10434
rect 7974 10376 10506 10432
rect 10562 10376 10567 10432
rect 7974 10374 10567 10376
rect 10501 10371 10567 10374
rect 11513 10434 11579 10437
rect 12014 10434 12020 10436
rect 11513 10432 12020 10434
rect 11513 10376 11518 10432
rect 11574 10376 12020 10432
rect 11513 10374 12020 10376
rect 11513 10371 11579 10374
rect 12014 10372 12020 10374
rect 12084 10372 12090 10436
rect 5874 10368 6194 10369
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6194 10368
rect 5874 10303 6194 10304
rect 10805 10368 11125 10369
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 10303 11125 10304
rect 11605 10298 11671 10301
rect 6318 10238 9690 10298
rect 4613 10162 4679 10165
rect 6318 10162 6378 10238
rect 4613 10160 6378 10162
rect 4613 10104 4618 10160
rect 4674 10104 6378 10160
rect 4613 10102 6378 10104
rect 9630 10162 9690 10238
rect 11605 10296 13048 10298
rect 11605 10240 11610 10296
rect 11666 10240 13048 10296
rect 11605 10238 13048 10240
rect 11605 10235 11671 10238
rect 10542 10162 10548 10164
rect 9630 10102 10548 10162
rect 4613 10099 4679 10102
rect 10542 10100 10548 10102
rect 10612 10162 10618 10164
rect 12382 10162 12388 10164
rect 10612 10102 12388 10162
rect 10612 10100 10618 10102
rect 12382 10100 12388 10102
rect 12452 10100 12458 10164
rect 12988 10162 13048 10238
rect 13813 10162 13879 10165
rect 12988 10160 13879 10162
rect 12988 10104 13818 10160
rect 13874 10104 13879 10160
rect 12988 10102 13879 10104
rect 13813 10099 13879 10102
rect 0 10026 480 10056
rect 2865 10026 2931 10029
rect 0 10024 2931 10026
rect 0 9968 2870 10024
rect 2926 9968 2931 10024
rect 0 9966 2931 9968
rect 0 9936 480 9966
rect 2865 9963 2931 9966
rect 3417 10026 3483 10029
rect 7465 10026 7531 10029
rect 3417 10024 7531 10026
rect 3417 9968 3422 10024
rect 3478 9968 7470 10024
rect 7526 9968 7531 10024
rect 3417 9966 7531 9968
rect 3417 9963 3483 9966
rect 7465 9963 7531 9966
rect 8109 10026 8175 10029
rect 15009 10026 15075 10029
rect 8109 10024 15075 10026
rect 8109 9968 8114 10024
rect 8170 9968 15014 10024
rect 15070 9968 15075 10024
rect 8109 9966 15075 9968
rect 8109 9963 8175 9966
rect 15009 9963 15075 9966
rect 1209 9890 1275 9893
rect 2497 9890 2563 9893
rect 1209 9888 2563 9890
rect 1209 9832 1214 9888
rect 1270 9832 2502 9888
rect 2558 9832 2563 9888
rect 1209 9830 2563 9832
rect 1209 9827 1275 9830
rect 2497 9827 2563 9830
rect 9397 9890 9463 9893
rect 10685 9890 10751 9893
rect 9397 9888 10751 9890
rect 9397 9832 9402 9888
rect 9458 9832 10690 9888
rect 10746 9832 10751 9888
rect 9397 9830 10751 9832
rect 9397 9827 9463 9830
rect 10685 9827 10751 9830
rect 11237 9890 11303 9893
rect 12157 9890 12223 9893
rect 11237 9888 12223 9890
rect 11237 9832 11242 9888
rect 11298 9832 12162 9888
rect 12218 9832 12223 9888
rect 11237 9830 12223 9832
rect 11237 9827 11303 9830
rect 12157 9827 12223 9830
rect 13721 9890 13787 9893
rect 16520 9890 17000 9920
rect 13721 9888 17000 9890
rect 13721 9832 13726 9888
rect 13782 9832 17000 9888
rect 13721 9830 17000 9832
rect 13721 9827 13787 9830
rect 3409 9824 3729 9825
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 9759 3729 9760
rect 8340 9824 8660 9825
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 9759 8660 9760
rect 13270 9824 13590 9825
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 16520 9800 17000 9830
rect 13270 9759 13590 9760
rect 6453 9754 6519 9757
rect 7741 9754 7807 9757
rect 6453 9752 7807 9754
rect 6453 9696 6458 9752
rect 6514 9696 7746 9752
rect 7802 9696 7807 9752
rect 6453 9694 7807 9696
rect 6453 9691 6519 9694
rect 7741 9691 7807 9694
rect 9029 9754 9095 9757
rect 10593 9754 10659 9757
rect 11605 9756 11671 9757
rect 11462 9754 11468 9756
rect 9029 9752 10242 9754
rect 9029 9696 9034 9752
rect 9090 9696 10242 9752
rect 9029 9694 10242 9696
rect 9029 9691 9095 9694
rect 2681 9618 2747 9621
rect 4613 9618 4679 9621
rect 2681 9616 4679 9618
rect 2681 9560 2686 9616
rect 2742 9560 4618 9616
rect 4674 9560 4679 9616
rect 2681 9558 4679 9560
rect 2681 9555 2747 9558
rect 4613 9555 4679 9558
rect 4981 9618 5047 9621
rect 10041 9618 10107 9621
rect 4981 9616 10107 9618
rect 4981 9560 4986 9616
rect 5042 9560 10046 9616
rect 10102 9560 10107 9616
rect 4981 9558 10107 9560
rect 10182 9618 10242 9694
rect 10593 9752 11468 9754
rect 10593 9696 10598 9752
rect 10654 9696 11468 9752
rect 10593 9694 11468 9696
rect 10593 9691 10659 9694
rect 11462 9692 11468 9694
rect 11532 9692 11538 9756
rect 11605 9752 11652 9756
rect 11716 9754 11722 9756
rect 11605 9696 11610 9752
rect 11605 9692 11652 9696
rect 11716 9694 11762 9754
rect 11716 9692 11722 9694
rect 11605 9691 11671 9692
rect 14181 9618 14247 9621
rect 14406 9618 14412 9620
rect 10182 9616 14412 9618
rect 10182 9560 14186 9616
rect 14242 9560 14412 9616
rect 10182 9558 14412 9560
rect 4981 9555 5047 9558
rect 10041 9555 10107 9558
rect 14181 9555 14247 9558
rect 14406 9556 14412 9558
rect 14476 9556 14482 9620
rect 2221 9482 2287 9485
rect 13629 9482 13695 9485
rect 2221 9480 13695 9482
rect 2221 9424 2226 9480
rect 2282 9424 13634 9480
rect 13690 9424 13695 9480
rect 2221 9422 13695 9424
rect 2221 9419 2287 9422
rect 13629 9419 13695 9422
rect 6269 9346 6335 9349
rect 10174 9346 10180 9348
rect 6269 9344 10180 9346
rect 6269 9288 6274 9344
rect 6330 9288 10180 9344
rect 6269 9286 10180 9288
rect 6269 9283 6335 9286
rect 10174 9284 10180 9286
rect 10244 9284 10250 9348
rect 5874 9280 6194 9281
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6194 9280
rect 5874 9215 6194 9216
rect 10805 9280 11125 9281
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 9215 11125 9216
rect 2998 9148 3004 9212
rect 3068 9210 3074 9212
rect 3509 9210 3575 9213
rect 6361 9212 6427 9213
rect 3068 9208 3575 9210
rect 3068 9152 3514 9208
rect 3570 9152 3575 9208
rect 3068 9150 3575 9152
rect 3068 9148 3074 9150
rect 3509 9147 3575 9150
rect 6310 9148 6316 9212
rect 6380 9210 6427 9212
rect 6380 9208 6472 9210
rect 6422 9152 6472 9208
rect 6380 9150 6472 9152
rect 6380 9148 6427 9150
rect 6678 9148 6684 9212
rect 6748 9210 6754 9212
rect 9121 9210 9187 9213
rect 6748 9208 9187 9210
rect 6748 9152 9126 9208
rect 9182 9152 9187 9208
rect 6748 9150 9187 9152
rect 6748 9148 6754 9150
rect 6361 9147 6427 9148
rect 9121 9147 9187 9150
rect 9673 9210 9739 9213
rect 10593 9210 10659 9213
rect 9673 9208 10659 9210
rect 9673 9152 9678 9208
rect 9734 9152 10598 9208
rect 10654 9152 10659 9208
rect 9673 9150 10659 9152
rect 9673 9147 9739 9150
rect 10593 9147 10659 9150
rect 13261 9210 13327 9213
rect 14222 9210 14228 9212
rect 13261 9208 14228 9210
rect 13261 9152 13266 9208
rect 13322 9152 14228 9208
rect 13261 9150 14228 9152
rect 13261 9147 13327 9150
rect 14222 9148 14228 9150
rect 14292 9210 14298 9212
rect 14549 9210 14615 9213
rect 14292 9208 14615 9210
rect 14292 9152 14554 9208
rect 14610 9152 14615 9208
rect 14292 9150 14615 9152
rect 14292 9148 14298 9150
rect 14549 9147 14615 9150
rect 0 9074 480 9104
rect 2773 9074 2839 9077
rect 4613 9074 4679 9077
rect 13629 9074 13695 9077
rect 0 9072 2839 9074
rect 0 9016 2778 9072
rect 2834 9016 2839 9072
rect 0 9014 2839 9016
rect 0 8984 480 9014
rect 2773 9011 2839 9014
rect 3374 9014 4538 9074
rect 2681 8938 2747 8941
rect 3374 8938 3434 9014
rect 2681 8936 3434 8938
rect 2681 8880 2686 8936
rect 2742 8880 3434 8936
rect 2681 8878 3434 8880
rect 4478 8938 4538 9014
rect 4613 9072 13695 9074
rect 4613 9016 4618 9072
rect 4674 9016 13634 9072
rect 13690 9016 13695 9072
rect 4613 9014 13695 9016
rect 4613 9011 4679 9014
rect 13629 9011 13695 9014
rect 13353 8938 13419 8941
rect 4478 8936 13419 8938
rect 4478 8880 13358 8936
rect 13414 8880 13419 8936
rect 4478 8878 13419 8880
rect 2681 8875 2747 8878
rect 13353 8875 13419 8878
rect 8017 8802 8083 8805
rect 4662 8800 8083 8802
rect 4662 8744 8022 8800
rect 8078 8744 8083 8800
rect 4662 8742 8083 8744
rect 3409 8736 3729 8737
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 8671 3729 8672
rect 1945 8530 2011 8533
rect 4662 8530 4722 8742
rect 8017 8739 8083 8742
rect 8753 8802 8819 8805
rect 9489 8802 9555 8805
rect 10041 8802 10107 8805
rect 8753 8800 10107 8802
rect 8753 8744 8758 8800
rect 8814 8744 9494 8800
rect 9550 8744 10046 8800
rect 10102 8744 10107 8800
rect 8753 8742 10107 8744
rect 8753 8739 8819 8742
rect 9489 8739 9555 8742
rect 10041 8739 10107 8742
rect 10685 8802 10751 8805
rect 12382 8802 12388 8804
rect 10685 8800 12388 8802
rect 10685 8744 10690 8800
rect 10746 8744 12388 8800
rect 10685 8742 12388 8744
rect 10685 8739 10751 8742
rect 12382 8740 12388 8742
rect 12452 8740 12458 8804
rect 8340 8736 8660 8737
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 8671 8660 8672
rect 13270 8736 13590 8737
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 8671 13590 8672
rect 5073 8666 5139 8669
rect 5073 8664 8264 8666
rect 5073 8608 5078 8664
rect 5134 8608 8264 8664
rect 5073 8606 8264 8608
rect 5073 8603 5139 8606
rect 1945 8528 4722 8530
rect 1945 8472 1950 8528
rect 2006 8472 4722 8528
rect 1945 8470 4722 8472
rect 4981 8530 5047 8533
rect 6269 8530 6335 8533
rect 4981 8528 6335 8530
rect 4981 8472 4986 8528
rect 5042 8472 6274 8528
rect 6330 8472 6335 8528
rect 4981 8470 6335 8472
rect 1945 8467 2011 8470
rect 4981 8467 5047 8470
rect 6269 8467 6335 8470
rect 6494 8468 6500 8532
rect 6564 8530 6570 8532
rect 7557 8530 7623 8533
rect 8017 8532 8083 8533
rect 6564 8528 7623 8530
rect 6564 8472 7562 8528
rect 7618 8472 7623 8528
rect 6564 8470 7623 8472
rect 6564 8468 6570 8470
rect 7557 8467 7623 8470
rect 7966 8468 7972 8532
rect 8036 8530 8083 8532
rect 8204 8530 8264 8606
rect 9990 8604 9996 8668
rect 10060 8666 10066 8668
rect 11646 8666 11652 8668
rect 10060 8606 11652 8666
rect 10060 8604 10066 8606
rect 11646 8604 11652 8606
rect 11716 8604 11722 8668
rect 11881 8666 11947 8669
rect 12014 8666 12020 8668
rect 11881 8664 12020 8666
rect 11881 8608 11886 8664
rect 11942 8608 12020 8664
rect 11881 8606 12020 8608
rect 11881 8603 11947 8606
rect 12014 8604 12020 8606
rect 12084 8604 12090 8668
rect 9622 8530 9628 8532
rect 8036 8528 8128 8530
rect 8078 8472 8128 8528
rect 8036 8470 8128 8472
rect 8204 8470 9628 8530
rect 8036 8468 8083 8470
rect 9622 8468 9628 8470
rect 9692 8468 9698 8532
rect 10225 8530 10291 8533
rect 12617 8530 12683 8533
rect 10225 8528 12683 8530
rect 10225 8472 10230 8528
rect 10286 8472 12622 8528
rect 12678 8472 12683 8528
rect 10225 8470 12683 8472
rect 8017 8467 8083 8468
rect 10225 8467 10291 8470
rect 12617 8467 12683 8470
rect 4889 8394 4955 8397
rect 5717 8394 5783 8397
rect 6729 8394 6795 8397
rect 15009 8394 15075 8397
rect 4889 8392 6332 8394
rect 4889 8336 4894 8392
rect 4950 8336 5722 8392
rect 5778 8336 6332 8392
rect 4889 8334 6332 8336
rect 4889 8331 4955 8334
rect 5717 8331 5783 8334
rect 6272 8258 6332 8334
rect 6729 8392 15075 8394
rect 6729 8336 6734 8392
rect 6790 8336 15014 8392
rect 15070 8336 15075 8392
rect 6729 8334 15075 8336
rect 6729 8331 6795 8334
rect 15009 8331 15075 8334
rect 9254 8258 9260 8260
rect 6272 8198 9260 8258
rect 9254 8196 9260 8198
rect 9324 8196 9330 8260
rect 15101 8258 15167 8261
rect 11286 8256 15167 8258
rect 11286 8200 15106 8256
rect 15162 8200 15167 8256
rect 11286 8198 15167 8200
rect 5874 8192 6194 8193
rect 0 8122 480 8152
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6194 8192
rect 5874 8127 6194 8128
rect 10805 8192 11125 8193
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 8127 11125 8128
rect 3049 8122 3115 8125
rect 0 8120 3115 8122
rect 0 8064 3054 8120
rect 3110 8064 3115 8120
rect 0 8062 3115 8064
rect 0 8032 480 8062
rect 3049 8059 3115 8062
rect 5257 8122 5323 8125
rect 5625 8122 5691 8125
rect 5257 8120 5691 8122
rect 5257 8064 5262 8120
rect 5318 8064 5630 8120
rect 5686 8064 5691 8120
rect 5257 8062 5691 8064
rect 5257 8059 5323 8062
rect 5625 8059 5691 8062
rect 6269 8122 6335 8125
rect 9673 8122 9739 8125
rect 6269 8120 9739 8122
rect 6269 8064 6274 8120
rect 6330 8064 9678 8120
rect 9734 8064 9739 8120
rect 6269 8062 9739 8064
rect 6269 8059 6335 8062
rect 9673 8059 9739 8062
rect 933 7986 999 7989
rect 1393 7986 1459 7989
rect 11286 7986 11346 8198
rect 15101 8195 15167 8198
rect 11881 8124 11947 8125
rect 11830 8060 11836 8124
rect 11900 8122 11947 8124
rect 11900 8120 11992 8122
rect 11942 8064 11992 8120
rect 11900 8062 11992 8064
rect 11900 8060 11947 8062
rect 11881 8059 11947 8060
rect 933 7984 11346 7986
rect 933 7928 938 7984
rect 994 7928 1398 7984
rect 1454 7928 11346 7984
rect 933 7926 11346 7928
rect 933 7923 999 7926
rect 1393 7923 1459 7926
rect 11830 7924 11836 7988
rect 11900 7986 11906 7988
rect 12433 7986 12499 7989
rect 11900 7984 12499 7986
rect 11900 7928 12438 7984
rect 12494 7928 12499 7984
rect 11900 7926 12499 7928
rect 11900 7924 11906 7926
rect 12433 7923 12499 7926
rect 2129 7850 2195 7853
rect 7373 7850 7439 7853
rect 2129 7848 7439 7850
rect 2129 7792 2134 7848
rect 2190 7792 7378 7848
rect 7434 7792 7439 7848
rect 2129 7790 7439 7792
rect 2129 7787 2195 7790
rect 7373 7787 7439 7790
rect 7925 7850 7991 7853
rect 11145 7850 11211 7853
rect 11973 7850 12039 7853
rect 12566 7850 12572 7852
rect 7925 7848 12572 7850
rect 7925 7792 7930 7848
rect 7986 7792 11150 7848
rect 11206 7792 11978 7848
rect 12034 7792 12572 7848
rect 7925 7790 12572 7792
rect 7925 7787 7991 7790
rect 11145 7787 11211 7790
rect 11973 7787 12039 7790
rect 12566 7788 12572 7790
rect 12636 7788 12642 7852
rect 5206 7652 5212 7716
rect 5276 7714 5282 7716
rect 5809 7714 5875 7717
rect 5276 7712 5875 7714
rect 5276 7656 5814 7712
rect 5870 7656 5875 7712
rect 5276 7654 5875 7656
rect 5276 7652 5282 7654
rect 5809 7651 5875 7654
rect 6729 7714 6795 7717
rect 7966 7714 7972 7716
rect 6729 7712 7972 7714
rect 6729 7656 6734 7712
rect 6790 7656 7972 7712
rect 6729 7654 7972 7656
rect 6729 7651 6795 7654
rect 7966 7652 7972 7654
rect 8036 7652 8042 7716
rect 9254 7652 9260 7716
rect 9324 7714 9330 7716
rect 9581 7714 9647 7717
rect 9324 7712 9647 7714
rect 9324 7656 9586 7712
rect 9642 7656 9647 7712
rect 9324 7654 9647 7656
rect 9324 7652 9330 7654
rect 9581 7651 9647 7654
rect 9765 7714 9831 7717
rect 11421 7714 11487 7717
rect 9765 7712 11487 7714
rect 9765 7656 9770 7712
rect 9826 7656 11426 7712
rect 11482 7656 11487 7712
rect 9765 7654 11487 7656
rect 9765 7651 9831 7654
rect 11421 7651 11487 7654
rect 3409 7648 3729 7649
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 7583 3729 7584
rect 8340 7648 8660 7649
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 7583 8660 7584
rect 13270 7648 13590 7649
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 7583 13590 7584
rect 2589 7578 2655 7581
rect 3233 7578 3299 7581
rect 2589 7576 3299 7578
rect 2589 7520 2594 7576
rect 2650 7520 3238 7576
rect 3294 7520 3299 7576
rect 2589 7518 3299 7520
rect 2589 7515 2655 7518
rect 3233 7515 3299 7518
rect 4797 7580 4863 7581
rect 4797 7576 4844 7580
rect 4908 7578 4914 7580
rect 5349 7578 5415 7581
rect 7281 7578 7347 7581
rect 7649 7580 7715 7581
rect 7598 7578 7604 7580
rect 4797 7520 4802 7576
rect 4797 7516 4844 7520
rect 4908 7518 4954 7578
rect 5349 7576 7347 7578
rect 5349 7520 5354 7576
rect 5410 7520 7286 7576
rect 7342 7520 7347 7576
rect 5349 7518 7347 7520
rect 7558 7518 7604 7578
rect 7668 7576 7715 7580
rect 7710 7520 7715 7576
rect 4908 7516 4914 7518
rect 4797 7515 4863 7516
rect 5349 7515 5415 7518
rect 7281 7515 7347 7518
rect 7598 7516 7604 7518
rect 7668 7516 7715 7520
rect 7649 7515 7715 7516
rect 9213 7578 9279 7581
rect 11697 7578 11763 7581
rect 9213 7576 11763 7578
rect 9213 7520 9218 7576
rect 9274 7520 11702 7576
rect 11758 7520 11763 7576
rect 9213 7518 11763 7520
rect 9213 7515 9279 7518
rect 11697 7515 11763 7518
rect 3049 7442 3115 7445
rect 4889 7442 4955 7445
rect 3049 7440 4955 7442
rect 3049 7384 3054 7440
rect 3110 7384 4894 7440
rect 4950 7384 4955 7440
rect 3049 7382 4955 7384
rect 3049 7379 3115 7382
rect 4889 7379 4955 7382
rect 5022 7380 5028 7444
rect 5092 7442 5098 7444
rect 6494 7442 6500 7444
rect 5092 7382 6500 7442
rect 5092 7380 5098 7382
rect 6494 7380 6500 7382
rect 6564 7380 6570 7444
rect 6637 7442 6703 7445
rect 11053 7442 11119 7445
rect 6637 7440 11119 7442
rect 6637 7384 6642 7440
rect 6698 7384 11058 7440
rect 11114 7384 11119 7440
rect 6637 7382 11119 7384
rect 6637 7379 6703 7382
rect 11053 7379 11119 7382
rect 11421 7442 11487 7445
rect 14365 7442 14431 7445
rect 11421 7440 14431 7442
rect 11421 7384 11426 7440
rect 11482 7384 14370 7440
rect 14426 7384 14431 7440
rect 11421 7382 14431 7384
rect 11421 7379 11487 7382
rect 14365 7379 14431 7382
rect 1853 7306 1919 7309
rect 11973 7306 12039 7309
rect 1853 7304 12039 7306
rect 1853 7248 1858 7304
rect 1914 7248 11978 7304
rect 12034 7248 12039 7304
rect 1853 7246 12039 7248
rect 1853 7243 1919 7246
rect 11973 7243 12039 7246
rect 13118 7244 13124 7308
rect 13188 7306 13194 7308
rect 15561 7306 15627 7309
rect 13188 7304 15627 7306
rect 13188 7248 15566 7304
rect 15622 7248 15627 7304
rect 13188 7246 15627 7248
rect 13188 7244 13194 7246
rect 15561 7243 15627 7246
rect 0 7170 480 7200
rect 749 7170 815 7173
rect 0 7168 815 7170
rect 0 7112 754 7168
rect 810 7112 815 7168
rect 0 7110 815 7112
rect 0 7080 480 7110
rect 749 7107 815 7110
rect 6453 7170 6519 7173
rect 7230 7170 7236 7172
rect 6453 7168 7236 7170
rect 6453 7112 6458 7168
rect 6514 7112 7236 7168
rect 6453 7110 7236 7112
rect 6453 7107 6519 7110
rect 7230 7108 7236 7110
rect 7300 7170 7306 7172
rect 7373 7170 7439 7173
rect 7300 7168 7439 7170
rect 7300 7112 7378 7168
rect 7434 7112 7439 7168
rect 7300 7110 7439 7112
rect 7300 7108 7306 7110
rect 7373 7107 7439 7110
rect 7557 7170 7623 7173
rect 8109 7170 8175 7173
rect 7557 7168 8175 7170
rect 7557 7112 7562 7168
rect 7618 7112 8114 7168
rect 8170 7112 8175 7168
rect 7557 7110 8175 7112
rect 7557 7107 7623 7110
rect 8109 7107 8175 7110
rect 8661 7170 8727 7173
rect 10225 7170 10291 7173
rect 8661 7168 10291 7170
rect 8661 7112 8666 7168
rect 8722 7112 10230 7168
rect 10286 7112 10291 7168
rect 8661 7110 10291 7112
rect 8661 7107 8727 7110
rect 10225 7107 10291 7110
rect 12249 7170 12315 7173
rect 14038 7170 14044 7172
rect 12249 7168 14044 7170
rect 12249 7112 12254 7168
rect 12310 7112 14044 7168
rect 12249 7110 14044 7112
rect 12249 7107 12315 7110
rect 14038 7108 14044 7110
rect 14108 7108 14114 7172
rect 5874 7104 6194 7105
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6194 7104
rect 5874 7039 6194 7040
rect 10805 7104 11125 7105
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 7039 11125 7040
rect 6494 6972 6500 7036
rect 6564 7034 6570 7036
rect 9765 7034 9831 7037
rect 6564 7032 9831 7034
rect 6564 6976 9770 7032
rect 9826 6976 9831 7032
rect 6564 6974 9831 6976
rect 6564 6972 6570 6974
rect 9765 6971 9831 6974
rect 11240 6974 12404 7034
rect 2221 6898 2287 6901
rect 7598 6898 7604 6900
rect 2221 6896 7604 6898
rect 2221 6840 2226 6896
rect 2282 6840 7604 6896
rect 2221 6838 7604 6840
rect 2221 6835 2287 6838
rect 7598 6836 7604 6838
rect 7668 6836 7674 6900
rect 7966 6836 7972 6900
rect 8036 6898 8042 6900
rect 8109 6898 8175 6901
rect 11240 6898 11300 6974
rect 8036 6896 11300 6898
rect 8036 6840 8114 6896
rect 8170 6840 11300 6896
rect 8036 6838 11300 6840
rect 8036 6836 8042 6838
rect 8109 6835 8175 6838
rect 11646 6836 11652 6900
rect 11716 6898 11722 6900
rect 12157 6898 12223 6901
rect 11716 6896 12223 6898
rect 11716 6840 12162 6896
rect 12218 6840 12223 6896
rect 11716 6838 12223 6840
rect 12344 6898 12404 6974
rect 12566 6972 12572 7036
rect 12636 7034 12642 7036
rect 12709 7034 12775 7037
rect 13905 7034 13971 7037
rect 12636 7032 13971 7034
rect 12636 6976 12714 7032
rect 12770 6976 13910 7032
rect 13966 6976 13971 7032
rect 12636 6974 13971 6976
rect 12636 6972 12642 6974
rect 12709 6971 12775 6974
rect 13905 6971 13971 6974
rect 12617 6898 12683 6901
rect 12344 6896 12683 6898
rect 12344 6840 12622 6896
rect 12678 6840 12683 6896
rect 12344 6838 12683 6840
rect 11716 6836 11722 6838
rect 12157 6835 12223 6838
rect 12617 6835 12683 6838
rect 13670 6836 13676 6900
rect 13740 6898 13746 6900
rect 13997 6898 14063 6901
rect 13740 6896 14063 6898
rect 13740 6840 14002 6896
rect 14058 6840 14063 6896
rect 13740 6838 14063 6840
rect 13740 6836 13746 6838
rect 13997 6835 14063 6838
rect 4889 6760 4955 6765
rect 4889 6704 4894 6760
rect 4950 6704 4955 6760
rect 4889 6699 4955 6704
rect 5257 6762 5323 6765
rect 5257 6760 9736 6762
rect 5257 6704 5262 6760
rect 5318 6704 9736 6760
rect 5257 6702 9736 6704
rect 5257 6699 5323 6702
rect 4892 6626 4952 6699
rect 5809 6626 5875 6629
rect 4892 6624 5875 6626
rect 4892 6568 5814 6624
rect 5870 6568 5875 6624
rect 4892 6566 5875 6568
rect 5809 6563 5875 6566
rect 6913 6626 6979 6629
rect 7046 6626 7052 6628
rect 6913 6624 7052 6626
rect 6913 6568 6918 6624
rect 6974 6568 7052 6624
rect 6913 6566 7052 6568
rect 6913 6563 6979 6566
rect 7046 6564 7052 6566
rect 7116 6564 7122 6628
rect 9676 6626 9736 6702
rect 9806 6700 9812 6764
rect 9876 6762 9882 6764
rect 13721 6762 13787 6765
rect 9876 6760 13787 6762
rect 9876 6704 13726 6760
rect 13782 6704 13787 6760
rect 9876 6702 13787 6704
rect 9876 6700 9882 6702
rect 13721 6699 13787 6702
rect 12709 6626 12775 6629
rect 9676 6624 12775 6626
rect 9676 6568 12714 6624
rect 12770 6568 12775 6624
rect 9676 6566 12775 6568
rect 12709 6563 12775 6566
rect 3409 6560 3729 6561
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 3049 6492 3115 6493
rect 2998 6428 3004 6492
rect 3068 6490 3115 6492
rect 6637 6490 6703 6493
rect 7966 6490 7972 6492
rect 3068 6488 3160 6490
rect 3110 6432 3160 6488
rect 3068 6430 3160 6432
rect 6637 6488 7972 6490
rect 6637 6432 6642 6488
rect 6698 6432 7972 6488
rect 6637 6430 7972 6432
rect 3068 6428 3115 6430
rect 3049 6427 3115 6428
rect 6637 6427 6703 6430
rect 7966 6428 7972 6430
rect 8036 6428 8042 6492
rect 8753 6490 8819 6493
rect 9213 6490 9279 6493
rect 8753 6488 9279 6490
rect 8753 6432 8758 6488
rect 8814 6432 9218 6488
rect 9274 6432 9279 6488
rect 8753 6430 9279 6432
rect 8753 6427 8819 6430
rect 9213 6427 9279 6430
rect 9806 6428 9812 6492
rect 9876 6490 9882 6492
rect 11053 6490 11119 6493
rect 9876 6488 11119 6490
rect 9876 6432 11058 6488
rect 11114 6432 11119 6488
rect 9876 6430 11119 6432
rect 9876 6428 9882 6430
rect 11053 6427 11119 6430
rect 3785 6354 3851 6357
rect 6177 6354 6243 6357
rect 3785 6352 6243 6354
rect 3785 6296 3790 6352
rect 3846 6296 6182 6352
rect 6238 6296 6243 6352
rect 3785 6294 6243 6296
rect 3785 6291 3851 6294
rect 6177 6291 6243 6294
rect 6310 6292 6316 6356
rect 6380 6354 6386 6356
rect 12801 6354 12867 6357
rect 6380 6352 12867 6354
rect 6380 6296 12806 6352
rect 12862 6296 12867 6352
rect 6380 6294 12867 6296
rect 6380 6292 6386 6294
rect 12801 6291 12867 6294
rect 12985 6354 13051 6357
rect 13854 6354 13860 6356
rect 12985 6352 13860 6354
rect 12985 6296 12990 6352
rect 13046 6296 13860 6352
rect 12985 6294 13860 6296
rect 12985 6291 13051 6294
rect 13854 6292 13860 6294
rect 13924 6292 13930 6356
rect 0 6218 480 6248
rect 4286 6218 4292 6220
rect 0 6158 4292 6218
rect 0 6128 480 6158
rect 4286 6156 4292 6158
rect 4356 6156 4362 6220
rect 4429 6218 4495 6221
rect 9121 6218 9187 6221
rect 15009 6218 15075 6221
rect 4429 6216 9187 6218
rect 4429 6160 4434 6216
rect 4490 6160 9126 6216
rect 9182 6160 9187 6216
rect 4429 6158 9187 6160
rect 4429 6155 4495 6158
rect 9121 6155 9187 6158
rect 9400 6216 15075 6218
rect 9400 6160 15014 6216
rect 15070 6160 15075 6216
rect 9400 6158 15075 6160
rect 2405 6082 2471 6085
rect 5717 6082 5783 6085
rect 2405 6080 5783 6082
rect 2405 6024 2410 6080
rect 2466 6024 5722 6080
rect 5778 6024 5783 6080
rect 2405 6022 5783 6024
rect 2405 6019 2471 6022
rect 5717 6019 5783 6022
rect 6821 6082 6887 6085
rect 9400 6082 9460 6158
rect 15009 6155 15075 6158
rect 6821 6080 9460 6082
rect 6821 6024 6826 6080
rect 6882 6024 9460 6080
rect 6821 6022 9460 6024
rect 11329 6082 11395 6085
rect 13629 6082 13695 6085
rect 11329 6080 13695 6082
rect 11329 6024 11334 6080
rect 11390 6024 13634 6080
rect 13690 6024 13695 6080
rect 11329 6022 13695 6024
rect 6821 6019 6887 6022
rect 11329 6019 11395 6022
rect 13629 6019 13695 6022
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 6361 5946 6427 5949
rect 7741 5946 7807 5949
rect 6361 5944 7807 5946
rect 6361 5888 6366 5944
rect 6422 5888 7746 5944
rect 7802 5888 7807 5944
rect 6361 5886 7807 5888
rect 6361 5883 6427 5886
rect 7741 5883 7807 5886
rect 7966 5884 7972 5948
rect 8036 5946 8042 5948
rect 8569 5946 8635 5949
rect 8036 5944 8635 5946
rect 8036 5888 8574 5944
rect 8630 5888 8635 5944
rect 8036 5886 8635 5888
rect 8036 5884 8042 5886
rect 8569 5883 8635 5886
rect 9397 5946 9463 5949
rect 10225 5946 10291 5949
rect 9397 5944 10291 5946
rect 9397 5888 9402 5944
rect 9458 5888 10230 5944
rect 10286 5888 10291 5944
rect 9397 5886 10291 5888
rect 9397 5883 9463 5886
rect 10225 5883 10291 5886
rect 11329 5946 11395 5949
rect 11830 5946 11836 5948
rect 11329 5944 11836 5946
rect 11329 5888 11334 5944
rect 11390 5888 11836 5944
rect 11329 5886 11836 5888
rect 11329 5883 11395 5886
rect 11830 5884 11836 5886
rect 11900 5884 11906 5948
rect 12566 5884 12572 5948
rect 12636 5946 12642 5948
rect 12709 5946 12775 5949
rect 12636 5944 12775 5946
rect 12636 5888 12714 5944
rect 12770 5888 12775 5944
rect 12636 5886 12775 5888
rect 12636 5884 12642 5886
rect 12709 5883 12775 5886
rect 12934 5884 12940 5948
rect 13004 5946 13010 5948
rect 14181 5946 14247 5949
rect 13004 5944 14247 5946
rect 13004 5888 14186 5944
rect 14242 5888 14247 5944
rect 13004 5886 14247 5888
rect 13004 5884 13010 5886
rect 14181 5883 14247 5886
rect 14365 5946 14431 5949
rect 16520 5946 17000 5976
rect 14365 5944 17000 5946
rect 14365 5888 14370 5944
rect 14426 5888 17000 5944
rect 14365 5886 17000 5888
rect 14365 5883 14431 5886
rect 16520 5856 17000 5886
rect 1393 5810 1459 5813
rect 7414 5810 7420 5812
rect 1393 5808 7420 5810
rect 1393 5752 1398 5808
rect 1454 5752 7420 5808
rect 1393 5750 7420 5752
rect 1393 5747 1459 5750
rect 7414 5748 7420 5750
rect 7484 5748 7490 5812
rect 7598 5748 7604 5812
rect 7668 5810 7674 5812
rect 14641 5810 14707 5813
rect 7668 5808 14707 5810
rect 7668 5752 14646 5808
rect 14702 5752 14707 5808
rect 7668 5750 14707 5752
rect 7668 5748 7674 5750
rect 14641 5747 14707 5750
rect 2773 5674 2839 5677
rect 5349 5676 5415 5677
rect 2773 5672 5274 5674
rect 2773 5616 2778 5672
rect 2834 5616 5274 5672
rect 2773 5614 5274 5616
rect 2773 5611 2839 5614
rect 5214 5538 5274 5614
rect 5349 5672 5396 5676
rect 5460 5674 5466 5676
rect 5717 5674 5783 5677
rect 7782 5674 7788 5676
rect 5349 5616 5354 5672
rect 5349 5612 5396 5616
rect 5460 5614 5506 5674
rect 5717 5672 7788 5674
rect 5717 5616 5722 5672
rect 5778 5616 7788 5672
rect 5717 5614 7788 5616
rect 5460 5612 5466 5614
rect 5349 5611 5415 5612
rect 5717 5611 5783 5614
rect 7782 5612 7788 5614
rect 7852 5612 7858 5676
rect 9121 5674 9187 5677
rect 10225 5674 10291 5677
rect 10961 5674 11027 5677
rect 8158 5614 8816 5674
rect 7782 5538 7788 5540
rect 5214 5478 7788 5538
rect 7782 5476 7788 5478
rect 7852 5476 7858 5540
rect 3409 5472 3729 5473
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 4470 5340 4476 5404
rect 4540 5402 4546 5404
rect 4797 5402 4863 5405
rect 4540 5400 4863 5402
rect 4540 5344 4802 5400
rect 4858 5344 4863 5400
rect 4540 5342 4863 5344
rect 4540 5340 4546 5342
rect 4797 5339 4863 5342
rect 5349 5402 5415 5405
rect 8158 5402 8218 5614
rect 8756 5538 8816 5614
rect 9121 5672 10058 5674
rect 9121 5616 9126 5672
rect 9182 5616 10058 5672
rect 9121 5614 10058 5616
rect 9121 5611 9187 5614
rect 9070 5538 9076 5540
rect 8756 5478 9076 5538
rect 9070 5476 9076 5478
rect 9140 5476 9146 5540
rect 9998 5538 10058 5614
rect 10225 5672 11027 5674
rect 10225 5616 10230 5672
rect 10286 5616 10966 5672
rect 11022 5616 11027 5672
rect 10225 5614 11027 5616
rect 10225 5611 10291 5614
rect 10961 5611 11027 5614
rect 11237 5674 11303 5677
rect 12198 5674 12204 5676
rect 11237 5672 12204 5674
rect 11237 5616 11242 5672
rect 11298 5616 12204 5672
rect 11237 5614 12204 5616
rect 11237 5611 11303 5614
rect 12198 5612 12204 5614
rect 12268 5612 12274 5676
rect 12341 5674 12407 5677
rect 14273 5674 14339 5677
rect 12341 5672 14339 5674
rect 12341 5616 12346 5672
rect 12402 5616 14278 5672
rect 14334 5616 14339 5672
rect 12341 5614 14339 5616
rect 12341 5611 12407 5614
rect 14273 5611 14339 5614
rect 10317 5538 10383 5541
rect 9998 5536 10383 5538
rect 9998 5480 10322 5536
rect 10378 5480 10383 5536
rect 9998 5478 10383 5480
rect 10317 5475 10383 5478
rect 10685 5538 10751 5541
rect 11646 5538 11652 5540
rect 10685 5536 11652 5538
rect 10685 5480 10690 5536
rect 10746 5480 11652 5536
rect 10685 5478 11652 5480
rect 10685 5475 10751 5478
rect 11646 5476 11652 5478
rect 11716 5476 11722 5540
rect 11789 5538 11855 5541
rect 12198 5538 12204 5540
rect 11789 5536 12204 5538
rect 11789 5480 11794 5536
rect 11850 5480 12204 5536
rect 11789 5478 12204 5480
rect 11789 5475 11855 5478
rect 12198 5476 12204 5478
rect 12268 5476 12274 5540
rect 12525 5536 12591 5541
rect 12525 5480 12530 5536
rect 12586 5480 12591 5536
rect 12525 5475 12591 5480
rect 12801 5538 12867 5541
rect 12985 5538 13051 5541
rect 12801 5536 13051 5538
rect 12801 5480 12806 5536
rect 12862 5480 12990 5536
rect 13046 5480 13051 5536
rect 12801 5478 13051 5480
rect 12801 5475 12867 5478
rect 12985 5475 13051 5478
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 5349 5400 8218 5402
rect 5349 5344 5354 5400
rect 5410 5344 8218 5400
rect 5349 5342 8218 5344
rect 5349 5339 5415 5342
rect 9622 5340 9628 5404
rect 9692 5402 9698 5404
rect 12528 5402 12588 5475
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 9692 5342 12588 5402
rect 9692 5340 9698 5342
rect 0 5266 480 5296
rect 841 5266 907 5269
rect 0 5264 907 5266
rect 0 5208 846 5264
rect 902 5208 907 5264
rect 0 5206 907 5208
rect 0 5176 480 5206
rect 841 5203 907 5206
rect 2497 5266 2563 5269
rect 9121 5266 9187 5269
rect 2497 5264 9187 5266
rect 2497 5208 2502 5264
rect 2558 5208 9126 5264
rect 9182 5208 9187 5264
rect 2497 5206 9187 5208
rect 2497 5203 2563 5206
rect 9121 5203 9187 5206
rect 10409 5266 10475 5269
rect 13169 5266 13235 5269
rect 13813 5266 13879 5269
rect 10409 5264 13879 5266
rect 10409 5208 10414 5264
rect 10470 5208 13174 5264
rect 13230 5208 13818 5264
rect 13874 5208 13879 5264
rect 10409 5206 13879 5208
rect 10409 5203 10475 5206
rect 13169 5203 13235 5206
rect 13813 5203 13879 5206
rect 1393 5130 1459 5133
rect 3509 5130 3575 5133
rect 6637 5130 6703 5133
rect 1393 5128 3434 5130
rect 1393 5072 1398 5128
rect 1454 5072 3434 5128
rect 1393 5070 3434 5072
rect 1393 5067 1459 5070
rect 3374 4994 3434 5070
rect 3509 5128 6703 5130
rect 3509 5072 3514 5128
rect 3570 5072 6642 5128
rect 6698 5072 6703 5128
rect 3509 5070 6703 5072
rect 3509 5067 3575 5070
rect 6637 5067 6703 5070
rect 7281 5130 7347 5133
rect 9622 5130 9628 5132
rect 7281 5128 9628 5130
rect 7281 5072 7286 5128
rect 7342 5072 9628 5128
rect 7281 5070 9628 5072
rect 7281 5067 7347 5070
rect 9622 5068 9628 5070
rect 9692 5068 9698 5132
rect 13629 5130 13695 5133
rect 9814 5128 13695 5130
rect 9814 5072 13634 5128
rect 13690 5072 13695 5128
rect 9814 5070 13695 5072
rect 5349 4994 5415 4997
rect 3374 4992 5415 4994
rect 3374 4936 5354 4992
rect 5410 4936 5415 4992
rect 3374 4934 5415 4936
rect 5349 4931 5415 4934
rect 7189 4994 7255 4997
rect 9814 4994 9874 5070
rect 13629 5067 13695 5070
rect 7189 4992 9874 4994
rect 7189 4936 7194 4992
rect 7250 4936 9874 4992
rect 7189 4934 9874 4936
rect 7189 4931 7255 4934
rect 10174 4932 10180 4996
rect 10244 4994 10250 4996
rect 10409 4994 10475 4997
rect 10244 4992 10475 4994
rect 10244 4936 10414 4992
rect 10470 4936 10475 4992
rect 10244 4934 10475 4936
rect 10244 4932 10250 4934
rect 10409 4931 10475 4934
rect 12566 4932 12572 4996
rect 12636 4994 12642 4996
rect 13261 4994 13327 4997
rect 13445 4994 13511 4997
rect 12636 4992 13511 4994
rect 12636 4936 13266 4992
rect 13322 4936 13450 4992
rect 13506 4936 13511 4992
rect 12636 4934 13511 4936
rect 12636 4932 12642 4934
rect 13261 4931 13327 4934
rect 13445 4931 13511 4934
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 1669 4858 1735 4861
rect 10133 4860 10199 4861
rect 5022 4858 5028 4860
rect 1669 4856 5028 4858
rect 1669 4800 1674 4856
rect 1730 4800 5028 4856
rect 1669 4798 5028 4800
rect 1669 4795 1735 4798
rect 5022 4796 5028 4798
rect 5092 4796 5098 4860
rect 9622 4858 9628 4860
rect 6272 4798 9628 4858
rect 4102 4660 4108 4724
rect 4172 4722 4178 4724
rect 6272 4722 6332 4798
rect 9622 4796 9628 4798
rect 9692 4796 9698 4860
rect 10133 4856 10180 4860
rect 10244 4858 10250 4860
rect 11237 4858 11303 4861
rect 13353 4858 13419 4861
rect 10133 4800 10138 4856
rect 10133 4796 10180 4800
rect 10244 4798 10290 4858
rect 11237 4856 13419 4858
rect 11237 4800 11242 4856
rect 11298 4800 13358 4856
rect 13414 4800 13419 4856
rect 11237 4798 13419 4800
rect 10244 4796 10250 4798
rect 10133 4795 10199 4796
rect 11237 4795 11303 4798
rect 13353 4795 13419 4798
rect 4172 4662 6332 4722
rect 4172 4660 4178 4662
rect 7414 4660 7420 4724
rect 7484 4722 7490 4724
rect 11973 4722 12039 4725
rect 7484 4720 12039 4722
rect 7484 4664 11978 4720
rect 12034 4664 12039 4720
rect 7484 4662 12039 4664
rect 7484 4660 7490 4662
rect 11973 4659 12039 4662
rect 12341 4722 12407 4725
rect 12801 4722 12867 4725
rect 12341 4720 12867 4722
rect 12341 4664 12346 4720
rect 12402 4664 12806 4720
rect 12862 4664 12867 4720
rect 12341 4662 12867 4664
rect 12341 4659 12407 4662
rect 12801 4659 12867 4662
rect 12934 4660 12940 4724
rect 13004 4722 13010 4724
rect 13721 4722 13787 4725
rect 13004 4720 13787 4722
rect 13004 4664 13726 4720
rect 13782 4664 13787 4720
rect 13004 4662 13787 4664
rect 13004 4660 13010 4662
rect 13721 4659 13787 4662
rect 2865 4586 2931 4589
rect 12433 4586 12499 4589
rect 14222 4586 14228 4588
rect 2865 4584 12499 4586
rect 2865 4528 2870 4584
rect 2926 4528 12438 4584
rect 12494 4528 12499 4584
rect 2865 4526 12499 4528
rect 2865 4523 2931 4526
rect 12433 4523 12499 4526
rect 12988 4526 14228 4586
rect 4705 4450 4771 4453
rect 6821 4450 6887 4453
rect 4705 4448 6887 4450
rect 4705 4392 4710 4448
rect 4766 4392 6826 4448
rect 6882 4392 6887 4448
rect 4705 4390 6887 4392
rect 4705 4387 4771 4390
rect 6821 4387 6887 4390
rect 7005 4450 7071 4453
rect 8753 4450 8819 4453
rect 9029 4450 9095 4453
rect 9254 4450 9260 4452
rect 7005 4448 8172 4450
rect 7005 4392 7010 4448
rect 7066 4392 8172 4448
rect 7005 4390 8172 4392
rect 7005 4387 7071 4390
rect 3409 4384 3729 4385
rect 0 4314 480 4344
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 2865 4314 2931 4317
rect 0 4312 2931 4314
rect 0 4256 2870 4312
rect 2926 4256 2931 4312
rect 0 4254 2931 4256
rect 0 4224 480 4254
rect 2865 4251 2931 4254
rect 4153 4314 4219 4317
rect 4797 4316 4863 4317
rect 4470 4314 4476 4316
rect 4153 4312 4476 4314
rect 4153 4256 4158 4312
rect 4214 4256 4476 4312
rect 4153 4254 4476 4256
rect 4153 4251 4219 4254
rect 4470 4252 4476 4254
rect 4540 4252 4546 4316
rect 4797 4314 4844 4316
rect 4752 4312 4844 4314
rect 4752 4256 4802 4312
rect 4752 4254 4844 4256
rect 4797 4252 4844 4254
rect 4908 4252 4914 4316
rect 4981 4314 5047 4317
rect 7649 4314 7715 4317
rect 4981 4312 7715 4314
rect 4981 4256 4986 4312
rect 5042 4256 7654 4312
rect 7710 4256 7715 4312
rect 4981 4254 7715 4256
rect 4797 4251 4863 4252
rect 4981 4251 5047 4254
rect 7649 4251 7715 4254
rect 7782 4252 7788 4316
rect 7852 4314 7858 4316
rect 7852 4254 8034 4314
rect 7852 4252 7858 4254
rect 1853 4178 1919 4181
rect 3509 4178 3575 4181
rect 1853 4176 3575 4178
rect 1853 4120 1858 4176
rect 1914 4120 3514 4176
rect 3570 4120 3575 4176
rect 1853 4118 3575 4120
rect 1853 4115 1919 4118
rect 3509 4115 3575 4118
rect 3693 4178 3759 4181
rect 7782 4178 7788 4180
rect 3693 4176 7788 4178
rect 3693 4120 3698 4176
rect 3754 4120 7788 4176
rect 3693 4118 7788 4120
rect 3693 4115 3759 4118
rect 7782 4116 7788 4118
rect 7852 4116 7858 4180
rect 1669 4042 1735 4045
rect 4153 4042 4219 4045
rect 1669 4040 4219 4042
rect 1669 3984 1674 4040
rect 1730 3984 4158 4040
rect 4214 3984 4219 4040
rect 1669 3982 4219 3984
rect 1669 3979 1735 3982
rect 4153 3979 4219 3982
rect 4286 3980 4292 4044
rect 4356 4042 4362 4044
rect 6269 4042 6335 4045
rect 4356 4040 6335 4042
rect 4356 3984 6274 4040
rect 6330 3984 6335 4040
rect 4356 3982 6335 3984
rect 4356 3980 4362 3982
rect 6269 3979 6335 3982
rect 6545 4042 6611 4045
rect 7046 4042 7052 4044
rect 6545 4040 7052 4042
rect 6545 3984 6550 4040
rect 6606 3984 7052 4040
rect 6545 3982 7052 3984
rect 6545 3979 6611 3982
rect 7046 3980 7052 3982
rect 7116 3980 7122 4044
rect 7230 3980 7236 4044
rect 7300 4042 7306 4044
rect 7557 4042 7623 4045
rect 7300 4040 7623 4042
rect 7300 3984 7562 4040
rect 7618 3984 7623 4040
rect 7300 3982 7623 3984
rect 7974 4042 8034 4254
rect 8112 4178 8172 4390
rect 8753 4448 9260 4450
rect 8753 4392 8758 4448
rect 8814 4392 9034 4448
rect 9090 4392 9260 4448
rect 8753 4390 9260 4392
rect 8753 4387 8819 4390
rect 9029 4387 9095 4390
rect 9254 4388 9260 4390
rect 9324 4388 9330 4452
rect 9673 4450 9739 4453
rect 9673 4448 12818 4450
rect 9673 4392 9678 4448
rect 9734 4392 12818 4448
rect 9673 4390 12818 4392
rect 9673 4387 9739 4390
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 8753 4314 8819 4317
rect 9070 4314 9076 4316
rect 8753 4312 9076 4314
rect 8753 4256 8758 4312
rect 8814 4256 9076 4312
rect 8753 4254 9076 4256
rect 8753 4251 8819 4254
rect 9070 4252 9076 4254
rect 9140 4252 9146 4316
rect 9673 4314 9739 4317
rect 11053 4314 11119 4317
rect 9673 4312 11119 4314
rect 9673 4256 9678 4312
rect 9734 4256 11058 4312
rect 11114 4256 11119 4312
rect 9673 4254 11119 4256
rect 9673 4251 9739 4254
rect 11053 4251 11119 4254
rect 11513 4314 11579 4317
rect 11697 4314 11763 4317
rect 11513 4312 11763 4314
rect 11513 4256 11518 4312
rect 11574 4256 11702 4312
rect 11758 4256 11763 4312
rect 11513 4254 11763 4256
rect 11513 4251 11579 4254
rect 11697 4251 11763 4254
rect 12014 4252 12020 4316
rect 12084 4314 12090 4316
rect 12617 4314 12683 4317
rect 12084 4312 12683 4314
rect 12084 4256 12622 4312
rect 12678 4256 12683 4312
rect 12084 4254 12683 4256
rect 12084 4252 12090 4254
rect 12617 4251 12683 4254
rect 8293 4178 8359 4181
rect 8112 4176 8359 4178
rect 8112 4120 8298 4176
rect 8354 4120 8359 4176
rect 8112 4118 8359 4120
rect 8293 4115 8359 4118
rect 8569 4178 8635 4181
rect 9489 4178 9555 4181
rect 10409 4180 10475 4181
rect 8569 4176 9555 4178
rect 8569 4120 8574 4176
rect 8630 4120 9494 4176
rect 9550 4120 9555 4176
rect 8569 4118 9555 4120
rect 8569 4115 8635 4118
rect 9489 4115 9555 4118
rect 10358 4116 10364 4180
rect 10428 4178 10475 4180
rect 10869 4178 10935 4181
rect 12525 4178 12591 4181
rect 10428 4176 10520 4178
rect 10470 4120 10520 4176
rect 10428 4118 10520 4120
rect 10869 4176 12591 4178
rect 10869 4120 10874 4176
rect 10930 4120 12530 4176
rect 12586 4120 12591 4176
rect 10869 4118 12591 4120
rect 10428 4116 10475 4118
rect 10409 4115 10475 4116
rect 10869 4115 10935 4118
rect 12525 4115 12591 4118
rect 8477 4042 8543 4045
rect 11462 4042 11468 4044
rect 7974 4040 11468 4042
rect 7974 3984 8482 4040
rect 8538 3984 11468 4040
rect 7974 3982 11468 3984
rect 7300 3980 7306 3982
rect 7557 3979 7623 3982
rect 8477 3979 8543 3982
rect 11462 3980 11468 3982
rect 11532 4042 11538 4044
rect 12065 4042 12131 4045
rect 11532 4040 12131 4042
rect 11532 3984 12070 4040
rect 12126 3984 12131 4040
rect 11532 3982 12131 3984
rect 12758 4042 12818 4390
rect 12988 4181 13048 4526
rect 14222 4524 14228 4526
rect 14292 4524 14298 4588
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 4319 13590 4320
rect 12985 4176 13051 4181
rect 12985 4120 12990 4176
rect 13046 4120 13051 4176
rect 12985 4115 13051 4120
rect 13261 4042 13327 4045
rect 12758 4040 13327 4042
rect 12758 3984 13266 4040
rect 13322 3984 13327 4040
rect 12758 3982 13327 3984
rect 11532 3980 11538 3982
rect 12065 3979 12131 3982
rect 13261 3979 13327 3982
rect 1853 3906 1919 3909
rect 5574 3906 5580 3908
rect 1853 3904 5580 3906
rect 1853 3848 1858 3904
rect 1914 3848 5580 3904
rect 1853 3846 5580 3848
rect 1853 3843 1919 3846
rect 5574 3844 5580 3846
rect 5644 3844 5650 3908
rect 6729 3906 6795 3909
rect 10133 3906 10199 3909
rect 6729 3904 10199 3906
rect 6729 3848 6734 3904
rect 6790 3848 10138 3904
rect 10194 3848 10199 3904
rect 6729 3846 10199 3848
rect 6729 3843 6795 3846
rect 10133 3843 10199 3846
rect 11462 3844 11468 3908
rect 11532 3906 11538 3908
rect 11697 3906 11763 3909
rect 11532 3904 11763 3906
rect 11532 3848 11702 3904
rect 11758 3848 11763 3904
rect 11532 3846 11763 3848
rect 11532 3844 11538 3846
rect 11697 3843 11763 3846
rect 12014 3844 12020 3908
rect 12084 3906 12090 3908
rect 15009 3906 15075 3909
rect 12084 3904 15075 3906
rect 12084 3848 15014 3904
rect 15070 3848 15075 3904
rect 12084 3846 15075 3848
rect 12084 3844 12090 3846
rect 15009 3843 15075 3846
rect 5874 3840 6194 3841
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 3233 3770 3299 3773
rect 5574 3770 5580 3772
rect 3233 3768 5580 3770
rect 3233 3712 3238 3768
rect 3294 3712 5580 3768
rect 3233 3710 5580 3712
rect 3233 3707 3299 3710
rect 5574 3708 5580 3710
rect 5644 3708 5650 3772
rect 9806 3708 9812 3772
rect 9876 3770 9882 3772
rect 9949 3770 10015 3773
rect 9876 3768 10015 3770
rect 9876 3712 9954 3768
rect 10010 3712 10015 3768
rect 9876 3710 10015 3712
rect 9876 3708 9882 3710
rect 9949 3707 10015 3710
rect 12198 3708 12204 3772
rect 12268 3770 12274 3772
rect 13629 3770 13695 3773
rect 12268 3768 13695 3770
rect 12268 3712 13634 3768
rect 13690 3712 13695 3768
rect 12268 3710 13695 3712
rect 12268 3708 12274 3710
rect 13629 3707 13695 3710
rect 3182 3572 3188 3636
rect 3252 3634 3258 3636
rect 3509 3634 3575 3637
rect 3252 3632 3575 3634
rect 3252 3576 3514 3632
rect 3570 3576 3575 3632
rect 3252 3574 3575 3576
rect 3252 3572 3258 3574
rect 3509 3571 3575 3574
rect 3918 3572 3924 3636
rect 3988 3634 3994 3636
rect 9305 3634 9371 3637
rect 12566 3634 12572 3636
rect 3988 3574 9138 3634
rect 3988 3572 3994 3574
rect 3233 3500 3299 3501
rect 3182 3498 3188 3500
rect 3142 3438 3188 3498
rect 3252 3496 3299 3500
rect 3294 3440 3299 3496
rect 3182 3436 3188 3438
rect 3252 3436 3299 3440
rect 3233 3435 3299 3436
rect 3417 3498 3483 3501
rect 4521 3498 4587 3501
rect 5022 3498 5028 3500
rect 3417 3496 3986 3498
rect 3417 3440 3422 3496
rect 3478 3440 3986 3496
rect 3417 3438 3986 3440
rect 3417 3435 3483 3438
rect 0 3362 480 3392
rect 1669 3362 1735 3365
rect 0 3360 1735 3362
rect 0 3304 1674 3360
rect 1730 3304 1735 3360
rect 0 3302 1735 3304
rect 3926 3362 3986 3438
rect 4521 3496 5028 3498
rect 4521 3440 4526 3496
rect 4582 3440 5028 3496
rect 4521 3438 5028 3440
rect 4521 3435 4587 3438
rect 5022 3436 5028 3438
rect 5092 3436 5098 3500
rect 5349 3498 5415 3501
rect 9078 3498 9138 3574
rect 9305 3632 12572 3634
rect 9305 3576 9310 3632
rect 9366 3576 12572 3632
rect 9305 3574 12572 3576
rect 9305 3571 9371 3574
rect 12566 3572 12572 3574
rect 12636 3572 12642 3636
rect 12893 3634 12959 3637
rect 13118 3634 13124 3636
rect 12893 3632 13124 3634
rect 12893 3576 12898 3632
rect 12954 3576 13124 3632
rect 12893 3574 13124 3576
rect 12893 3571 12959 3574
rect 13118 3572 13124 3574
rect 13188 3572 13194 3636
rect 12157 3498 12223 3501
rect 14549 3498 14615 3501
rect 5349 3496 9000 3498
rect 5349 3440 5354 3496
rect 5410 3440 9000 3496
rect 5349 3438 9000 3440
rect 9078 3496 12223 3498
rect 9078 3440 12162 3496
rect 12218 3440 12223 3496
rect 9078 3438 12223 3440
rect 5349 3435 5415 3438
rect 6729 3362 6795 3365
rect 3926 3360 6795 3362
rect 3926 3304 6734 3360
rect 6790 3304 6795 3360
rect 3926 3302 6795 3304
rect 8940 3362 9000 3438
rect 12157 3435 12223 3438
rect 12344 3496 14615 3498
rect 12344 3440 14554 3496
rect 14610 3440 14615 3496
rect 12344 3438 14615 3440
rect 12344 3362 12404 3438
rect 14549 3435 14615 3438
rect 8940 3302 12404 3362
rect 12801 3362 12867 3365
rect 13077 3362 13143 3365
rect 12801 3360 13143 3362
rect 12801 3304 12806 3360
rect 12862 3304 13082 3360
rect 13138 3304 13143 3360
rect 12801 3302 13143 3304
rect 0 3272 480 3302
rect 1669 3299 1735 3302
rect 6729 3299 6795 3302
rect 12801 3299 12867 3302
rect 13077 3299 13143 3302
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 3231 13590 3232
rect 3877 3228 3943 3229
rect 3877 3226 3924 3228
rect 3832 3224 3924 3226
rect 3832 3168 3882 3224
rect 3832 3166 3924 3168
rect 3877 3164 3924 3166
rect 3988 3164 3994 3228
rect 4245 3226 4311 3229
rect 5349 3226 5415 3229
rect 4245 3224 5415 3226
rect 4245 3168 4250 3224
rect 4306 3168 5354 3224
rect 5410 3168 5415 3224
rect 4245 3166 5415 3168
rect 3877 3163 3943 3164
rect 4245 3163 4311 3166
rect 5349 3163 5415 3166
rect 5574 3164 5580 3228
rect 5644 3226 5650 3228
rect 8109 3226 8175 3229
rect 5644 3224 8175 3226
rect 5644 3168 8114 3224
rect 8170 3168 8175 3224
rect 5644 3166 8175 3168
rect 5644 3164 5650 3166
rect 8109 3163 8175 3166
rect 9070 3164 9076 3228
rect 9140 3226 9146 3228
rect 11278 3226 11284 3228
rect 9140 3166 11284 3226
rect 9140 3164 9146 3166
rect 11278 3164 11284 3166
rect 11348 3164 11354 3228
rect 11462 3164 11468 3228
rect 11532 3226 11538 3228
rect 11973 3226 12039 3229
rect 11532 3224 12039 3226
rect 11532 3168 11978 3224
rect 12034 3168 12039 3224
rect 11532 3166 12039 3168
rect 11532 3164 11538 3166
rect 11973 3163 12039 3166
rect 12382 3164 12388 3228
rect 12452 3226 12458 3228
rect 13077 3226 13143 3229
rect 12452 3224 13143 3226
rect 12452 3168 13082 3224
rect 13138 3168 13143 3224
rect 12452 3166 13143 3168
rect 12452 3164 12458 3166
rect 13077 3163 13143 3166
rect 13813 3226 13879 3229
rect 14406 3226 14412 3228
rect 13813 3224 14412 3226
rect 13813 3168 13818 3224
rect 13874 3168 14412 3224
rect 13813 3166 14412 3168
rect 13813 3163 13879 3166
rect 14406 3164 14412 3166
rect 14476 3164 14482 3228
rect 3509 3090 3575 3093
rect 12014 3090 12020 3092
rect 3509 3088 12020 3090
rect 3509 3032 3514 3088
rect 3570 3032 12020 3088
rect 3509 3030 12020 3032
rect 3509 3027 3575 3030
rect 12014 3028 12020 3030
rect 12084 3028 12090 3092
rect 12157 3090 12223 3093
rect 14181 3090 14247 3093
rect 12157 3088 14247 3090
rect 12157 3032 12162 3088
rect 12218 3032 14186 3088
rect 14242 3032 14247 3088
rect 12157 3030 14247 3032
rect 12157 3027 12223 3030
rect 14181 3027 14247 3030
rect 2681 2954 2747 2957
rect 13721 2954 13787 2957
rect 2681 2952 13787 2954
rect 2681 2896 2686 2952
rect 2742 2896 13726 2952
rect 13782 2896 13787 2952
rect 2681 2894 13787 2896
rect 2681 2891 2747 2894
rect 13721 2891 13787 2894
rect 3049 2818 3115 2821
rect 3417 2818 3483 2821
rect 3969 2820 4035 2821
rect 3918 2818 3924 2820
rect 3049 2816 3483 2818
rect 3049 2760 3054 2816
rect 3110 2760 3422 2816
rect 3478 2760 3483 2816
rect 3049 2758 3483 2760
rect 3878 2758 3924 2818
rect 3988 2816 4035 2820
rect 4030 2760 4035 2816
rect 3049 2755 3115 2758
rect 3417 2755 3483 2758
rect 3918 2756 3924 2758
rect 3988 2756 4035 2760
rect 4470 2756 4476 2820
rect 4540 2818 4546 2820
rect 5441 2818 5507 2821
rect 4540 2816 5507 2818
rect 4540 2760 5446 2816
rect 5502 2760 5507 2816
rect 4540 2758 5507 2760
rect 4540 2756 4546 2758
rect 3969 2755 4035 2756
rect 5441 2755 5507 2758
rect 6729 2818 6795 2821
rect 8886 2818 8892 2820
rect 6729 2816 8892 2818
rect 6729 2760 6734 2816
rect 6790 2760 8892 2816
rect 6729 2758 8892 2760
rect 6729 2755 6795 2758
rect 8886 2756 8892 2758
rect 8956 2756 8962 2820
rect 9622 2756 9628 2820
rect 9692 2818 9698 2820
rect 10409 2818 10475 2821
rect 10593 2820 10659 2821
rect 9692 2816 10475 2818
rect 9692 2760 10414 2816
rect 10470 2760 10475 2816
rect 9692 2758 10475 2760
rect 9692 2756 9698 2758
rect 10409 2755 10475 2758
rect 10542 2756 10548 2820
rect 10612 2818 10659 2820
rect 10612 2816 10704 2818
rect 10654 2760 10704 2816
rect 10612 2758 10704 2760
rect 10612 2756 10659 2758
rect 11462 2756 11468 2820
rect 11532 2818 11538 2820
rect 11605 2818 11671 2821
rect 11789 2820 11855 2821
rect 11789 2818 11836 2820
rect 11532 2816 11671 2818
rect 11532 2760 11610 2816
rect 11666 2760 11671 2816
rect 11532 2758 11671 2760
rect 11744 2816 11836 2818
rect 11744 2760 11794 2816
rect 11744 2758 11836 2760
rect 11532 2756 11538 2758
rect 10593 2755 10659 2756
rect 11605 2755 11671 2758
rect 11789 2756 11836 2758
rect 11900 2756 11906 2820
rect 13721 2818 13787 2821
rect 15009 2818 15075 2821
rect 13721 2816 15075 2818
rect 13721 2760 13726 2816
rect 13782 2760 15014 2816
rect 15070 2760 15075 2816
rect 13721 2758 15075 2760
rect 11789 2755 11855 2756
rect 13721 2755 13787 2758
rect 15009 2755 15075 2758
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 3141 2682 3207 2685
rect 4654 2682 4660 2684
rect 3141 2680 4660 2682
rect 3141 2624 3146 2680
rect 3202 2624 4660 2680
rect 3141 2622 4660 2624
rect 3141 2619 3207 2622
rect 4654 2620 4660 2622
rect 4724 2620 4730 2684
rect 5206 2620 5212 2684
rect 5276 2682 5282 2684
rect 5625 2682 5691 2685
rect 5276 2680 5691 2682
rect 5276 2624 5630 2680
rect 5686 2624 5691 2680
rect 5276 2622 5691 2624
rect 5276 2620 5282 2622
rect 5625 2619 5691 2622
rect 6678 2620 6684 2684
rect 6748 2682 6754 2684
rect 6821 2682 6887 2685
rect 6748 2680 6887 2682
rect 6748 2624 6826 2680
rect 6882 2624 6887 2680
rect 6748 2622 6887 2624
rect 6748 2620 6754 2622
rect 6821 2619 6887 2622
rect 8017 2682 8083 2685
rect 8150 2682 8156 2684
rect 8017 2680 8156 2682
rect 8017 2624 8022 2680
rect 8078 2624 8156 2680
rect 8017 2622 8156 2624
rect 8017 2619 8083 2622
rect 8150 2620 8156 2622
rect 8220 2620 8226 2684
rect 9305 2682 9371 2685
rect 8342 2680 9371 2682
rect 8342 2624 9310 2680
rect 9366 2624 9371 2680
rect 8342 2622 9371 2624
rect 1301 2546 1367 2549
rect 4613 2546 4679 2549
rect 7465 2546 7531 2549
rect 8342 2546 8402 2622
rect 9305 2619 9371 2622
rect 10174 2620 10180 2684
rect 10244 2682 10250 2684
rect 10317 2682 10383 2685
rect 12157 2682 12223 2685
rect 10244 2680 10383 2682
rect 10244 2624 10322 2680
rect 10378 2624 10383 2680
rect 10244 2622 10383 2624
rect 10244 2620 10250 2622
rect 10317 2619 10383 2622
rect 11332 2680 12223 2682
rect 11332 2624 12162 2680
rect 12218 2624 12223 2680
rect 11332 2622 12223 2624
rect 1301 2544 8402 2546
rect 1301 2488 1306 2544
rect 1362 2488 4618 2544
rect 4674 2488 7470 2544
rect 7526 2488 8402 2544
rect 1301 2486 8402 2488
rect 8845 2546 8911 2549
rect 11332 2546 11392 2622
rect 12157 2619 12223 2622
rect 12617 2682 12683 2685
rect 13997 2684 14063 2685
rect 12750 2682 12756 2684
rect 12617 2680 12756 2682
rect 12617 2624 12622 2680
rect 12678 2624 12756 2680
rect 12617 2622 12756 2624
rect 12617 2619 12683 2622
rect 12750 2620 12756 2622
rect 12820 2620 12826 2684
rect 13997 2682 14044 2684
rect 13952 2680 14044 2682
rect 13952 2624 14002 2680
rect 13952 2622 14044 2624
rect 13997 2620 14044 2622
rect 14108 2620 14114 2684
rect 13997 2619 14063 2620
rect 8845 2544 11392 2546
rect 8845 2488 8850 2544
rect 8906 2488 11392 2544
rect 8845 2486 11392 2488
rect 11513 2546 11579 2549
rect 13813 2546 13879 2549
rect 11513 2544 13879 2546
rect 11513 2488 11518 2544
rect 11574 2488 13818 2544
rect 13874 2488 13879 2544
rect 11513 2486 13879 2488
rect 1301 2483 1367 2486
rect 4613 2483 4679 2486
rect 7465 2483 7531 2486
rect 8845 2483 8911 2486
rect 11513 2483 11579 2486
rect 13813 2483 13879 2486
rect 0 2410 480 2440
rect 5349 2410 5415 2413
rect 6862 2410 6868 2412
rect 0 2408 6868 2410
rect 0 2352 5354 2408
rect 5410 2352 6868 2408
rect 0 2350 6868 2352
rect 0 2320 480 2350
rect 5349 2347 5415 2350
rect 6862 2348 6868 2350
rect 6932 2348 6938 2412
rect 7557 2410 7623 2413
rect 12525 2410 12591 2413
rect 7557 2408 12591 2410
rect 7557 2352 7562 2408
rect 7618 2352 12530 2408
rect 12586 2352 12591 2408
rect 7557 2350 12591 2352
rect 7557 2347 7623 2350
rect 12525 2347 12591 2350
rect 4337 2274 4403 2277
rect 7598 2274 7604 2276
rect 4337 2272 7604 2274
rect 4337 2216 4342 2272
rect 4398 2216 7604 2272
rect 4337 2214 7604 2216
rect 4337 2211 4403 2214
rect 7598 2212 7604 2214
rect 7668 2212 7674 2276
rect 7782 2212 7788 2276
rect 7852 2274 7858 2276
rect 7925 2274 7991 2277
rect 7852 2272 7991 2274
rect 7852 2216 7930 2272
rect 7986 2216 7991 2272
rect 7852 2214 7991 2216
rect 7852 2212 7858 2214
rect 7925 2211 7991 2214
rect 9254 2212 9260 2276
rect 9324 2274 9330 2276
rect 11329 2274 11395 2277
rect 9324 2272 11395 2274
rect 9324 2216 11334 2272
rect 11390 2216 11395 2272
rect 9324 2214 11395 2216
rect 9324 2212 9330 2214
rect 11329 2211 11395 2214
rect 11462 2212 11468 2276
rect 11532 2274 11538 2276
rect 12801 2274 12867 2277
rect 13813 2276 13879 2277
rect 13813 2274 13860 2276
rect 11532 2272 12867 2274
rect 11532 2216 12806 2272
rect 12862 2216 12867 2272
rect 11532 2214 12867 2216
rect 13768 2272 13860 2274
rect 13768 2216 13818 2272
rect 13768 2214 13860 2216
rect 11532 2212 11538 2214
rect 12801 2211 12867 2214
rect 13813 2212 13860 2214
rect 13924 2212 13930 2276
rect 13813 2211 13879 2212
rect 3409 2208 3729 2209
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
rect 8753 2138 8819 2141
rect 12198 2138 12204 2140
rect 8753 2136 12204 2138
rect 8753 2080 8758 2136
rect 8814 2080 12204 2136
rect 8753 2078 12204 2080
rect 8753 2075 8819 2078
rect 12198 2076 12204 2078
rect 12268 2076 12274 2140
rect 1853 2002 1919 2005
rect 14089 2002 14155 2005
rect 1853 2000 14155 2002
rect 1853 1944 1858 2000
rect 1914 1944 14094 2000
rect 14150 1944 14155 2000
rect 1853 1942 14155 1944
rect 1853 1939 1919 1942
rect 14089 1939 14155 1942
rect 15561 2002 15627 2005
rect 16520 2002 17000 2032
rect 15561 2000 17000 2002
rect 15561 1944 15566 2000
rect 15622 1944 17000 2000
rect 15561 1942 17000 1944
rect 15561 1939 15627 1942
rect 16520 1912 17000 1942
rect 3918 1804 3924 1868
rect 3988 1866 3994 1868
rect 11513 1866 11579 1869
rect 3988 1864 11579 1866
rect 3988 1808 11518 1864
rect 11574 1808 11579 1864
rect 3988 1806 11579 1808
rect 3988 1804 3994 1806
rect 11513 1803 11579 1806
rect 3509 1730 3575 1733
rect 4102 1730 4108 1732
rect 3509 1728 4108 1730
rect 3509 1672 3514 1728
rect 3570 1672 4108 1728
rect 3509 1670 4108 1672
rect 3509 1667 3575 1670
rect 4102 1668 4108 1670
rect 4172 1668 4178 1732
rect 5390 1668 5396 1732
rect 5460 1730 5466 1732
rect 14273 1730 14339 1733
rect 5460 1728 14339 1730
rect 5460 1672 14278 1728
rect 14334 1672 14339 1728
rect 5460 1670 14339 1672
rect 5460 1668 5466 1670
rect 14273 1667 14339 1670
rect 4981 1594 5047 1597
rect 8937 1594 9003 1597
rect 4981 1592 9003 1594
rect 4981 1536 4986 1592
rect 5042 1536 8942 1592
rect 8998 1536 9003 1592
rect 4981 1534 9003 1536
rect 4981 1531 5047 1534
rect 8937 1531 9003 1534
rect 11646 1532 11652 1596
rect 11716 1594 11722 1596
rect 14273 1594 14339 1597
rect 11716 1592 14339 1594
rect 11716 1536 14278 1592
rect 14334 1536 14339 1592
rect 11716 1534 14339 1536
rect 11716 1532 11722 1534
rect 14273 1531 14339 1534
rect 0 1458 480 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 480 1398
rect 2773 1395 2839 1398
rect 3182 1396 3188 1460
rect 3252 1458 3258 1460
rect 9070 1458 9076 1460
rect 3252 1398 9076 1458
rect 3252 1396 3258 1398
rect 9070 1396 9076 1398
rect 9140 1396 9146 1460
rect 10358 1396 10364 1460
rect 10428 1458 10434 1460
rect 15101 1458 15167 1461
rect 10428 1456 15167 1458
rect 10428 1400 15106 1456
rect 15162 1400 15167 1456
rect 10428 1398 15167 1400
rect 10428 1396 10434 1398
rect 15101 1395 15167 1398
rect 2221 1322 2287 1325
rect 7414 1322 7420 1324
rect 2221 1320 7420 1322
rect 2221 1264 2226 1320
rect 2282 1264 7420 1320
rect 2221 1262 7420 1264
rect 2221 1259 2287 1262
rect 7414 1260 7420 1262
rect 7484 1260 7490 1324
rect 9397 1322 9463 1325
rect 12934 1322 12940 1324
rect 9397 1320 12940 1322
rect 9397 1264 9402 1320
rect 9458 1264 12940 1320
rect 9397 1262 12940 1264
rect 9397 1259 9463 1262
rect 12934 1260 12940 1262
rect 13004 1260 13010 1324
rect 5533 1186 5599 1189
rect 6310 1186 6316 1188
rect 5533 1184 6316 1186
rect 5533 1128 5538 1184
rect 5594 1128 6316 1184
rect 5533 1126 6316 1128
rect 5533 1123 5599 1126
rect 6310 1124 6316 1126
rect 6380 1124 6386 1188
rect 7966 1124 7972 1188
rect 8036 1186 8042 1188
rect 9673 1186 9739 1189
rect 12893 1186 12959 1189
rect 13670 1186 13676 1188
rect 8036 1184 13676 1186
rect 8036 1128 9678 1184
rect 9734 1128 12898 1184
rect 12954 1128 13676 1184
rect 8036 1126 13676 1128
rect 8036 1124 8042 1126
rect 9673 1123 9739 1126
rect 12893 1123 12959 1126
rect 13670 1124 13676 1126
rect 13740 1124 13746 1188
rect 6177 1050 6243 1053
rect 9990 1050 9996 1052
rect 6177 1048 9996 1050
rect 6177 992 6182 1048
rect 6238 992 9996 1048
rect 6177 990 9996 992
rect 6177 987 6243 990
rect 9990 988 9996 990
rect 10060 1050 10066 1052
rect 10133 1050 10199 1053
rect 10060 1048 10199 1050
rect 10060 992 10138 1048
rect 10194 992 10199 1048
rect 10060 990 10199 992
rect 10060 988 10066 990
rect 10133 987 10199 990
rect 0 506 480 536
rect 1117 506 1183 509
rect 0 504 1183 506
rect 0 448 1122 504
rect 1178 448 1183 504
rect 0 446 1183 448
rect 0 416 480 446
rect 1117 443 1183 446
<< via3 >>
rect 8892 17716 8956 17780
rect 8156 17580 8220 17644
rect 10364 17444 10428 17508
rect 3417 17436 3481 17440
rect 3417 17380 3421 17436
rect 3421 17380 3477 17436
rect 3477 17380 3481 17436
rect 3417 17376 3481 17380
rect 3497 17436 3561 17440
rect 3497 17380 3501 17436
rect 3501 17380 3557 17436
rect 3557 17380 3561 17436
rect 3497 17376 3561 17380
rect 3577 17436 3641 17440
rect 3577 17380 3581 17436
rect 3581 17380 3637 17436
rect 3637 17380 3641 17436
rect 3577 17376 3641 17380
rect 3657 17436 3721 17440
rect 3657 17380 3661 17436
rect 3661 17380 3717 17436
rect 3717 17380 3721 17436
rect 3657 17376 3721 17380
rect 8348 17436 8412 17440
rect 8348 17380 8352 17436
rect 8352 17380 8408 17436
rect 8408 17380 8412 17436
rect 8348 17376 8412 17380
rect 8428 17436 8492 17440
rect 8428 17380 8432 17436
rect 8432 17380 8488 17436
rect 8488 17380 8492 17436
rect 8428 17376 8492 17380
rect 8508 17436 8572 17440
rect 8508 17380 8512 17436
rect 8512 17380 8568 17436
rect 8568 17380 8572 17436
rect 8508 17376 8572 17380
rect 8588 17436 8652 17440
rect 8588 17380 8592 17436
rect 8592 17380 8648 17436
rect 8648 17380 8652 17436
rect 8588 17376 8652 17380
rect 13278 17436 13342 17440
rect 13278 17380 13282 17436
rect 13282 17380 13338 17436
rect 13338 17380 13342 17436
rect 13278 17376 13342 17380
rect 13358 17436 13422 17440
rect 13358 17380 13362 17436
rect 13362 17380 13418 17436
rect 13418 17380 13422 17436
rect 13358 17376 13422 17380
rect 13438 17436 13502 17440
rect 13438 17380 13442 17436
rect 13442 17380 13498 17436
rect 13498 17380 13502 17436
rect 13438 17376 13502 17380
rect 13518 17436 13582 17440
rect 13518 17380 13522 17436
rect 13522 17380 13578 17436
rect 13578 17380 13582 17436
rect 13518 17376 13582 17380
rect 7972 17172 8036 17236
rect 10548 16900 10612 16964
rect 5882 16892 5946 16896
rect 5882 16836 5886 16892
rect 5886 16836 5942 16892
rect 5942 16836 5946 16892
rect 5882 16832 5946 16836
rect 5962 16892 6026 16896
rect 5962 16836 5966 16892
rect 5966 16836 6022 16892
rect 6022 16836 6026 16892
rect 5962 16832 6026 16836
rect 6042 16892 6106 16896
rect 6042 16836 6046 16892
rect 6046 16836 6102 16892
rect 6102 16836 6106 16892
rect 6042 16832 6106 16836
rect 6122 16892 6186 16896
rect 6122 16836 6126 16892
rect 6126 16836 6182 16892
rect 6182 16836 6186 16892
rect 6122 16832 6186 16836
rect 10813 16892 10877 16896
rect 10813 16836 10817 16892
rect 10817 16836 10873 16892
rect 10873 16836 10877 16892
rect 10813 16832 10877 16836
rect 10893 16892 10957 16896
rect 10893 16836 10897 16892
rect 10897 16836 10953 16892
rect 10953 16836 10957 16892
rect 10893 16832 10957 16836
rect 10973 16892 11037 16896
rect 10973 16836 10977 16892
rect 10977 16836 11033 16892
rect 11033 16836 11037 16892
rect 10973 16832 11037 16836
rect 11053 16892 11117 16896
rect 11053 16836 11057 16892
rect 11057 16836 11113 16892
rect 11113 16836 11117 16892
rect 11053 16832 11117 16836
rect 10180 16764 10244 16828
rect 9812 16688 9876 16692
rect 9812 16632 9826 16688
rect 9826 16632 9876 16688
rect 9812 16628 9876 16632
rect 9628 16492 9692 16556
rect 3417 16348 3481 16352
rect 3417 16292 3421 16348
rect 3421 16292 3477 16348
rect 3477 16292 3481 16348
rect 3417 16288 3481 16292
rect 3497 16348 3561 16352
rect 3497 16292 3501 16348
rect 3501 16292 3557 16348
rect 3557 16292 3561 16348
rect 3497 16288 3561 16292
rect 3577 16348 3641 16352
rect 3577 16292 3581 16348
rect 3581 16292 3637 16348
rect 3637 16292 3641 16348
rect 3577 16288 3641 16292
rect 3657 16348 3721 16352
rect 3657 16292 3661 16348
rect 3661 16292 3717 16348
rect 3717 16292 3721 16348
rect 3657 16288 3721 16292
rect 8348 16348 8412 16352
rect 8348 16292 8352 16348
rect 8352 16292 8408 16348
rect 8408 16292 8412 16348
rect 8348 16288 8412 16292
rect 8428 16348 8492 16352
rect 8428 16292 8432 16348
rect 8432 16292 8488 16348
rect 8488 16292 8492 16348
rect 8428 16288 8492 16292
rect 8508 16348 8572 16352
rect 8508 16292 8512 16348
rect 8512 16292 8568 16348
rect 8568 16292 8572 16348
rect 8508 16288 8572 16292
rect 8588 16348 8652 16352
rect 8588 16292 8592 16348
rect 8592 16292 8648 16348
rect 8648 16292 8652 16348
rect 8588 16288 8652 16292
rect 13278 16348 13342 16352
rect 13278 16292 13282 16348
rect 13282 16292 13338 16348
rect 13338 16292 13342 16348
rect 13278 16288 13342 16292
rect 13358 16348 13422 16352
rect 13358 16292 13362 16348
rect 13362 16292 13418 16348
rect 13418 16292 13422 16348
rect 13358 16288 13422 16292
rect 13438 16348 13502 16352
rect 13438 16292 13442 16348
rect 13442 16292 13498 16348
rect 13498 16292 13502 16348
rect 13438 16288 13502 16292
rect 13518 16348 13582 16352
rect 13518 16292 13522 16348
rect 13522 16292 13578 16348
rect 13578 16292 13582 16348
rect 13518 16288 13582 16292
rect 9076 16220 9140 16284
rect 9996 16220 10060 16284
rect 12940 16220 13004 16284
rect 11652 15812 11716 15876
rect 5882 15804 5946 15808
rect 5882 15748 5886 15804
rect 5886 15748 5942 15804
rect 5942 15748 5946 15804
rect 5882 15744 5946 15748
rect 5962 15804 6026 15808
rect 5962 15748 5966 15804
rect 5966 15748 6022 15804
rect 6022 15748 6026 15804
rect 5962 15744 6026 15748
rect 6042 15804 6106 15808
rect 6042 15748 6046 15804
rect 6046 15748 6102 15804
rect 6102 15748 6106 15804
rect 6042 15744 6106 15748
rect 6122 15804 6186 15808
rect 6122 15748 6126 15804
rect 6126 15748 6182 15804
rect 6182 15748 6186 15804
rect 6122 15744 6186 15748
rect 10813 15804 10877 15808
rect 10813 15748 10817 15804
rect 10817 15748 10873 15804
rect 10873 15748 10877 15804
rect 10813 15744 10877 15748
rect 10893 15804 10957 15808
rect 10893 15748 10897 15804
rect 10897 15748 10953 15804
rect 10953 15748 10957 15804
rect 10893 15744 10957 15748
rect 10973 15804 11037 15808
rect 10973 15748 10977 15804
rect 10977 15748 11033 15804
rect 11033 15748 11037 15804
rect 10973 15744 11037 15748
rect 11053 15804 11117 15808
rect 11053 15748 11057 15804
rect 11057 15748 11113 15804
rect 11113 15748 11117 15804
rect 11053 15744 11117 15748
rect 11284 15676 11348 15740
rect 7788 15600 7852 15604
rect 7788 15544 7802 15600
rect 7802 15544 7852 15600
rect 7788 15540 7852 15544
rect 8156 15540 8220 15604
rect 3188 15404 3252 15468
rect 4660 15328 4724 15332
rect 4660 15272 4674 15328
rect 4674 15272 4724 15328
rect 4660 15268 4724 15272
rect 3417 15260 3481 15264
rect 3417 15204 3421 15260
rect 3421 15204 3477 15260
rect 3477 15204 3481 15260
rect 3417 15200 3481 15204
rect 3497 15260 3561 15264
rect 3497 15204 3501 15260
rect 3501 15204 3557 15260
rect 3557 15204 3561 15260
rect 3497 15200 3561 15204
rect 3577 15260 3641 15264
rect 3577 15204 3581 15260
rect 3581 15204 3637 15260
rect 3637 15204 3641 15260
rect 3577 15200 3641 15204
rect 3657 15260 3721 15264
rect 3657 15204 3661 15260
rect 3661 15204 3717 15260
rect 3717 15204 3721 15260
rect 3657 15200 3721 15204
rect 2820 15056 2884 15060
rect 2820 15000 2834 15056
rect 2834 15000 2884 15056
rect 2820 14996 2884 15000
rect 7420 15268 7484 15332
rect 10364 15404 10428 15468
rect 9444 15268 9508 15332
rect 12756 15268 12820 15332
rect 8348 15260 8412 15264
rect 8348 15204 8352 15260
rect 8352 15204 8408 15260
rect 8408 15204 8412 15260
rect 8348 15200 8412 15204
rect 8428 15260 8492 15264
rect 8428 15204 8432 15260
rect 8432 15204 8488 15260
rect 8488 15204 8492 15260
rect 8428 15200 8492 15204
rect 8508 15260 8572 15264
rect 8508 15204 8512 15260
rect 8512 15204 8568 15260
rect 8568 15204 8572 15260
rect 8508 15200 8572 15204
rect 8588 15260 8652 15264
rect 8588 15204 8592 15260
rect 8592 15204 8648 15260
rect 8648 15204 8652 15260
rect 8588 15200 8652 15204
rect 13278 15260 13342 15264
rect 13278 15204 13282 15260
rect 13282 15204 13338 15260
rect 13338 15204 13342 15260
rect 13278 15200 13342 15204
rect 13358 15260 13422 15264
rect 13358 15204 13362 15260
rect 13362 15204 13418 15260
rect 13418 15204 13422 15260
rect 13358 15200 13422 15204
rect 13438 15260 13502 15264
rect 13438 15204 13442 15260
rect 13442 15204 13498 15260
rect 13498 15204 13502 15260
rect 13438 15200 13502 15204
rect 13518 15260 13582 15264
rect 13518 15204 13522 15260
rect 13522 15204 13578 15260
rect 13578 15204 13582 15260
rect 13518 15200 13582 15204
rect 8892 15132 8956 15196
rect 9996 15132 10060 15196
rect 10364 15132 10428 15196
rect 12204 15132 12268 15196
rect 10364 14860 10428 14924
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 6122 14716 6186 14720
rect 6122 14660 6126 14716
rect 6126 14660 6182 14716
rect 6182 14660 6186 14716
rect 6122 14656 6186 14660
rect 9996 14588 10060 14652
rect 13860 14724 13924 14788
rect 10813 14716 10877 14720
rect 10813 14660 10817 14716
rect 10817 14660 10873 14716
rect 10873 14660 10877 14716
rect 10813 14656 10877 14660
rect 10893 14716 10957 14720
rect 10893 14660 10897 14716
rect 10897 14660 10953 14716
rect 10953 14660 10957 14716
rect 10893 14656 10957 14660
rect 10973 14716 11037 14720
rect 10973 14660 10977 14716
rect 10977 14660 11033 14716
rect 11033 14660 11037 14716
rect 10973 14656 11037 14660
rect 11053 14716 11117 14720
rect 11053 14660 11057 14716
rect 11057 14660 11113 14716
rect 11113 14660 11117 14716
rect 11053 14656 11117 14660
rect 12940 14452 13004 14516
rect 10364 14316 10428 14380
rect 10180 14240 10244 14244
rect 10180 14184 10194 14240
rect 10194 14184 10244 14240
rect 10180 14180 10244 14184
rect 10548 14180 10612 14244
rect 3417 14172 3481 14176
rect 3417 14116 3421 14172
rect 3421 14116 3477 14172
rect 3477 14116 3481 14172
rect 3417 14112 3481 14116
rect 3497 14172 3561 14176
rect 3497 14116 3501 14172
rect 3501 14116 3557 14172
rect 3557 14116 3561 14172
rect 3497 14112 3561 14116
rect 3577 14172 3641 14176
rect 3577 14116 3581 14172
rect 3581 14116 3637 14172
rect 3637 14116 3641 14172
rect 3577 14112 3641 14116
rect 3657 14172 3721 14176
rect 3657 14116 3661 14172
rect 3661 14116 3717 14172
rect 3717 14116 3721 14172
rect 3657 14112 3721 14116
rect 8348 14172 8412 14176
rect 8348 14116 8352 14172
rect 8352 14116 8408 14172
rect 8408 14116 8412 14172
rect 8348 14112 8412 14116
rect 8428 14172 8492 14176
rect 8428 14116 8432 14172
rect 8432 14116 8488 14172
rect 8488 14116 8492 14172
rect 8428 14112 8492 14116
rect 8508 14172 8572 14176
rect 8508 14116 8512 14172
rect 8512 14116 8568 14172
rect 8568 14116 8572 14172
rect 8508 14112 8572 14116
rect 8588 14172 8652 14176
rect 8588 14116 8592 14172
rect 8592 14116 8648 14172
rect 8648 14116 8652 14172
rect 8588 14112 8652 14116
rect 13278 14172 13342 14176
rect 13278 14116 13282 14172
rect 13282 14116 13338 14172
rect 13338 14116 13342 14172
rect 13278 14112 13342 14116
rect 13358 14172 13422 14176
rect 13358 14116 13362 14172
rect 13362 14116 13418 14172
rect 13418 14116 13422 14172
rect 13358 14112 13422 14116
rect 13438 14172 13502 14176
rect 13438 14116 13442 14172
rect 13442 14116 13498 14172
rect 13498 14116 13502 14172
rect 13438 14112 13502 14116
rect 13518 14172 13582 14176
rect 13518 14116 13522 14172
rect 13522 14116 13578 14172
rect 13578 14116 13582 14172
rect 13518 14112 13582 14116
rect 8892 13772 8956 13836
rect 10180 13772 10244 13836
rect 12388 13772 12452 13836
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 6122 13628 6186 13632
rect 6122 13572 6126 13628
rect 6126 13572 6182 13628
rect 6182 13572 6186 13628
rect 6122 13568 6186 13572
rect 10813 13628 10877 13632
rect 10813 13572 10817 13628
rect 10817 13572 10873 13628
rect 10873 13572 10877 13628
rect 10813 13568 10877 13572
rect 10893 13628 10957 13632
rect 10893 13572 10897 13628
rect 10897 13572 10953 13628
rect 10953 13572 10957 13628
rect 10893 13568 10957 13572
rect 10973 13628 11037 13632
rect 10973 13572 10977 13628
rect 10977 13572 11033 13628
rect 11033 13572 11037 13628
rect 10973 13568 11037 13572
rect 11053 13628 11117 13632
rect 11053 13572 11057 13628
rect 11057 13572 11113 13628
rect 11113 13572 11117 13628
rect 11053 13568 11117 13572
rect 2820 13500 2884 13564
rect 11836 13500 11900 13564
rect 3417 13084 3481 13088
rect 3417 13028 3421 13084
rect 3421 13028 3477 13084
rect 3477 13028 3481 13084
rect 3417 13024 3481 13028
rect 3497 13084 3561 13088
rect 3497 13028 3501 13084
rect 3501 13028 3557 13084
rect 3557 13028 3561 13084
rect 3497 13024 3561 13028
rect 3577 13084 3641 13088
rect 3577 13028 3581 13084
rect 3581 13028 3637 13084
rect 3637 13028 3641 13084
rect 3577 13024 3641 13028
rect 3657 13084 3721 13088
rect 3657 13028 3661 13084
rect 3661 13028 3717 13084
rect 3717 13028 3721 13084
rect 3657 13024 3721 13028
rect 8348 13084 8412 13088
rect 8348 13028 8352 13084
rect 8352 13028 8408 13084
rect 8408 13028 8412 13084
rect 8348 13024 8412 13028
rect 8428 13084 8492 13088
rect 8428 13028 8432 13084
rect 8432 13028 8488 13084
rect 8488 13028 8492 13084
rect 8428 13024 8492 13028
rect 8508 13084 8572 13088
rect 8508 13028 8512 13084
rect 8512 13028 8568 13084
rect 8568 13028 8572 13084
rect 8508 13024 8572 13028
rect 8588 13084 8652 13088
rect 8588 13028 8592 13084
rect 8592 13028 8648 13084
rect 8648 13028 8652 13084
rect 8588 13024 8652 13028
rect 13278 13084 13342 13088
rect 13278 13028 13282 13084
rect 13282 13028 13338 13084
rect 13338 13028 13342 13084
rect 13278 13024 13342 13028
rect 13358 13084 13422 13088
rect 13358 13028 13362 13084
rect 13362 13028 13418 13084
rect 13418 13028 13422 13084
rect 13358 13024 13422 13028
rect 13438 13084 13502 13088
rect 13438 13028 13442 13084
rect 13442 13028 13498 13084
rect 13498 13028 13502 13084
rect 13438 13024 13502 13028
rect 13518 13084 13582 13088
rect 13518 13028 13522 13084
rect 13522 13028 13578 13084
rect 13578 13028 13582 13084
rect 13518 13024 13582 13028
rect 7972 12956 8036 13020
rect 10180 12956 10244 13020
rect 10548 12956 10612 13020
rect 9628 12548 9692 12612
rect 10548 12548 10612 12612
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 6122 12540 6186 12544
rect 6122 12484 6126 12540
rect 6126 12484 6182 12540
rect 6182 12484 6186 12540
rect 6122 12480 6186 12484
rect 10813 12540 10877 12544
rect 10813 12484 10817 12540
rect 10817 12484 10873 12540
rect 10873 12484 10877 12540
rect 10813 12480 10877 12484
rect 10893 12540 10957 12544
rect 10893 12484 10897 12540
rect 10897 12484 10953 12540
rect 10953 12484 10957 12540
rect 10893 12480 10957 12484
rect 10973 12540 11037 12544
rect 10973 12484 10977 12540
rect 10977 12484 11033 12540
rect 11033 12484 11037 12540
rect 10973 12480 11037 12484
rect 11053 12540 11117 12544
rect 11053 12484 11057 12540
rect 11057 12484 11113 12540
rect 11113 12484 11117 12540
rect 11053 12480 11117 12484
rect 7788 12412 7852 12476
rect 12572 12412 12636 12476
rect 3188 12276 3252 12340
rect 3188 12140 3252 12204
rect 3417 11996 3481 12000
rect 3417 11940 3421 11996
rect 3421 11940 3477 11996
rect 3477 11940 3481 11996
rect 3417 11936 3481 11940
rect 3497 11996 3561 12000
rect 3497 11940 3501 11996
rect 3501 11940 3557 11996
rect 3557 11940 3561 11996
rect 3497 11936 3561 11940
rect 3577 11996 3641 12000
rect 3577 11940 3581 11996
rect 3581 11940 3637 11996
rect 3637 11940 3641 11996
rect 3577 11936 3641 11940
rect 3657 11996 3721 12000
rect 3657 11940 3661 11996
rect 3661 11940 3717 11996
rect 3717 11940 3721 11996
rect 3657 11936 3721 11940
rect 8348 11996 8412 12000
rect 8348 11940 8352 11996
rect 8352 11940 8408 11996
rect 8408 11940 8412 11996
rect 8348 11936 8412 11940
rect 8428 11996 8492 12000
rect 8428 11940 8432 11996
rect 8432 11940 8488 11996
rect 8488 11940 8492 11996
rect 8428 11936 8492 11940
rect 8508 11996 8572 12000
rect 8508 11940 8512 11996
rect 8512 11940 8568 11996
rect 8568 11940 8572 11996
rect 8508 11936 8572 11940
rect 8588 11996 8652 12000
rect 8588 11940 8592 11996
rect 8592 11940 8648 11996
rect 8648 11940 8652 11996
rect 8588 11936 8652 11940
rect 4476 11868 4540 11932
rect 5580 11868 5644 11932
rect 10180 12140 10244 12204
rect 11284 12200 11348 12204
rect 11284 12144 11334 12200
rect 11334 12144 11348 12200
rect 11284 12140 11348 12144
rect 12020 12140 12084 12204
rect 9260 12004 9324 12068
rect 13278 11996 13342 12000
rect 13278 11940 13282 11996
rect 13282 11940 13338 11996
rect 13338 11940 13342 11996
rect 13278 11936 13342 11940
rect 13358 11996 13422 12000
rect 13358 11940 13362 11996
rect 13362 11940 13418 11996
rect 13418 11940 13422 11996
rect 13358 11936 13422 11940
rect 13438 11996 13502 12000
rect 13438 11940 13442 11996
rect 13442 11940 13498 11996
rect 13498 11940 13502 11996
rect 13438 11936 13502 11940
rect 13518 11996 13582 12000
rect 13518 11940 13522 11996
rect 13522 11940 13578 11996
rect 13578 11940 13582 11996
rect 13518 11936 13582 11940
rect 13124 11868 13188 11932
rect 6868 11732 6932 11796
rect 9996 11732 10060 11796
rect 6868 11460 6932 11524
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 6122 11452 6186 11456
rect 6122 11396 6126 11452
rect 6126 11396 6182 11452
rect 6182 11396 6186 11452
rect 6122 11392 6186 11396
rect 10813 11452 10877 11456
rect 10813 11396 10817 11452
rect 10817 11396 10873 11452
rect 10873 11396 10877 11452
rect 10813 11392 10877 11396
rect 10893 11452 10957 11456
rect 10893 11396 10897 11452
rect 10897 11396 10953 11452
rect 10953 11396 10957 11452
rect 10893 11392 10957 11396
rect 10973 11452 11037 11456
rect 10973 11396 10977 11452
rect 10977 11396 11033 11452
rect 11033 11396 11037 11452
rect 10973 11392 11037 11396
rect 11053 11452 11117 11456
rect 11053 11396 11057 11452
rect 11057 11396 11113 11452
rect 11113 11396 11117 11452
rect 11053 11392 11117 11396
rect 11284 11324 11348 11388
rect 9996 11112 10060 11116
rect 9996 11056 10010 11112
rect 10010 11056 10060 11112
rect 9996 11052 10060 11056
rect 3417 10908 3481 10912
rect 3417 10852 3421 10908
rect 3421 10852 3477 10908
rect 3477 10852 3481 10908
rect 3417 10848 3481 10852
rect 3497 10908 3561 10912
rect 3497 10852 3501 10908
rect 3501 10852 3557 10908
rect 3557 10852 3561 10908
rect 3497 10848 3561 10852
rect 3577 10908 3641 10912
rect 3577 10852 3581 10908
rect 3581 10852 3637 10908
rect 3637 10852 3641 10908
rect 3577 10848 3641 10852
rect 3657 10908 3721 10912
rect 3657 10852 3661 10908
rect 3661 10852 3717 10908
rect 3717 10852 3721 10908
rect 3657 10848 3721 10852
rect 8348 10908 8412 10912
rect 8348 10852 8352 10908
rect 8352 10852 8408 10908
rect 8408 10852 8412 10908
rect 8348 10848 8412 10852
rect 8428 10908 8492 10912
rect 8428 10852 8432 10908
rect 8432 10852 8488 10908
rect 8488 10852 8492 10908
rect 8428 10848 8492 10852
rect 8508 10908 8572 10912
rect 8508 10852 8512 10908
rect 8512 10852 8568 10908
rect 8568 10852 8572 10908
rect 8508 10848 8572 10852
rect 8588 10908 8652 10912
rect 8588 10852 8592 10908
rect 8592 10852 8648 10908
rect 8648 10852 8652 10908
rect 8588 10848 8652 10852
rect 13278 10908 13342 10912
rect 13278 10852 13282 10908
rect 13282 10852 13338 10908
rect 13338 10852 13342 10908
rect 13278 10848 13342 10852
rect 13358 10908 13422 10912
rect 13358 10852 13362 10908
rect 13362 10852 13418 10908
rect 13418 10852 13422 10908
rect 13358 10848 13422 10852
rect 13438 10908 13502 10912
rect 13438 10852 13442 10908
rect 13442 10852 13498 10908
rect 13498 10852 13502 10908
rect 13438 10848 13502 10852
rect 13518 10908 13582 10912
rect 13518 10852 13522 10908
rect 13522 10852 13578 10908
rect 13578 10852 13582 10908
rect 13518 10848 13582 10852
rect 9444 10780 9508 10844
rect 8156 10508 8220 10572
rect 12020 10372 12084 10436
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 6122 10364 6186 10368
rect 6122 10308 6126 10364
rect 6126 10308 6182 10364
rect 6182 10308 6186 10364
rect 6122 10304 6186 10308
rect 10813 10364 10877 10368
rect 10813 10308 10817 10364
rect 10817 10308 10873 10364
rect 10873 10308 10877 10364
rect 10813 10304 10877 10308
rect 10893 10364 10957 10368
rect 10893 10308 10897 10364
rect 10897 10308 10953 10364
rect 10953 10308 10957 10364
rect 10893 10304 10957 10308
rect 10973 10364 11037 10368
rect 10973 10308 10977 10364
rect 10977 10308 11033 10364
rect 11033 10308 11037 10364
rect 10973 10304 11037 10308
rect 11053 10364 11117 10368
rect 11053 10308 11057 10364
rect 11057 10308 11113 10364
rect 11113 10308 11117 10364
rect 11053 10304 11117 10308
rect 10548 10100 10612 10164
rect 12388 10100 12452 10164
rect 3417 9820 3481 9824
rect 3417 9764 3421 9820
rect 3421 9764 3477 9820
rect 3477 9764 3481 9820
rect 3417 9760 3481 9764
rect 3497 9820 3561 9824
rect 3497 9764 3501 9820
rect 3501 9764 3557 9820
rect 3557 9764 3561 9820
rect 3497 9760 3561 9764
rect 3577 9820 3641 9824
rect 3577 9764 3581 9820
rect 3581 9764 3637 9820
rect 3637 9764 3641 9820
rect 3577 9760 3641 9764
rect 3657 9820 3721 9824
rect 3657 9764 3661 9820
rect 3661 9764 3717 9820
rect 3717 9764 3721 9820
rect 3657 9760 3721 9764
rect 8348 9820 8412 9824
rect 8348 9764 8352 9820
rect 8352 9764 8408 9820
rect 8408 9764 8412 9820
rect 8348 9760 8412 9764
rect 8428 9820 8492 9824
rect 8428 9764 8432 9820
rect 8432 9764 8488 9820
rect 8488 9764 8492 9820
rect 8428 9760 8492 9764
rect 8508 9820 8572 9824
rect 8508 9764 8512 9820
rect 8512 9764 8568 9820
rect 8568 9764 8572 9820
rect 8508 9760 8572 9764
rect 8588 9820 8652 9824
rect 8588 9764 8592 9820
rect 8592 9764 8648 9820
rect 8648 9764 8652 9820
rect 8588 9760 8652 9764
rect 13278 9820 13342 9824
rect 13278 9764 13282 9820
rect 13282 9764 13338 9820
rect 13338 9764 13342 9820
rect 13278 9760 13342 9764
rect 13358 9820 13422 9824
rect 13358 9764 13362 9820
rect 13362 9764 13418 9820
rect 13418 9764 13422 9820
rect 13358 9760 13422 9764
rect 13438 9820 13502 9824
rect 13438 9764 13442 9820
rect 13442 9764 13498 9820
rect 13498 9764 13502 9820
rect 13438 9760 13502 9764
rect 13518 9820 13582 9824
rect 13518 9764 13522 9820
rect 13522 9764 13578 9820
rect 13578 9764 13582 9820
rect 13518 9760 13582 9764
rect 11468 9692 11532 9756
rect 11652 9752 11716 9756
rect 11652 9696 11666 9752
rect 11666 9696 11716 9752
rect 11652 9692 11716 9696
rect 14412 9556 14476 9620
rect 10180 9284 10244 9348
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 6122 9276 6186 9280
rect 6122 9220 6126 9276
rect 6126 9220 6182 9276
rect 6182 9220 6186 9276
rect 6122 9216 6186 9220
rect 10813 9276 10877 9280
rect 10813 9220 10817 9276
rect 10817 9220 10873 9276
rect 10873 9220 10877 9276
rect 10813 9216 10877 9220
rect 10893 9276 10957 9280
rect 10893 9220 10897 9276
rect 10897 9220 10953 9276
rect 10953 9220 10957 9276
rect 10893 9216 10957 9220
rect 10973 9276 11037 9280
rect 10973 9220 10977 9276
rect 10977 9220 11033 9276
rect 11033 9220 11037 9276
rect 10973 9216 11037 9220
rect 11053 9276 11117 9280
rect 11053 9220 11057 9276
rect 11057 9220 11113 9276
rect 11113 9220 11117 9276
rect 11053 9216 11117 9220
rect 3004 9148 3068 9212
rect 6316 9208 6380 9212
rect 6316 9152 6366 9208
rect 6366 9152 6380 9208
rect 6316 9148 6380 9152
rect 6684 9148 6748 9212
rect 14228 9148 14292 9212
rect 3417 8732 3481 8736
rect 3417 8676 3421 8732
rect 3421 8676 3477 8732
rect 3477 8676 3481 8732
rect 3417 8672 3481 8676
rect 3497 8732 3561 8736
rect 3497 8676 3501 8732
rect 3501 8676 3557 8732
rect 3557 8676 3561 8732
rect 3497 8672 3561 8676
rect 3577 8732 3641 8736
rect 3577 8676 3581 8732
rect 3581 8676 3637 8732
rect 3637 8676 3641 8732
rect 3577 8672 3641 8676
rect 3657 8732 3721 8736
rect 3657 8676 3661 8732
rect 3661 8676 3717 8732
rect 3717 8676 3721 8732
rect 3657 8672 3721 8676
rect 12388 8740 12452 8804
rect 8348 8732 8412 8736
rect 8348 8676 8352 8732
rect 8352 8676 8408 8732
rect 8408 8676 8412 8732
rect 8348 8672 8412 8676
rect 8428 8732 8492 8736
rect 8428 8676 8432 8732
rect 8432 8676 8488 8732
rect 8488 8676 8492 8732
rect 8428 8672 8492 8676
rect 8508 8732 8572 8736
rect 8508 8676 8512 8732
rect 8512 8676 8568 8732
rect 8568 8676 8572 8732
rect 8508 8672 8572 8676
rect 8588 8732 8652 8736
rect 8588 8676 8592 8732
rect 8592 8676 8648 8732
rect 8648 8676 8652 8732
rect 8588 8672 8652 8676
rect 13278 8732 13342 8736
rect 13278 8676 13282 8732
rect 13282 8676 13338 8732
rect 13338 8676 13342 8732
rect 13278 8672 13342 8676
rect 13358 8732 13422 8736
rect 13358 8676 13362 8732
rect 13362 8676 13418 8732
rect 13418 8676 13422 8732
rect 13358 8672 13422 8676
rect 13438 8732 13502 8736
rect 13438 8676 13442 8732
rect 13442 8676 13498 8732
rect 13498 8676 13502 8732
rect 13438 8672 13502 8676
rect 13518 8732 13582 8736
rect 13518 8676 13522 8732
rect 13522 8676 13578 8732
rect 13578 8676 13582 8732
rect 13518 8672 13582 8676
rect 6500 8468 6564 8532
rect 7972 8528 8036 8532
rect 9996 8604 10060 8668
rect 11652 8604 11716 8668
rect 12020 8604 12084 8668
rect 7972 8472 8022 8528
rect 8022 8472 8036 8528
rect 7972 8468 8036 8472
rect 9628 8468 9692 8532
rect 9260 8196 9324 8260
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 6122 8188 6186 8192
rect 6122 8132 6126 8188
rect 6126 8132 6182 8188
rect 6182 8132 6186 8188
rect 6122 8128 6186 8132
rect 10813 8188 10877 8192
rect 10813 8132 10817 8188
rect 10817 8132 10873 8188
rect 10873 8132 10877 8188
rect 10813 8128 10877 8132
rect 10893 8188 10957 8192
rect 10893 8132 10897 8188
rect 10897 8132 10953 8188
rect 10953 8132 10957 8188
rect 10893 8128 10957 8132
rect 10973 8188 11037 8192
rect 10973 8132 10977 8188
rect 10977 8132 11033 8188
rect 11033 8132 11037 8188
rect 10973 8128 11037 8132
rect 11053 8188 11117 8192
rect 11053 8132 11057 8188
rect 11057 8132 11113 8188
rect 11113 8132 11117 8188
rect 11053 8128 11117 8132
rect 11836 8120 11900 8124
rect 11836 8064 11886 8120
rect 11886 8064 11900 8120
rect 11836 8060 11900 8064
rect 11836 7924 11900 7988
rect 12572 7788 12636 7852
rect 5212 7652 5276 7716
rect 7972 7652 8036 7716
rect 9260 7652 9324 7716
rect 3417 7644 3481 7648
rect 3417 7588 3421 7644
rect 3421 7588 3477 7644
rect 3477 7588 3481 7644
rect 3417 7584 3481 7588
rect 3497 7644 3561 7648
rect 3497 7588 3501 7644
rect 3501 7588 3557 7644
rect 3557 7588 3561 7644
rect 3497 7584 3561 7588
rect 3577 7644 3641 7648
rect 3577 7588 3581 7644
rect 3581 7588 3637 7644
rect 3637 7588 3641 7644
rect 3577 7584 3641 7588
rect 3657 7644 3721 7648
rect 3657 7588 3661 7644
rect 3661 7588 3717 7644
rect 3717 7588 3721 7644
rect 3657 7584 3721 7588
rect 8348 7644 8412 7648
rect 8348 7588 8352 7644
rect 8352 7588 8408 7644
rect 8408 7588 8412 7644
rect 8348 7584 8412 7588
rect 8428 7644 8492 7648
rect 8428 7588 8432 7644
rect 8432 7588 8488 7644
rect 8488 7588 8492 7644
rect 8428 7584 8492 7588
rect 8508 7644 8572 7648
rect 8508 7588 8512 7644
rect 8512 7588 8568 7644
rect 8568 7588 8572 7644
rect 8508 7584 8572 7588
rect 8588 7644 8652 7648
rect 8588 7588 8592 7644
rect 8592 7588 8648 7644
rect 8648 7588 8652 7644
rect 8588 7584 8652 7588
rect 13278 7644 13342 7648
rect 13278 7588 13282 7644
rect 13282 7588 13338 7644
rect 13338 7588 13342 7644
rect 13278 7584 13342 7588
rect 13358 7644 13422 7648
rect 13358 7588 13362 7644
rect 13362 7588 13418 7644
rect 13418 7588 13422 7644
rect 13358 7584 13422 7588
rect 13438 7644 13502 7648
rect 13438 7588 13442 7644
rect 13442 7588 13498 7644
rect 13498 7588 13502 7644
rect 13438 7584 13502 7588
rect 13518 7644 13582 7648
rect 13518 7588 13522 7644
rect 13522 7588 13578 7644
rect 13578 7588 13582 7644
rect 13518 7584 13582 7588
rect 4844 7576 4908 7580
rect 4844 7520 4858 7576
rect 4858 7520 4908 7576
rect 4844 7516 4908 7520
rect 7604 7576 7668 7580
rect 7604 7520 7654 7576
rect 7654 7520 7668 7576
rect 7604 7516 7668 7520
rect 5028 7380 5092 7444
rect 6500 7380 6564 7444
rect 13124 7244 13188 7308
rect 7236 7108 7300 7172
rect 14044 7108 14108 7172
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 6122 7100 6186 7104
rect 6122 7044 6126 7100
rect 6126 7044 6182 7100
rect 6182 7044 6186 7100
rect 6122 7040 6186 7044
rect 10813 7100 10877 7104
rect 10813 7044 10817 7100
rect 10817 7044 10873 7100
rect 10873 7044 10877 7100
rect 10813 7040 10877 7044
rect 10893 7100 10957 7104
rect 10893 7044 10897 7100
rect 10897 7044 10953 7100
rect 10953 7044 10957 7100
rect 10893 7040 10957 7044
rect 10973 7100 11037 7104
rect 10973 7044 10977 7100
rect 10977 7044 11033 7100
rect 11033 7044 11037 7100
rect 10973 7040 11037 7044
rect 11053 7100 11117 7104
rect 11053 7044 11057 7100
rect 11057 7044 11113 7100
rect 11113 7044 11117 7100
rect 11053 7040 11117 7044
rect 6500 6972 6564 7036
rect 7604 6836 7668 6900
rect 7972 6836 8036 6900
rect 11652 6836 11716 6900
rect 12572 6972 12636 7036
rect 13676 6836 13740 6900
rect 7052 6564 7116 6628
rect 9812 6700 9876 6764
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 3004 6488 3068 6492
rect 3004 6432 3054 6488
rect 3054 6432 3068 6488
rect 3004 6428 3068 6432
rect 7972 6428 8036 6492
rect 9812 6428 9876 6492
rect 6316 6292 6380 6356
rect 13860 6292 13924 6356
rect 4292 6156 4356 6220
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 7972 5884 8036 5948
rect 11836 5884 11900 5948
rect 12572 5884 12636 5948
rect 12940 5884 13004 5948
rect 7420 5748 7484 5812
rect 7604 5748 7668 5812
rect 5396 5672 5460 5676
rect 5396 5616 5410 5672
rect 5410 5616 5460 5672
rect 5396 5612 5460 5616
rect 7788 5612 7852 5676
rect 7788 5476 7852 5540
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 4476 5340 4540 5404
rect 9076 5476 9140 5540
rect 12204 5612 12268 5676
rect 11652 5476 11716 5540
rect 12204 5476 12268 5540
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 9628 5340 9692 5404
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 9628 5068 9692 5132
rect 10180 4932 10244 4996
rect 12572 4932 12636 4996
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 5028 4796 5092 4860
rect 4108 4660 4172 4724
rect 9628 4796 9692 4860
rect 10180 4856 10244 4860
rect 10180 4800 10194 4856
rect 10194 4800 10244 4856
rect 10180 4796 10244 4800
rect 7420 4660 7484 4724
rect 12940 4660 13004 4724
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 4476 4252 4540 4316
rect 4844 4312 4908 4316
rect 4844 4256 4858 4312
rect 4858 4256 4908 4312
rect 4844 4252 4908 4256
rect 7788 4252 7852 4316
rect 7788 4116 7852 4180
rect 4292 3980 4356 4044
rect 7052 3980 7116 4044
rect 7236 3980 7300 4044
rect 9260 4388 9324 4452
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 9076 4252 9140 4316
rect 12020 4252 12084 4316
rect 10364 4176 10428 4180
rect 10364 4120 10414 4176
rect 10414 4120 10428 4176
rect 10364 4116 10428 4120
rect 11468 3980 11532 4044
rect 14228 4524 14292 4588
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 5580 3844 5644 3908
rect 11468 3844 11532 3908
rect 12020 3844 12084 3908
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 5580 3708 5644 3772
rect 9812 3708 9876 3772
rect 12204 3708 12268 3772
rect 3188 3572 3252 3636
rect 3924 3572 3988 3636
rect 3188 3496 3252 3500
rect 3188 3440 3238 3496
rect 3238 3440 3252 3496
rect 3188 3436 3252 3440
rect 5028 3436 5092 3500
rect 12572 3572 12636 3636
rect 13124 3572 13188 3636
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 3924 3224 3988 3228
rect 3924 3168 3938 3224
rect 3938 3168 3988 3224
rect 3924 3164 3988 3168
rect 5580 3164 5644 3228
rect 9076 3164 9140 3228
rect 11284 3164 11348 3228
rect 11468 3164 11532 3228
rect 12388 3164 12452 3228
rect 14412 3164 14476 3228
rect 12020 3028 12084 3092
rect 3924 2816 3988 2820
rect 3924 2760 3974 2816
rect 3974 2760 3988 2816
rect 3924 2756 3988 2760
rect 4476 2756 4540 2820
rect 8892 2756 8956 2820
rect 9628 2756 9692 2820
rect 10548 2816 10612 2820
rect 10548 2760 10598 2816
rect 10598 2760 10612 2816
rect 10548 2756 10612 2760
rect 11468 2756 11532 2820
rect 11836 2816 11900 2820
rect 11836 2760 11850 2816
rect 11850 2760 11900 2816
rect 11836 2756 11900 2760
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 4660 2620 4724 2684
rect 5212 2620 5276 2684
rect 6684 2620 6748 2684
rect 8156 2620 8220 2684
rect 10180 2620 10244 2684
rect 12756 2620 12820 2684
rect 14044 2680 14108 2684
rect 14044 2624 14058 2680
rect 14058 2624 14108 2680
rect 14044 2620 14108 2624
rect 6868 2348 6932 2412
rect 7604 2212 7668 2276
rect 7788 2212 7852 2276
rect 9260 2212 9324 2276
rect 11468 2212 11532 2276
rect 13860 2272 13924 2276
rect 13860 2216 13874 2272
rect 13874 2216 13924 2272
rect 13860 2212 13924 2216
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
rect 12204 2076 12268 2140
rect 3924 1804 3988 1868
rect 4108 1668 4172 1732
rect 5396 1668 5460 1732
rect 11652 1532 11716 1596
rect 3188 1396 3252 1460
rect 9076 1396 9140 1460
rect 10364 1396 10428 1460
rect 7420 1260 7484 1324
rect 12940 1260 13004 1324
rect 6316 1124 6380 1188
rect 7972 1124 8036 1188
rect 13676 1124 13740 1188
rect 9996 988 10060 1052
<< metal4 >>
rect 8891 17780 8957 17781
rect 8891 17716 8892 17780
rect 8956 17716 8957 17780
rect 8891 17715 8957 17716
rect 8155 17644 8221 17645
rect 8155 17580 8156 17644
rect 8220 17580 8221 17644
rect 8155 17579 8221 17580
rect 3409 17440 3729 17456
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 16352 3729 17376
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3187 15468 3253 15469
rect 3187 15404 3188 15468
rect 3252 15404 3253 15468
rect 3187 15403 3253 15404
rect 2819 15060 2885 15061
rect 2819 14996 2820 15060
rect 2884 14996 2885 15060
rect 2819 14995 2885 14996
rect 2822 13565 2882 14995
rect 2819 13564 2885 13565
rect 2819 13500 2820 13564
rect 2884 13500 2885 13564
rect 2819 13499 2885 13500
rect 3190 12341 3250 15403
rect 3409 15264 3729 16288
rect 5874 16896 6195 17456
rect 7971 17236 8037 17237
rect 7971 17172 7972 17236
rect 8036 17172 8037 17236
rect 7971 17171 8037 17172
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6195 16896
rect 5874 15808 6195 16832
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6195 15808
rect 4659 15332 4725 15333
rect 4659 15268 4660 15332
rect 4724 15268 4725 15332
rect 4659 15267 4725 15268
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 14176 3729 15200
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 13088 3729 14112
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3187 12340 3253 12341
rect 3187 12276 3188 12340
rect 3252 12276 3253 12340
rect 3187 12275 3253 12276
rect 3187 12204 3253 12205
rect 3187 12140 3188 12204
rect 3252 12140 3253 12204
rect 3187 12139 3253 12140
rect 3003 9212 3069 9213
rect 3003 9148 3004 9212
rect 3068 9148 3069 9212
rect 3003 9147 3069 9148
rect 3006 6493 3066 9147
rect 3003 6492 3069 6493
rect 3003 6428 3004 6492
rect 3068 6428 3069 6492
rect 3003 6427 3069 6428
rect 3190 3637 3250 12139
rect 3409 12000 3729 13024
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 10912 3729 11936
rect 4475 11932 4541 11933
rect 4475 11868 4476 11932
rect 4540 11868 4541 11932
rect 4475 11867 4541 11868
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 9824 3729 10848
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 8736 3729 9760
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 7648 3729 8672
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 6560 3729 7584
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 5472 3729 6496
rect 4291 6220 4357 6221
rect 4291 6156 4292 6220
rect 4356 6156 4357 6220
rect 4291 6155 4357 6156
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 4107 4724 4173 4725
rect 4107 4660 4108 4724
rect 4172 4660 4173 4724
rect 4107 4659 4173 4660
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3187 3636 3253 3637
rect 3187 3572 3188 3636
rect 3252 3572 3253 3636
rect 3187 3571 3253 3572
rect 3187 3500 3253 3501
rect 3187 3436 3188 3500
rect 3252 3436 3253 3500
rect 3187 3435 3253 3436
rect 3190 1461 3250 3435
rect 3409 3296 3729 4320
rect 3923 3636 3989 3637
rect 3923 3572 3924 3636
rect 3988 3572 3989 3636
rect 3923 3571 3989 3572
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 2208 3729 3232
rect 3926 3229 3986 3571
rect 3923 3228 3989 3229
rect 3923 3164 3924 3228
rect 3988 3164 3989 3228
rect 3923 3163 3989 3164
rect 3923 2820 3989 2821
rect 3923 2756 3924 2820
rect 3988 2756 3989 2820
rect 3923 2755 3989 2756
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 3926 1869 3986 2755
rect 3923 1868 3989 1869
rect 3923 1804 3924 1868
rect 3988 1804 3989 1868
rect 3923 1803 3989 1804
rect 4110 1733 4170 4659
rect 4294 4045 4354 6155
rect 4478 5405 4538 11867
rect 4475 5404 4541 5405
rect 4475 5340 4476 5404
rect 4540 5340 4541 5404
rect 4475 5339 4541 5340
rect 4475 4316 4541 4317
rect 4475 4252 4476 4316
rect 4540 4252 4541 4316
rect 4475 4251 4541 4252
rect 4291 4044 4357 4045
rect 4291 3980 4292 4044
rect 4356 3980 4357 4044
rect 4291 3979 4357 3980
rect 4478 2821 4538 4251
rect 4475 2820 4541 2821
rect 4475 2756 4476 2820
rect 4540 2756 4541 2820
rect 4475 2755 4541 2756
rect 4662 2685 4722 15267
rect 5874 14720 6195 15744
rect 7787 15604 7853 15605
rect 7787 15540 7788 15604
rect 7852 15540 7853 15604
rect 7787 15539 7853 15540
rect 7419 15332 7485 15333
rect 7419 15268 7420 15332
rect 7484 15268 7485 15332
rect 7419 15267 7485 15268
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6195 14720
rect 5874 13632 6195 14656
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6195 13632
rect 5874 12544 6195 13568
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6195 12544
rect 5579 11932 5645 11933
rect 5579 11868 5580 11932
rect 5644 11868 5645 11932
rect 5579 11867 5645 11868
rect 5211 7716 5277 7717
rect 5211 7652 5212 7716
rect 5276 7652 5277 7716
rect 5211 7651 5277 7652
rect 4843 7580 4909 7581
rect 4843 7516 4844 7580
rect 4908 7516 4909 7580
rect 4843 7515 4909 7516
rect 4846 4317 4906 7515
rect 5027 7444 5093 7445
rect 5027 7380 5028 7444
rect 5092 7380 5093 7444
rect 5027 7379 5093 7380
rect 5030 4861 5090 7379
rect 5027 4860 5093 4861
rect 5027 4796 5028 4860
rect 5092 4796 5093 4860
rect 5027 4795 5093 4796
rect 4843 4316 4909 4317
rect 4843 4252 4844 4316
rect 4908 4252 4909 4316
rect 4843 4251 4909 4252
rect 5030 3501 5090 4795
rect 5027 3500 5093 3501
rect 5027 3436 5028 3500
rect 5092 3436 5093 3500
rect 5027 3435 5093 3436
rect 5214 2685 5274 7651
rect 5395 5676 5461 5677
rect 5395 5612 5396 5676
rect 5460 5612 5461 5676
rect 5395 5611 5461 5612
rect 4659 2684 4725 2685
rect 4659 2620 4660 2684
rect 4724 2620 4725 2684
rect 4659 2619 4725 2620
rect 5211 2684 5277 2685
rect 5211 2620 5212 2684
rect 5276 2620 5277 2684
rect 5211 2619 5277 2620
rect 5398 1733 5458 5611
rect 5582 3909 5642 11867
rect 5874 11456 6195 12480
rect 6867 11796 6933 11797
rect 6867 11732 6868 11796
rect 6932 11732 6933 11796
rect 6867 11731 6933 11732
rect 6870 11525 6930 11731
rect 6867 11524 6933 11525
rect 6867 11460 6868 11524
rect 6932 11460 6933 11524
rect 6867 11459 6933 11460
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6195 11456
rect 5874 10368 6195 11392
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6195 10368
rect 5874 9280 6195 10304
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6195 9280
rect 5874 8192 6195 9216
rect 6315 9212 6381 9213
rect 6315 9148 6316 9212
rect 6380 9148 6381 9212
rect 6315 9147 6381 9148
rect 6683 9212 6749 9213
rect 6683 9148 6684 9212
rect 6748 9148 6749 9212
rect 6683 9147 6749 9148
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6195 8192
rect 5874 7104 6195 8128
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6195 7104
rect 5874 6016 6195 7040
rect 6318 6357 6378 9147
rect 6499 8532 6565 8533
rect 6499 8468 6500 8532
rect 6564 8468 6565 8532
rect 6499 8467 6565 8468
rect 6502 7445 6562 8467
rect 6499 7444 6565 7445
rect 6499 7380 6500 7444
rect 6564 7380 6565 7444
rect 6499 7379 6565 7380
rect 6499 7036 6565 7037
rect 6499 6972 6500 7036
rect 6564 6972 6565 7036
rect 6499 6971 6565 6972
rect 6315 6356 6381 6357
rect 6315 6292 6316 6356
rect 6380 6292 6381 6356
rect 6315 6291 6381 6292
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5579 3908 5645 3909
rect 5579 3844 5580 3908
rect 5644 3844 5645 3908
rect 5579 3843 5645 3844
rect 5874 3840 6195 4864
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5579 3772 5645 3773
rect 5579 3708 5580 3772
rect 5644 3708 5645 3772
rect 5579 3707 5645 3708
rect 5582 3229 5642 3707
rect 5579 3228 5645 3229
rect 5579 3164 5580 3228
rect 5644 3164 5645 3228
rect 5579 3163 5645 3164
rect 5874 2752 6195 3776
rect 6502 3090 6562 6971
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 5874 2128 6195 2688
rect 6318 3030 6562 3090
rect 4107 1732 4173 1733
rect 4107 1668 4108 1732
rect 4172 1668 4173 1732
rect 4107 1667 4173 1668
rect 5395 1732 5461 1733
rect 5395 1668 5396 1732
rect 5460 1668 5461 1732
rect 5395 1667 5461 1668
rect 3187 1460 3253 1461
rect 3187 1396 3188 1460
rect 3252 1396 3253 1460
rect 3187 1395 3253 1396
rect 6318 1189 6378 3030
rect 6686 2685 6746 9147
rect 6683 2684 6749 2685
rect 6683 2620 6684 2684
rect 6748 2620 6749 2684
rect 6683 2619 6749 2620
rect 6870 2413 6930 11459
rect 7235 7172 7301 7173
rect 7235 7108 7236 7172
rect 7300 7108 7301 7172
rect 7235 7107 7301 7108
rect 7051 6628 7117 6629
rect 7051 6564 7052 6628
rect 7116 6564 7117 6628
rect 7051 6563 7117 6564
rect 7054 4045 7114 6563
rect 7238 4045 7298 7107
rect 7422 5813 7482 15267
rect 7790 12477 7850 15539
rect 7974 13021 8034 17171
rect 8158 15605 8218 17579
rect 8340 17440 8660 17456
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 16352 8660 17376
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8155 15604 8221 15605
rect 8155 15540 8156 15604
rect 8220 15540 8221 15604
rect 8155 15539 8221 15540
rect 8340 15264 8660 16288
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 14176 8660 15200
rect 8894 15197 8954 17715
rect 10363 17508 10429 17509
rect 10363 17444 10364 17508
rect 10428 17444 10429 17508
rect 10363 17443 10429 17444
rect 10179 16828 10245 16829
rect 10179 16764 10180 16828
rect 10244 16764 10245 16828
rect 10179 16763 10245 16764
rect 9811 16692 9877 16693
rect 9811 16628 9812 16692
rect 9876 16628 9877 16692
rect 9811 16627 9877 16628
rect 9627 16556 9693 16557
rect 9627 16492 9628 16556
rect 9692 16492 9693 16556
rect 9627 16491 9693 16492
rect 9075 16284 9141 16285
rect 9075 16220 9076 16284
rect 9140 16220 9141 16284
rect 9075 16219 9141 16220
rect 8891 15196 8957 15197
rect 8891 15132 8892 15196
rect 8956 15132 8957 15196
rect 8891 15131 8957 15132
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 13088 8660 14112
rect 8891 13836 8957 13837
rect 8891 13772 8892 13836
rect 8956 13772 8957 13836
rect 8891 13771 8957 13772
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 7971 13020 8037 13021
rect 7971 12956 7972 13020
rect 8036 12956 8037 13020
rect 7971 12955 8037 12956
rect 7787 12476 7853 12477
rect 7787 12412 7788 12476
rect 7852 12412 7853 12476
rect 7787 12411 7853 12412
rect 7974 8533 8034 12955
rect 8340 12000 8660 13024
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 10912 8660 11936
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8155 10572 8221 10573
rect 8155 10508 8156 10572
rect 8220 10508 8221 10572
rect 8155 10507 8221 10508
rect 7971 8532 8037 8533
rect 7971 8530 7972 8532
rect 7790 8470 7972 8530
rect 7603 7580 7669 7581
rect 7603 7516 7604 7580
rect 7668 7516 7669 7580
rect 7603 7515 7669 7516
rect 7606 6901 7666 7515
rect 7603 6900 7669 6901
rect 7603 6836 7604 6900
rect 7668 6836 7669 6900
rect 7603 6835 7669 6836
rect 7419 5812 7485 5813
rect 7419 5748 7420 5812
rect 7484 5748 7485 5812
rect 7419 5747 7485 5748
rect 7603 5812 7669 5813
rect 7603 5748 7604 5812
rect 7668 5748 7669 5812
rect 7603 5747 7669 5748
rect 7419 4724 7485 4725
rect 7419 4660 7420 4724
rect 7484 4660 7485 4724
rect 7419 4659 7485 4660
rect 7051 4044 7117 4045
rect 7051 3980 7052 4044
rect 7116 3980 7117 4044
rect 7051 3979 7117 3980
rect 7235 4044 7301 4045
rect 7235 3980 7236 4044
rect 7300 3980 7301 4044
rect 7235 3979 7301 3980
rect 6867 2412 6933 2413
rect 6867 2348 6868 2412
rect 6932 2348 6933 2412
rect 6867 2347 6933 2348
rect 7422 1325 7482 4659
rect 7606 2277 7666 5747
rect 7790 5677 7850 8470
rect 7971 8468 7972 8470
rect 8036 8468 8037 8532
rect 7971 8467 8037 8468
rect 7971 7716 8037 7717
rect 7971 7652 7972 7716
rect 8036 7652 8037 7716
rect 7971 7651 8037 7652
rect 7974 6901 8034 7651
rect 7971 6900 8037 6901
rect 7971 6836 7972 6900
rect 8036 6836 8037 6900
rect 7971 6835 8037 6836
rect 7971 6492 8037 6493
rect 7971 6428 7972 6492
rect 8036 6428 8037 6492
rect 7971 6427 8037 6428
rect 7974 5949 8034 6427
rect 7971 5948 8037 5949
rect 7971 5884 7972 5948
rect 8036 5884 8037 5948
rect 7971 5883 8037 5884
rect 7787 5676 7853 5677
rect 7787 5612 7788 5676
rect 7852 5674 7853 5676
rect 7852 5614 8034 5674
rect 7852 5612 7853 5614
rect 7787 5611 7853 5612
rect 7787 5540 7853 5541
rect 7787 5476 7788 5540
rect 7852 5476 7853 5540
rect 7787 5475 7853 5476
rect 7790 4317 7850 5475
rect 7787 4316 7853 4317
rect 7787 4252 7788 4316
rect 7852 4252 7853 4316
rect 7787 4251 7853 4252
rect 7787 4180 7853 4181
rect 7787 4116 7788 4180
rect 7852 4116 7853 4180
rect 7787 4115 7853 4116
rect 7790 2277 7850 4115
rect 7603 2276 7669 2277
rect 7603 2212 7604 2276
rect 7668 2212 7669 2276
rect 7603 2211 7669 2212
rect 7787 2276 7853 2277
rect 7787 2212 7788 2276
rect 7852 2212 7853 2276
rect 7787 2211 7853 2212
rect 7419 1324 7485 1325
rect 7419 1260 7420 1324
rect 7484 1260 7485 1324
rect 7419 1259 7485 1260
rect 7974 1189 8034 5614
rect 8158 2685 8218 10507
rect 8340 9824 8660 10848
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 8736 8660 9760
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 7648 8660 8672
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 6560 8660 7584
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 5472 8660 6496
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 3296 8660 4320
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8155 2684 8221 2685
rect 8155 2620 8156 2684
rect 8220 2620 8221 2684
rect 8155 2619 8221 2620
rect 8340 2208 8660 3232
rect 8894 2821 8954 13771
rect 9078 5541 9138 16219
rect 9443 15332 9509 15333
rect 9443 15268 9444 15332
rect 9508 15268 9509 15332
rect 9443 15267 9509 15268
rect 9259 12068 9325 12069
rect 9259 12004 9260 12068
rect 9324 12004 9325 12068
rect 9259 12003 9325 12004
rect 9262 8261 9322 12003
rect 9446 10845 9506 15267
rect 9630 12613 9690 16491
rect 9627 12612 9693 12613
rect 9627 12548 9628 12612
rect 9692 12548 9693 12612
rect 9627 12547 9693 12548
rect 9443 10844 9509 10845
rect 9443 10780 9444 10844
rect 9508 10780 9509 10844
rect 9443 10779 9509 10780
rect 9627 8532 9693 8533
rect 9627 8468 9628 8532
rect 9692 8468 9693 8532
rect 9627 8467 9693 8468
rect 9259 8260 9325 8261
rect 9259 8196 9260 8260
rect 9324 8196 9325 8260
rect 9259 8195 9325 8196
rect 9259 7716 9325 7717
rect 9259 7652 9260 7716
rect 9324 7652 9325 7716
rect 9259 7651 9325 7652
rect 9075 5540 9141 5541
rect 9075 5476 9076 5540
rect 9140 5476 9141 5540
rect 9075 5475 9141 5476
rect 9262 4722 9322 7651
rect 9630 6490 9690 8467
rect 9814 6765 9874 16627
rect 9995 16284 10061 16285
rect 9995 16220 9996 16284
rect 10060 16220 10061 16284
rect 9995 16219 10061 16220
rect 9998 15197 10058 16219
rect 9995 15196 10061 15197
rect 9995 15132 9996 15196
rect 10060 15132 10061 15196
rect 9995 15131 10061 15132
rect 9995 14652 10061 14653
rect 9995 14588 9996 14652
rect 10060 14588 10061 14652
rect 9995 14587 10061 14588
rect 9998 11797 10058 14587
rect 10182 14245 10242 16763
rect 10366 15469 10426 17443
rect 10547 16964 10613 16965
rect 10547 16900 10548 16964
rect 10612 16900 10613 16964
rect 10547 16899 10613 16900
rect 10363 15468 10429 15469
rect 10363 15404 10364 15468
rect 10428 15404 10429 15468
rect 10363 15403 10429 15404
rect 10363 15196 10429 15197
rect 10363 15132 10364 15196
rect 10428 15132 10429 15196
rect 10363 15131 10429 15132
rect 10366 14925 10426 15131
rect 10363 14924 10429 14925
rect 10363 14860 10364 14924
rect 10428 14860 10429 14924
rect 10363 14859 10429 14860
rect 10363 14380 10429 14381
rect 10363 14316 10364 14380
rect 10428 14316 10429 14380
rect 10363 14315 10429 14316
rect 10179 14244 10245 14245
rect 10179 14180 10180 14244
rect 10244 14180 10245 14244
rect 10179 14179 10245 14180
rect 10179 13836 10245 13837
rect 10179 13772 10180 13836
rect 10244 13772 10245 13836
rect 10179 13771 10245 13772
rect 10182 13021 10242 13771
rect 10179 13020 10245 13021
rect 10179 12956 10180 13020
rect 10244 12956 10245 13020
rect 10179 12955 10245 12956
rect 10179 12204 10245 12205
rect 10179 12140 10180 12204
rect 10244 12140 10245 12204
rect 10179 12139 10245 12140
rect 9995 11796 10061 11797
rect 9995 11732 9996 11796
rect 10060 11732 10061 11796
rect 9995 11731 10061 11732
rect 9995 11116 10061 11117
rect 9995 11052 9996 11116
rect 10060 11052 10061 11116
rect 9995 11051 10061 11052
rect 9998 8669 10058 11051
rect 10182 9349 10242 12139
rect 10179 9348 10245 9349
rect 10179 9284 10180 9348
rect 10244 9284 10245 9348
rect 10179 9283 10245 9284
rect 9995 8668 10061 8669
rect 9995 8604 9996 8668
rect 10060 8604 10061 8668
rect 9995 8603 10061 8604
rect 9811 6764 9877 6765
rect 9811 6700 9812 6764
rect 9876 6700 9877 6764
rect 9811 6699 9877 6700
rect 9811 6492 9877 6493
rect 9811 6490 9812 6492
rect 9630 6430 9812 6490
rect 9811 6428 9812 6430
rect 9876 6428 9877 6492
rect 9811 6427 9877 6428
rect 9627 5404 9693 5405
rect 9627 5340 9628 5404
rect 9692 5340 9693 5404
rect 9627 5339 9693 5340
rect 9630 5133 9690 5339
rect 9627 5132 9693 5133
rect 9627 5068 9628 5132
rect 9692 5068 9693 5132
rect 9627 5067 9693 5068
rect 9627 4860 9693 4861
rect 9627 4796 9628 4860
rect 9692 4796 9693 4860
rect 9627 4795 9693 4796
rect 9078 4662 9322 4722
rect 9078 4317 9138 4662
rect 9259 4452 9325 4453
rect 9259 4388 9260 4452
rect 9324 4388 9325 4452
rect 9259 4387 9325 4388
rect 9075 4316 9141 4317
rect 9075 4252 9076 4316
rect 9140 4252 9141 4316
rect 9075 4251 9141 4252
rect 9075 3228 9141 3229
rect 9075 3164 9076 3228
rect 9140 3164 9141 3228
rect 9075 3163 9141 3164
rect 8891 2820 8957 2821
rect 8891 2756 8892 2820
rect 8956 2756 8957 2820
rect 8891 2755 8957 2756
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 9078 1461 9138 3163
rect 9262 2277 9322 4387
rect 9630 2821 9690 4795
rect 9814 3773 9874 6427
rect 9811 3772 9877 3773
rect 9811 3708 9812 3772
rect 9876 3708 9877 3772
rect 9811 3707 9877 3708
rect 9627 2820 9693 2821
rect 9627 2756 9628 2820
rect 9692 2756 9693 2820
rect 9627 2755 9693 2756
rect 9259 2276 9325 2277
rect 9259 2212 9260 2276
rect 9324 2212 9325 2276
rect 9259 2211 9325 2212
rect 9075 1460 9141 1461
rect 9075 1396 9076 1460
rect 9140 1396 9141 1460
rect 9075 1395 9141 1396
rect 6315 1188 6381 1189
rect 6315 1124 6316 1188
rect 6380 1124 6381 1188
rect 6315 1123 6381 1124
rect 7971 1188 8037 1189
rect 7971 1124 7972 1188
rect 8036 1124 8037 1188
rect 7971 1123 8037 1124
rect 9998 1053 10058 8603
rect 10182 4997 10242 9283
rect 10179 4996 10245 4997
rect 10179 4932 10180 4996
rect 10244 4932 10245 4996
rect 10179 4931 10245 4932
rect 10179 4860 10245 4861
rect 10179 4796 10180 4860
rect 10244 4796 10245 4860
rect 10179 4795 10245 4796
rect 10182 2685 10242 4795
rect 10366 4181 10426 14315
rect 10550 14245 10610 16899
rect 10805 16896 11125 17456
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 15808 11125 16832
rect 13270 17440 13590 17456
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 13270 16352 13590 17376
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 12939 16284 13005 16285
rect 12939 16220 12940 16284
rect 13004 16220 13005 16284
rect 12939 16219 13005 16220
rect 11651 15876 11717 15877
rect 11651 15812 11652 15876
rect 11716 15812 11717 15876
rect 11651 15811 11717 15812
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 14720 11125 15744
rect 11283 15740 11349 15741
rect 11283 15676 11284 15740
rect 11348 15676 11349 15740
rect 11283 15675 11349 15676
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10547 14244 10613 14245
rect 10547 14180 10548 14244
rect 10612 14180 10613 14244
rect 10547 14179 10613 14180
rect 10805 13632 11125 14656
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10547 13020 10613 13021
rect 10547 12956 10548 13020
rect 10612 12956 10613 13020
rect 10547 12955 10613 12956
rect 10550 12613 10610 12955
rect 10547 12612 10613 12613
rect 10547 12548 10548 12612
rect 10612 12548 10613 12612
rect 10547 12547 10613 12548
rect 10805 12544 11125 13568
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 11456 11125 12480
rect 11286 12205 11346 15675
rect 11283 12204 11349 12205
rect 11283 12140 11284 12204
rect 11348 12140 11349 12204
rect 11283 12139 11349 12140
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 10368 11125 11392
rect 11283 11388 11349 11389
rect 11283 11324 11284 11388
rect 11348 11324 11349 11388
rect 11283 11323 11349 11324
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10547 10164 10613 10165
rect 10547 10100 10548 10164
rect 10612 10100 10613 10164
rect 10547 10099 10613 10100
rect 10363 4180 10429 4181
rect 10363 4116 10364 4180
rect 10428 4116 10429 4180
rect 10363 4115 10429 4116
rect 10179 2684 10245 2685
rect 10179 2620 10180 2684
rect 10244 2620 10245 2684
rect 10179 2619 10245 2620
rect 10366 1461 10426 4115
rect 10550 2821 10610 10099
rect 10805 9280 11125 10304
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 8192 11125 9216
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 7104 11125 8128
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 6016 11125 7040
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 3840 11125 4864
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10547 2820 10613 2821
rect 10547 2756 10548 2820
rect 10612 2756 10613 2820
rect 10547 2755 10613 2756
rect 10805 2752 11125 3776
rect 11286 3229 11346 11323
rect 11654 9757 11714 15811
rect 12755 15332 12821 15333
rect 12755 15268 12756 15332
rect 12820 15268 12821 15332
rect 12755 15267 12821 15268
rect 12203 15196 12269 15197
rect 12203 15132 12204 15196
rect 12268 15132 12269 15196
rect 12203 15131 12269 15132
rect 11835 13564 11901 13565
rect 11835 13500 11836 13564
rect 11900 13500 11901 13564
rect 11835 13499 11901 13500
rect 11467 9756 11533 9757
rect 11467 9692 11468 9756
rect 11532 9692 11533 9756
rect 11467 9691 11533 9692
rect 11651 9756 11717 9757
rect 11651 9692 11652 9756
rect 11716 9692 11717 9756
rect 11651 9691 11717 9692
rect 11470 4045 11530 9691
rect 11651 8668 11717 8669
rect 11651 8604 11652 8668
rect 11716 8604 11717 8668
rect 11651 8603 11717 8604
rect 11654 6901 11714 8603
rect 11838 8125 11898 13499
rect 12019 12204 12085 12205
rect 12019 12140 12020 12204
rect 12084 12140 12085 12204
rect 12019 12139 12085 12140
rect 12022 10437 12082 12139
rect 12019 10436 12085 10437
rect 12019 10372 12020 10436
rect 12084 10372 12085 10436
rect 12019 10371 12085 10372
rect 12019 8668 12085 8669
rect 12019 8604 12020 8668
rect 12084 8604 12085 8668
rect 12019 8603 12085 8604
rect 11835 8124 11901 8125
rect 11835 8060 11836 8124
rect 11900 8060 11901 8124
rect 11835 8059 11901 8060
rect 11835 7988 11901 7989
rect 11835 7924 11836 7988
rect 11900 7924 11901 7988
rect 11835 7923 11901 7924
rect 11651 6900 11717 6901
rect 11651 6836 11652 6900
rect 11716 6836 11717 6900
rect 11651 6835 11717 6836
rect 11838 5949 11898 7923
rect 11835 5948 11901 5949
rect 11835 5884 11836 5948
rect 11900 5884 11901 5948
rect 11835 5883 11901 5884
rect 11651 5540 11717 5541
rect 11651 5476 11652 5540
rect 11716 5476 11717 5540
rect 11651 5475 11717 5476
rect 11467 4044 11533 4045
rect 11467 3980 11468 4044
rect 11532 3980 11533 4044
rect 11467 3979 11533 3980
rect 11467 3908 11533 3909
rect 11467 3844 11468 3908
rect 11532 3844 11533 3908
rect 11467 3843 11533 3844
rect 11470 3229 11530 3843
rect 11283 3228 11349 3229
rect 11283 3164 11284 3228
rect 11348 3164 11349 3228
rect 11283 3163 11349 3164
rect 11467 3228 11533 3229
rect 11467 3164 11468 3228
rect 11532 3164 11533 3228
rect 11467 3163 11533 3164
rect 11467 2820 11533 2821
rect 11467 2756 11468 2820
rect 11532 2756 11533 2820
rect 11467 2755 11533 2756
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2128 11125 2688
rect 11470 2277 11530 2755
rect 11467 2276 11533 2277
rect 11467 2212 11468 2276
rect 11532 2212 11533 2276
rect 11467 2211 11533 2212
rect 11654 1597 11714 5475
rect 11838 2821 11898 5883
rect 12022 4317 12082 8603
rect 12206 5677 12266 15131
rect 12387 13836 12453 13837
rect 12387 13772 12388 13836
rect 12452 13772 12453 13836
rect 12387 13771 12453 13772
rect 12390 10165 12450 13771
rect 12571 12476 12637 12477
rect 12571 12412 12572 12476
rect 12636 12412 12637 12476
rect 12571 12411 12637 12412
rect 12387 10164 12453 10165
rect 12387 10100 12388 10164
rect 12452 10100 12453 10164
rect 12387 10099 12453 10100
rect 12387 8804 12453 8805
rect 12387 8740 12388 8804
rect 12452 8740 12453 8804
rect 12387 8739 12453 8740
rect 12203 5676 12269 5677
rect 12203 5612 12204 5676
rect 12268 5612 12269 5676
rect 12203 5611 12269 5612
rect 12203 5540 12269 5541
rect 12203 5476 12204 5540
rect 12268 5476 12269 5540
rect 12203 5475 12269 5476
rect 12019 4316 12085 4317
rect 12019 4252 12020 4316
rect 12084 4252 12085 4316
rect 12019 4251 12085 4252
rect 12019 3908 12085 3909
rect 12019 3844 12020 3908
rect 12084 3844 12085 3908
rect 12019 3843 12085 3844
rect 12022 3093 12082 3843
rect 12206 3773 12266 5475
rect 12203 3772 12269 3773
rect 12203 3708 12204 3772
rect 12268 3708 12269 3772
rect 12203 3707 12269 3708
rect 12019 3092 12085 3093
rect 12019 3028 12020 3092
rect 12084 3028 12085 3092
rect 12019 3027 12085 3028
rect 11835 2820 11901 2821
rect 11835 2756 11836 2820
rect 11900 2756 11901 2820
rect 11835 2755 11901 2756
rect 12206 2141 12266 3707
rect 12390 3229 12450 8739
rect 12574 7853 12634 12411
rect 12571 7852 12637 7853
rect 12571 7788 12572 7852
rect 12636 7788 12637 7852
rect 12571 7787 12637 7788
rect 12571 7036 12637 7037
rect 12571 6972 12572 7036
rect 12636 6972 12637 7036
rect 12571 6971 12637 6972
rect 12574 5949 12634 6971
rect 12571 5948 12637 5949
rect 12571 5884 12572 5948
rect 12636 5884 12637 5948
rect 12571 5883 12637 5884
rect 12571 4996 12637 4997
rect 12571 4932 12572 4996
rect 12636 4932 12637 4996
rect 12571 4931 12637 4932
rect 12574 3637 12634 4931
rect 12571 3636 12637 3637
rect 12571 3572 12572 3636
rect 12636 3572 12637 3636
rect 12571 3571 12637 3572
rect 12387 3228 12453 3229
rect 12387 3164 12388 3228
rect 12452 3164 12453 3228
rect 12387 3163 12453 3164
rect 12758 2685 12818 15267
rect 12942 14517 13002 16219
rect 13270 15264 13590 16288
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 12939 14516 13005 14517
rect 12939 14452 12940 14516
rect 13004 14452 13005 14516
rect 12939 14451 13005 14452
rect 12942 5949 13002 14451
rect 13270 14176 13590 15200
rect 13859 14788 13925 14789
rect 13859 14724 13860 14788
rect 13924 14724 13925 14788
rect 13859 14723 13925 14724
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 13088 13590 14112
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 12000 13590 13024
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13123 11932 13189 11933
rect 13123 11868 13124 11932
rect 13188 11868 13189 11932
rect 13123 11867 13189 11868
rect 13126 7309 13186 11867
rect 13270 10912 13590 11936
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 9824 13590 10848
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 8736 13590 9760
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 7648 13590 8672
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13123 7308 13189 7309
rect 13123 7244 13124 7308
rect 13188 7244 13189 7308
rect 13123 7243 13189 7244
rect 13270 6560 13590 7584
rect 13675 6900 13741 6901
rect 13675 6836 13676 6900
rect 13740 6836 13741 6900
rect 13675 6835 13741 6836
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 12939 5948 13005 5949
rect 12939 5884 12940 5948
rect 13004 5946 13005 5948
rect 13004 5886 13186 5946
rect 13004 5884 13005 5886
rect 12939 5883 13005 5884
rect 12939 4724 13005 4725
rect 12939 4660 12940 4724
rect 13004 4660 13005 4724
rect 12939 4659 13005 4660
rect 12755 2684 12821 2685
rect 12755 2620 12756 2684
rect 12820 2620 12821 2684
rect 12755 2619 12821 2620
rect 12203 2140 12269 2141
rect 12203 2076 12204 2140
rect 12268 2076 12269 2140
rect 12203 2075 12269 2076
rect 11651 1596 11717 1597
rect 11651 1532 11652 1596
rect 11716 1532 11717 1596
rect 11651 1531 11717 1532
rect 10363 1460 10429 1461
rect 10363 1396 10364 1460
rect 10428 1396 10429 1460
rect 10363 1395 10429 1396
rect 12942 1325 13002 4659
rect 13126 3637 13186 5886
rect 13270 5472 13590 6496
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13123 3636 13189 3637
rect 13123 3572 13124 3636
rect 13188 3572 13189 3636
rect 13123 3571 13189 3572
rect 13270 3296 13590 4320
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 2208 13590 3232
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2128 13590 2144
rect 12939 1324 13005 1325
rect 12939 1260 12940 1324
rect 13004 1260 13005 1324
rect 12939 1259 13005 1260
rect 13678 1189 13738 6835
rect 13862 6357 13922 14723
rect 14411 9620 14477 9621
rect 14411 9556 14412 9620
rect 14476 9556 14477 9620
rect 14411 9555 14477 9556
rect 14227 9212 14293 9213
rect 14227 9148 14228 9212
rect 14292 9148 14293 9212
rect 14227 9147 14293 9148
rect 14043 7172 14109 7173
rect 14043 7108 14044 7172
rect 14108 7108 14109 7172
rect 14043 7107 14109 7108
rect 13859 6356 13925 6357
rect 13859 6292 13860 6356
rect 13924 6292 13925 6356
rect 13859 6291 13925 6292
rect 13862 2277 13922 6291
rect 14046 2685 14106 7107
rect 14230 4589 14290 9147
rect 14227 4588 14293 4589
rect 14227 4524 14228 4588
rect 14292 4524 14293 4588
rect 14227 4523 14293 4524
rect 14414 3229 14474 9555
rect 14411 3228 14477 3229
rect 14411 3164 14412 3228
rect 14476 3164 14477 3228
rect 14411 3163 14477 3164
rect 14043 2684 14109 2685
rect 14043 2620 14044 2684
rect 14108 2620 14109 2684
rect 14043 2619 14109 2620
rect 13859 2276 13925 2277
rect 13859 2212 13860 2276
rect 13924 2212 13925 2276
rect 13859 2211 13925 2212
rect 13675 1188 13741 1189
rect 13675 1124 13676 1188
rect 13740 1124 13741 1188
rect 13675 1123 13741 1124
rect 9995 1052 10061 1053
rect 9995 988 9996 1052
rect 10060 988 10061 1052
rect 9995 987 10061 988
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2852 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2852 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4232 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4324 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28
timestamp 1606256979
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 5428 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5520 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5060 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1606256979
transform 1 0 5152 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1606256979
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8188 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7636 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1606256979
transform 1 0 7728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 8096 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_80
timestamp 1606256979
transform 1 0 8464 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_87
timestamp 1606256979
transform 1 0 9108 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1606256979
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9016 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 8832 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 9200 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1606256979
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 10396 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _53_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10028 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1606256979
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1606256979
transform 1 0 11224 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1606256979
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp 1606256979
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14076 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14260 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1606256979
transform 1 0 13248 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1606256979
transform 1 0 13432 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1606256979
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1606256979
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_151
timestamp 1606256979
transform 1 0 14996 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2852 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2668 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_12
timestamp 1606256979
transform 1 0 2208 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_16
timestamp 1606256979
transform 1 0 2576 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1606256979
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1606256979
transform 1 0 4876 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 4968 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6164 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1606256979
transform 1 0 5796 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 7360 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8188 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_64
timestamp 1606256979
transform 1 0 6992 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 9016 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1606256979
transform 1 0 10488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606256979
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 10856 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12052 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1606256979
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13248 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1606256979
transform 1 0 12880 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1606256979
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1606256979
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2576 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 1564 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_14
timestamp 1606256979
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 4876 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4048 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5520 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_47
timestamp 1606256979
transform 1 0 5428 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1606256979
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1606256979
transform 1 0 8004 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1606256979
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 10396 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 8832 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 10028 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_93
timestamp 1606256979
transform 1 0 9660 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_100
timestamp 1606256979
transform 1 0 10304 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1606256979
transform 1 0 11224 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1606256979
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13616 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1606256979
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1606256979
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1606256979
transform 1 0 14444 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1606256979
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_153
timestamp 1606256979
transform 1 0 15180 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 2852 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1606256979
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1606256979
transform 1 0 4876 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6440 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 5244 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_54
timestamp 1606256979
transform 1 0 6072 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8280 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_74
timestamp 1606256979
transform 1 0 7912 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1606256979
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1606256979
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1606256979
transform 1 0 10488 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606256979
transform 1 0 11684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10856 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1606256979
transform 1 0 14444 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13248 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp 1606256979
transform 1 0 12880 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1606256979
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1606256979
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2484 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_12
timestamp 1606256979
transform 1 0 2208 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1606256979
transform 1 0 3312 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4876 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 3680 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1606256979
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1606256979
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_62
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7360 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1606256979
transform 1 0 9200 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10396 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_84
timestamp 1606256979
transform 1 0 8832 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_97
timestamp 1606256979
transform 1 0 10028 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11224 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp 1606256979
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13616 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1606256979
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1606256979
transform 1 0 14444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1606256979
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_153
timestamp 1606256979
transform 1 0 15180 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2760 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 1840 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2208 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1606256979
transform 1 0 1748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1606256979
transform 1 0 2668 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4876 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 3036 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4508 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606256979
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 1606256979
transform 1 0 4416 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1606256979
transform 1 0 4508 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 5704 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_46
timestamp 1606256979
transform 1 0 5336 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1606256979
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7636 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8648 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_66
timestamp 1606256979
transform 1 0 7176 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_70
timestamp 1606256979
transform 1 0 7544 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1606256979
transform 1 0 8280 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1606256979
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1606256979
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1606256979
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_102
timestamp 1606256979
transform 1 0 10488 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1606256979
transform 1 0 10120 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _21_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10856 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12052 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_115
timestamp 1606256979
transform 1 0 11684 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_111
timestamp 1606256979
transform 1 0 11316 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1606256979
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1606256979
transform 1 0 14444 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13248 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13616 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1606256979
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_128
timestamp 1606256979
transform 1 0 12880 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1606256979
transform 1 0 14076 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_134
timestamp 1606256979
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1606256979
transform 1 0 14444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1606256979
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1606256979
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1606256979
transform 1 0 15180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2116 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1606256979
transform 1 0 1748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1606256979
transform 1 0 4508 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606256979
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1606256979
transform 1 0 4416 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5796 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_46
timestamp 1606256979
transform 1 0 5336 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_50
timestamp 1606256979
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 7636 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_67
timestamp 1606256979
transform 1 0 7268 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1606256979
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1606256979
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_102
timestamp 1606256979
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10856 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1606256979
transform 1 0 12052 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_115
timestamp 1606256979
transform 1 0 11684 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1606256979
transform 1 0 14444 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1606256979
transform 1 0 13248 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1606256979
transform 1 0 12880 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1606256979
transform 1 0 14076 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1606256979
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1840 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1606256979
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_17
timestamp 1606256979
transform 1 0 2668 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4876 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 3036 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_37
timestamp 1606256979
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1606256979
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1606256979
transform 1 0 8280 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8648 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_81
timestamp 1606256979
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1606256979
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1606256979
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1606256979
transform 1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_111
timestamp 1606256979
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1606256979
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13616 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1606256979
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_145
timestamp 1606256979
transform 1 0 14444 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1606256979
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1606256979
transform 1 0 15180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2116 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1606256979
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1606256979
transform 1 0 4508 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606256979
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_36
timestamp 1606256979
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5704 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_46
timestamp 1606256979
transform 1 0 5336 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1606256979
transform 1 0 8004 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 8280 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1606256979
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_66
timestamp 1606256979
transform 1 0 7176 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_72
timestamp 1606256979
transform 1 0 7728 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1606256979
transform 1 0 9108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606256979
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1606256979
transform 1 0 11500 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_109
timestamp 1606256979
transform 1 0 11132 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_122
timestamp 1606256979
transform 1 0 12328 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12696 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13892 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1606256979
transform 1 0 13524 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp 1606256979
transform 1 0 14720 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1606256979
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 1564 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 2760 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_14
timestamp 1606256979
transform 1 0 2392 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4876 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3036 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_37
timestamp 1606256979
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1606256979
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8648 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_78
timestamp 1606256979
transform 1 0 8280 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10488 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_98
timestamp 1606256979
transform 1 0 10120 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1606256979
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1606256979
transform 1 0 13616 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp 1606256979
transform 1 0 13248 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_145
timestamp 1606256979
transform 1 0 14444 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1606256979
transform 1 0 14812 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1606256979
transform 1 0 15180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2116 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_7
timestamp 1606256979
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4232 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1606256979
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5704 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7544 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_66
timestamp 1606256979
transform 1 0 7176 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_86
timestamp 1606256979
transform 1 0 9016 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11500 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_109
timestamp 1606256979
transform 1 0 11132 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13340 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_129
timestamp 1606256979
transform 1 0 12972 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_142
timestamp 1606256979
transform 1 0 14168 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1606256979
transform 1 0 14536 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1606256979
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2116 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1606256979
transform 1 0 1840 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1606256979
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_17
timestamp 1606256979
transform 1 0 2668 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_7
timestamp 1606256979
transform 1 0 1748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 3036 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_37
timestamp 1606256979
transform 1 0 4508 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_41
timestamp 1606256979
transform 1 0 4876 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606256979
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5888 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5244 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 4968 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_48
timestamp 1606256979
transform 1 0 5520 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7728 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7176 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_14_68
timestamp 1606256979
transform 1 0 7360 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10488 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 9016 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1606256979
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11500 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1606256979
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1606256979
transform 1 0 11132 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_122
timestamp 1606256979
transform 1 0 12328 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13892 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13616 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1606256979
transform 1 0 12696 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1606256979
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1606256979
transform 1 0 14444 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1606256979
transform 1 0 13524 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1606256979
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1606256979
transform 1 0 15180 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1606256979
transform 1 0 14720 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1606256979
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1840 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1606256979
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_17
timestamp 1606256979
transform 1 0 2668 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4876 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3036 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_37
timestamp 1606256979
transform 1 0 4508 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1606256979
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8648 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp 1606256979
transform 1 0 8280 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10488 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_98
timestamp 1606256979
transform 1 0 10120 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1606256979
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13616 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1606256979
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_145
timestamp 1606256979
transform 1 0 14444 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1606256979
transform 1 0 14812 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1606256979
transform 1 0 15180 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2116 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606256979
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1606256979
transform 1 0 6256 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 5888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_48
timestamp 1606256979
transform 1 0 5520 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_55
timestamp 1606256979
transform 1 0 6164 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_59
timestamp 1606256979
transform 1 0 6532 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1606256979
transform 1 0 8740 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6900 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1606256979
transform 1 0 8372 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_86
timestamp 1606256979
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1606256979
transform 1 0 11500 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1606256979
transform 1 0 11132 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_122
timestamp 1606256979
transform 1 0 12328 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12696 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13892 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1606256979
transform 1 0 13524 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1606256979
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1606256979
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1606256979
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_17
timestamp 1606256979
transform 1 0 2668 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3036 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4876 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_37
timestamp 1606256979
transform 1 0 4508 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1606256979
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8648 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_78
timestamp 1606256979
transform 1 0 8280 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10488 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_98
timestamp 1606256979
transform 1 0 10120 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1606256979
transform 1 0 11684 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_111
timestamp 1606256979
transform 1 0 11316 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1606256979
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1606256979
transform 1 0 13616 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1606256979
transform 1 0 13248 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_145
timestamp 1606256979
transform 1 0 14444 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1606256979
transform 1 0 14812 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1606256979
transform 1 0 15180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1656 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4692 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606256979
transform 1 0 4324 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606256979
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_37
timestamp 1606256979
transform 1 0 4508 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 6532 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_55
timestamp 1606256979
transform 1 0 6164 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_62
timestamp 1606256979
transform 1 0 6808 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1606256979
transform 1 0 7084 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1606256979
transform 1 0 8280 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_74
timestamp 1606256979
transform 1 0 7912 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 10212 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606256979
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1606256979
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1606256979
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_96
timestamp 1606256979
transform 1 0 9936 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1606256979
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1606256979
transform 1 0 10856 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1606256979
transform 1 0 12052 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_115
timestamp 1606256979
transform 1 0 11684 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13248 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_128
timestamp 1606256979
transform 1 0 12880 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1606256979
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1606256979
transform 1 0 1564 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_14
timestamp 1606256979
transform 1 0 2392 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_17
timestamp 1606256979
transform 1 0 2668 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1606256979
transform 1 0 2760 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 3036 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4876 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_37
timestamp 1606256979
transform 1 0 4508 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1606256979
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_38
timestamp 1606256979
transform 1 0 4600 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4968 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6808 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1606256979
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1606256979
transform 1 0 6440 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1606256979
transform 1 0 8372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8648 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 8096 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_71
timestamp 1606256979
transform 1 0 7636 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_75
timestamp 1606256979
transform 1 0 8004 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1606256979
transform 1 0 8648 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_78
timestamp 1606256979
transform 1 0 8280 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1606256979
transform 1 0 9016 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1606256979
transform 1 0 9660 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1606256979
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 10304 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_89
timestamp 1606256979
transform 1 0 9292 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1606256979
transform 1 0 9936 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1606256979
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1606256979
transform 1 0 11500 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 11776 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_112
timestamp 1606256979
transform 1 0 11408 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_119
timestamp 1606256979
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_109
timestamp 1606256979
transform 1 0 11132 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_122
timestamp 1606256979
transform 1 0 12328 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 13616 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13616 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 12696 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1606256979
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_145
timestamp 1606256979
transform 1 0 14444 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_129
timestamp 1606256979
transform 1 0 12972 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_135
timestamp 1606256979
transform 1 0 13524 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1606256979
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2484 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_11
timestamp 1606256979
transform 1 0 2116 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4876 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1606256979
transform 1 0 3680 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_24
timestamp 1606256979
transform 1 0 3312 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_37
timestamp 1606256979
transform 1 0 4508 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1606256979
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8648 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_78
timestamp 1606256979
transform 1 0 8280 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1606256979
transform 1 0 10488 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1606256979
transform 1 0 10120 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 11684 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_111
timestamp 1606256979
transform 1 0 11316 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1606256979
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 13892 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_132
timestamp 1606256979
transform 1 0 13248 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_138
timestamp 1606256979
transform 1 0 13800 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_142
timestamp 1606256979
transform 1 0 14168 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_154
timestamp 1606256979
transform 1 0 15272 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2760 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1564 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_14
timestamp 1606256979
transform 1 0 2392 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1606256979
transform 1 0 4140 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606256979
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 5336 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_42
timestamp 1606256979
transform 1 0 4968 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_62
timestamp 1606256979
transform 1 0 6808 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 7176 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_82
timestamp 1606256979
transform 1 0 8648 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 9016 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1606256979
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1606256979
transform 1 0 10488 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12052 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1606256979
transform 1 0 10856 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_115
timestamp 1606256979
transform 1 0 11684 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1606256979
transform 1 0 13248 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_128
timestamp 1606256979
transform 1 0 12880 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1606256979
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1606256979
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1606256979
transform 1 0 1932 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1606256979
transform 1 0 1380 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_18
timestamp 1606256979
transform 1 0 2760 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4324 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1606256979
transform 1 0 3128 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_31
timestamp 1606256979
transform 1 0 3956 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5520 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_44
timestamp 1606256979
transform 1 0 5152 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1606256979
transform 1 0 6348 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1606256979
transform 1 0 8004 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1606256979
transform 1 0 8648 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_71
timestamp 1606256979
transform 1 0 7636 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_78
timestamp 1606256979
transform 1 0 8280 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9844 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1606256979
transform 1 0 9476 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_104
timestamp 1606256979
transform 1 0 10672 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606256979
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606256979
transform 1 0 11040 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_112 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11408 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1606256979
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606256979
transform 1 0 13892 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606256979
transform 1 0 13156 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_127
timestamp 1606256979
transform 1 0 12788 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_135
timestamp 1606256979
transform 1 0 13524 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_143
timestamp 1606256979
transform 1 0 14260 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1606256979
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1840 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1606256979
transform 1 0 2760 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1606256979
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1606256979
transform 1 0 1748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_14
timestamp 1606256979
transform 1 0 2392 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4140 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1606256979
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_32
timestamp 1606256979
transform 1 0 4048 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1606256979
transform 1 0 5336 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1606256979
transform 1 0 6532 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_42
timestamp 1606256979
transform 1 0 4968 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_55
timestamp 1606256979
transform 1 0 6164 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1606256979
transform 1 0 7728 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_68
timestamp 1606256979
transform 1 0 7360 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_81
timestamp 1606256979
transform 1 0 8556 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1606256979
transform 1 0 8924 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1606256979
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1606256979
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1606256979
transform 1 0 10488 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10856 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12052 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1606256979
transform 1 0 11684 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606256979
transform 1 0 13984 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606256979
transform 1 0 13248 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_128
timestamp 1606256979
transform 1 0 12880 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1606256979
transform 1 0 13616 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_144
timestamp 1606256979
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1606256979
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1606256979
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606256979
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2208 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_7
timestamp 1606256979
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_11
timestamp 1606256979
transform 1 0 2116 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_18
timestamp 1606256979
transform 1 0 2760 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1606256979
transform 1 0 4324 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 3128 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_31
timestamp 1606256979
transform 1 0 3956 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1606256979
transform 1 0 5520 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_44
timestamp 1606256979
transform 1 0 5152 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1606256979
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1606256979
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606256979
transform 1 0 8096 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6900 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_72
timestamp 1606256979
transform 1 0 7728 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_80
timestamp 1606256979
transform 1 0 8464 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9200 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1606256979
transform 1 0 10396 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1606256979
transform 1 0 10028 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606256979
transform 1 0 11592 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_110
timestamp 1606256979
transform 1 0 11224 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1606256979
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606256979
transform 1 0 13616 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606256979
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_134
timestamp 1606256979
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_140
timestamp 1606256979
transform 1 0 13984 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1606256979
transform 1 0 14628 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_146
timestamp 1606256979
transform 1 0 14536 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1606256979
transform 1 0 15180 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1606256979
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1606256979
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1606256979
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1606256979
transform 1 0 2116 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1840 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_14
timestamp 1606256979
transform 1 0 2392 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2760 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2484 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_30
timestamp 1606256979
transform 1 0 3864 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_24
timestamp 1606256979
transform 1 0 3312 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_26_28
timestamp 1606256979
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_21
timestamp 1606256979
transform 1 0 3036 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 3404 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_32
timestamp 1606256979
transform 1 0 4048 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_32
timestamp 1606256979
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4416 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4324 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606256979
transform 1 0 6164 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1606256979
transform 1 0 5612 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_51
timestamp 1606256979
transform 1 0 5796 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_59
timestamp 1606256979
transform 1 0 6532 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1606256979
transform 1 0 5244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_58
timestamp 1606256979
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1606256979
transform 1 0 8096 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6900 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1606256979
transform 1 0 7176 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1606256979
transform 1 0 8372 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_72
timestamp 1606256979
transform 1 0 7728 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_63
timestamp 1606256979
transform 1 0 6900 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_75
timestamp 1606256979
transform 1 0 8004 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_92
timestamp 1606256979
transform 1 0 9568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_88
timestamp 1606256979
transform 1 0 9200 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1606256979
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1606256979
transform 1 0 8924 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_103
timestamp 1606256979
transform 1 0 10580 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_102
timestamp 1606256979
transform 1 0 10488 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1606256979
transform 1 0 9752 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606256979
transform 1 0 10948 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606256979
transform 1 0 10856 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_111
timestamp 1606256979
transform 1 0 11316 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_110
timestamp 1606256979
transform 1 0 11224 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_118
timestamp 1606256979
transform 1 0 11960 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606256979
transform 1 0 11592 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606256979
transform 1 0 11684 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1606256979
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_119
timestamp 1606256979
transform 1 0 12052 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606256979
transform 1 0 12328 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606256979
transform 1 0 12604 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606256979
transform 1 0 13800 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606256979
transform 1 0 13064 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606256979
transform 1 0 13432 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_26_126
timestamp 1606256979
transform 1 0 12696 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_134
timestamp 1606256979
transform 1 0 13432 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_142
timestamp 1606256979
transform 1 0 14168 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_129
timestamp 1606256979
transform 1 0 12972 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_133
timestamp 1606256979
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1606256979
transform 1 0 14536 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 15824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 15824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1606256979
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1606256979
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_147
timestamp 1606256979
transform 1 0 14628 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1606256979
transform 1 0 15456 0 1 16864
box -38 -48 130 592
<< labels >>
rlabel metal2 s 202 19520 258 20000 6 IO_ISOL_N
port 0 nsew default input
rlabel metal3 s 0 1368 480 1488 6 ccff_head
port 1 nsew default input
rlabel metal3 s 16520 1912 17000 2032 6 ccff_tail
port 2 nsew default tristate
rlabel metal2 s 8482 0 8538 480 6 chany_bottom_in[0]
port 3 nsew default input
rlabel metal2 s 12622 0 12678 480 6 chany_bottom_in[10]
port 4 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[11]
port 5 nsew default input
rlabel metal2 s 13450 0 13506 480 6 chany_bottom_in[12]
port 6 nsew default input
rlabel metal2 s 13818 0 13874 480 6 chany_bottom_in[13]
port 7 nsew default input
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_in[14]
port 8 nsew default input
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_in[15]
port 9 nsew default input
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_in[16]
port 10 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_in[17]
port 11 nsew default input
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_in[18]
port 12 nsew default input
rlabel metal2 s 16302 0 16358 480 6 chany_bottom_in[19]
port 13 nsew default input
rlabel metal2 s 8850 0 8906 480 6 chany_bottom_in[1]
port 14 nsew default input
rlabel metal2 s 9310 0 9366 480 6 chany_bottom_in[2]
port 15 nsew default input
rlabel metal2 s 9678 0 9734 480 6 chany_bottom_in[3]
port 16 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[4]
port 17 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[5]
port 18 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[6]
port 19 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[7]
port 20 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[8]
port 21 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_in[9]
port 22 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 23 nsew default tristate
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_out[10]
port 24 nsew default tristate
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_out[11]
port 25 nsew default tristate
rlabel metal2 s 5170 0 5226 480 6 chany_bottom_out[12]
port 26 nsew default tristate
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_out[13]
port 27 nsew default tristate
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_out[14]
port 28 nsew default tristate
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_out[15]
port 29 nsew default tristate
rlabel metal2 s 6826 0 6882 480 6 chany_bottom_out[16]
port 30 nsew default tristate
rlabel metal2 s 7194 0 7250 480 6 chany_bottom_out[17]
port 31 nsew default tristate
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_out[18]
port 32 nsew default tristate
rlabel metal2 s 8022 0 8078 480 6 chany_bottom_out[19]
port 33 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 34 nsew default tristate
rlabel metal2 s 1030 0 1086 480 6 chany_bottom_out[2]
port 35 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 36 nsew default tristate
rlabel metal2 s 1858 0 1914 480 6 chany_bottom_out[4]
port 37 nsew default tristate
rlabel metal2 s 2226 0 2282 480 6 chany_bottom_out[5]
port 38 nsew default tristate
rlabel metal2 s 2686 0 2742 480 6 chany_bottom_out[6]
port 39 nsew default tristate
rlabel metal2 s 3054 0 3110 480 6 chany_bottom_out[7]
port 40 nsew default tristate
rlabel metal2 s 3514 0 3570 480 6 chany_bottom_out[8]
port 41 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 chany_bottom_out[9]
port 42 nsew default tristate
rlabel metal2 s 8666 19520 8722 20000 6 chany_top_in[0]
port 43 nsew default input
rlabel metal2 s 12714 19520 12770 20000 6 chany_top_in[10]
port 44 nsew default input
rlabel metal2 s 13082 19520 13138 20000 6 chany_top_in[11]
port 45 nsew default input
rlabel metal2 s 13542 19520 13598 20000 6 chany_top_in[12]
port 46 nsew default input
rlabel metal2 s 13910 19520 13966 20000 6 chany_top_in[13]
port 47 nsew default input
rlabel metal2 s 14370 19520 14426 20000 6 chany_top_in[14]
port 48 nsew default input
rlabel metal2 s 14738 19520 14794 20000 6 chany_top_in[15]
port 49 nsew default input
rlabel metal2 s 15106 19520 15162 20000 6 chany_top_in[16]
port 50 nsew default input
rlabel metal2 s 15566 19520 15622 20000 6 chany_top_in[17]
port 51 nsew default input
rlabel metal2 s 15934 19520 15990 20000 6 chany_top_in[18]
port 52 nsew default input
rlabel metal2 s 16394 19520 16450 20000 6 chany_top_in[19]
port 53 nsew default input
rlabel metal2 s 9034 19520 9090 20000 6 chany_top_in[1]
port 54 nsew default input
rlabel metal2 s 9494 19520 9550 20000 6 chany_top_in[2]
port 55 nsew default input
rlabel metal2 s 9862 19520 9918 20000 6 chany_top_in[3]
port 56 nsew default input
rlabel metal2 s 10322 19520 10378 20000 6 chany_top_in[4]
port 57 nsew default input
rlabel metal2 s 10690 19520 10746 20000 6 chany_top_in[5]
port 58 nsew default input
rlabel metal2 s 11058 19520 11114 20000 6 chany_top_in[6]
port 59 nsew default input
rlabel metal2 s 11518 19520 11574 20000 6 chany_top_in[7]
port 60 nsew default input
rlabel metal2 s 11886 19520 11942 20000 6 chany_top_in[8]
port 61 nsew default input
rlabel metal2 s 12346 19520 12402 20000 6 chany_top_in[9]
port 62 nsew default input
rlabel metal2 s 570 19520 626 20000 6 chany_top_out[0]
port 63 nsew default tristate
rlabel metal2 s 4618 19520 4674 20000 6 chany_top_out[10]
port 64 nsew default tristate
rlabel metal2 s 4986 19520 5042 20000 6 chany_top_out[11]
port 65 nsew default tristate
rlabel metal2 s 5446 19520 5502 20000 6 chany_top_out[12]
port 66 nsew default tristate
rlabel metal2 s 5814 19520 5870 20000 6 chany_top_out[13]
port 67 nsew default tristate
rlabel metal2 s 6274 19520 6330 20000 6 chany_top_out[14]
port 68 nsew default tristate
rlabel metal2 s 6642 19520 6698 20000 6 chany_top_out[15]
port 69 nsew default tristate
rlabel metal2 s 7010 19520 7066 20000 6 chany_top_out[16]
port 70 nsew default tristate
rlabel metal2 s 7470 19520 7526 20000 6 chany_top_out[17]
port 71 nsew default tristate
rlabel metal2 s 7838 19520 7894 20000 6 chany_top_out[18]
port 72 nsew default tristate
rlabel metal2 s 8298 19520 8354 20000 6 chany_top_out[19]
port 73 nsew default tristate
rlabel metal2 s 938 19520 994 20000 6 chany_top_out[1]
port 74 nsew default tristate
rlabel metal2 s 1398 19520 1454 20000 6 chany_top_out[2]
port 75 nsew default tristate
rlabel metal2 s 1766 19520 1822 20000 6 chany_top_out[3]
port 76 nsew default tristate
rlabel metal2 s 2226 19520 2282 20000 6 chany_top_out[4]
port 77 nsew default tristate
rlabel metal2 s 2594 19520 2650 20000 6 chany_top_out[5]
port 78 nsew default tristate
rlabel metal2 s 2962 19520 3018 20000 6 chany_top_out[6]
port 79 nsew default tristate
rlabel metal2 s 3422 19520 3478 20000 6 chany_top_out[7]
port 80 nsew default tristate
rlabel metal2 s 3790 19520 3846 20000 6 chany_top_out[8]
port 81 nsew default tristate
rlabel metal2 s 4250 19520 4306 20000 6 chany_top_out[9]
port 82 nsew default tristate
rlabel metal3 s 16520 9800 17000 9920 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 83 nsew default tristate
rlabel metal3 s 16520 13880 17000 14000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 84 nsew default input
rlabel metal3 s 16520 17824 17000 17944 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 85 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 left_grid_pin_16_
port 86 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 left_grid_pin_17_
port 87 nsew default tristate
rlabel metal3 s 0 5176 480 5296 6 left_grid_pin_18_
port 88 nsew default tristate
rlabel metal3 s 0 6128 480 6248 6 left_grid_pin_19_
port 89 nsew default tristate
rlabel metal3 s 0 7080 480 7200 6 left_grid_pin_20_
port 90 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 left_grid_pin_21_
port 91 nsew default tristate
rlabel metal3 s 0 8984 480 9104 6 left_grid_pin_22_
port 92 nsew default tristate
rlabel metal3 s 0 9936 480 10056 6 left_grid_pin_23_
port 93 nsew default tristate
rlabel metal3 s 0 10888 480 11008 6 left_grid_pin_24_
port 94 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 left_grid_pin_25_
port 95 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 left_grid_pin_26_
port 96 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 left_grid_pin_27_
port 97 nsew default tristate
rlabel metal3 s 0 14696 480 14816 6 left_grid_pin_28_
port 98 nsew default tristate
rlabel metal3 s 0 15648 480 15768 6 left_grid_pin_29_
port 99 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 left_grid_pin_30_
port 100 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 left_grid_pin_31_
port 101 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 left_width_0_height_0__pin_0_
port 102 nsew default input
rlabel metal3 s 0 416 480 536 6 left_width_0_height_0__pin_1_lower
port 103 nsew default tristate
rlabel metal3 s 0 19456 480 19576 6 left_width_0_height_0__pin_1_upper
port 104 nsew default tristate
rlabel metal2 s 16762 19520 16818 20000 6 prog_clk_0_N_out
port 105 nsew default tristate
rlabel metal2 s 16762 0 16818 480 6 prog_clk_0_S_out
port 106 nsew default tristate
rlabel metal3 s 0 2320 480 2440 6 prog_clk_0_W_in
port 107 nsew default input
rlabel metal3 s 16520 5856 17000 5976 6 right_grid_pin_0_
port 108 nsew default tristate
rlabel metal4 s 3409 2128 3729 17456 6 VPWR
port 109 nsew default input
rlabel metal4 s 5875 2128 6195 17456 6 VGND
port 110 nsew default input
<< properties >>
string FIXED_BBOX 0 0 17000 20000
<< end >>
