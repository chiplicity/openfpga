magic
tech sky130A
magscale 1 2
timestamp 1606930816
<< locali >>
rect 19107 18785 19291 18819
rect 19257 18751 19291 18785
rect 4997 18071 5031 18173
rect 5641 17051 5675 17289
rect 5583 17017 5675 17051
rect 18981 15895 19015 16065
rect 12725 15419 12759 15521
rect 8309 14807 8343 15045
rect 2697 14263 2731 14501
rect 16865 14263 16899 14569
rect 10609 13175 10643 13413
rect 17877 12835 17911 12937
rect 3893 12087 3927 12257
rect 8217 12155 8251 12393
rect 11345 12087 11379 12189
rect 17969 12087 18003 12257
rect 7389 11135 7423 11305
rect 8953 11067 8987 11237
rect 17509 11067 17543 11237
rect 7665 10455 7699 10693
rect 18981 10047 19015 10149
rect 13369 9911 13403 10013
rect 17325 9503 17359 9605
rect 19993 9367 20027 9537
rect 9413 8823 9447 8993
rect 13553 8823 13587 9129
rect 15025 8823 15059 8925
rect 17233 8891 17267 9129
rect 18153 8959 18187 9129
rect 6561 8483 6595 8585
rect 8401 8347 8435 8585
rect 18923 8585 19015 8619
rect 9321 8347 9355 8585
rect 18889 8347 18923 8449
rect 18981 8279 19015 8585
rect 21833 8075 21867 17153
rect 2145 7939 2179 8041
rect 13185 7735 13219 7837
rect 15025 7803 15059 8041
rect 14013 7191 14047 7293
rect 18889 7191 18923 7497
rect 18981 7191 19015 7293
rect 8217 6715 8251 6885
rect 10793 6647 10827 6749
rect 19073 6647 19107 6749
rect 5181 6171 5215 6341
rect 7481 6239 7515 6341
rect 9597 6103 9631 6273
rect 16865 6171 16899 6409
rect 19257 6239 19291 6409
rect 7021 5559 7055 5865
rect 8125 5627 8159 5797
rect 6653 5083 6687 5253
rect 10333 5151 10367 5321
rect 13461 5015 13495 5253
rect 10241 4471 10275 4777
rect 12265 4471 12299 4709
rect 16129 4675 16163 4777
rect 3709 4063 3743 4233
rect 6101 4063 6135 4233
rect 4169 3383 4203 3689
rect 12265 3383 12299 3689
rect 12541 2839 12575 3077
rect 15209 2295 15243 2397
<< viali >>
rect 8953 20009 8987 20043
rect 11161 20009 11195 20043
rect 13553 20009 13587 20043
rect 16405 20009 16439 20043
rect 1961 19941 1995 19975
rect 6377 19941 6411 19975
rect 11989 19941 12023 19975
rect 14749 19941 14783 19975
rect 17049 19941 17083 19975
rect 19165 19941 19199 19975
rect 20637 19941 20671 19975
rect 1685 19873 1719 19907
rect 2421 19873 2455 19907
rect 3433 19873 3467 19907
rect 4445 19873 4479 19907
rect 5457 19873 5491 19907
rect 6101 19873 6135 19907
rect 7196 19873 7230 19907
rect 10149 19873 10183 19907
rect 10977 19873 11011 19907
rect 11897 19873 11931 19907
rect 12633 19873 12667 19907
rect 12909 19873 12943 19907
rect 13369 19873 13403 19907
rect 13921 19873 13955 19907
rect 14473 19873 14507 19907
rect 15025 19873 15059 19907
rect 15669 19873 15703 19907
rect 16221 19873 16255 19907
rect 16773 19873 16807 19907
rect 17509 19873 17543 19907
rect 18337 19873 18371 19907
rect 18889 19873 18923 19907
rect 19625 19873 19659 19907
rect 20361 19873 20395 19907
rect 2697 19805 2731 19839
rect 4537 19805 4571 19839
rect 4721 19805 4755 19839
rect 5549 19805 5583 19839
rect 5733 19805 5767 19839
rect 6929 19805 6963 19839
rect 9045 19805 9079 19839
rect 9137 19805 9171 19839
rect 10241 19805 10275 19839
rect 10333 19805 10367 19839
rect 12081 19805 12115 19839
rect 15853 19805 15887 19839
rect 17785 19805 17819 19839
rect 19901 19805 19935 19839
rect 3617 19737 3651 19771
rect 9781 19737 9815 19771
rect 14105 19737 14139 19771
rect 15209 19737 15243 19771
rect 4077 19669 4111 19703
rect 5089 19669 5123 19703
rect 8309 19669 8343 19703
rect 8585 19669 8619 19703
rect 11529 19669 11563 19703
rect 18521 19669 18555 19703
rect 8401 19465 8435 19499
rect 10241 19465 10275 19499
rect 12449 19465 12483 19499
rect 15485 19465 15519 19499
rect 14657 19397 14691 19431
rect 3157 19329 3191 19363
rect 4353 19329 4387 19363
rect 7021 19329 7055 19363
rect 11989 19329 12023 19363
rect 13093 19329 13127 19363
rect 14289 19329 14323 19363
rect 15209 19329 15243 19363
rect 16037 19329 16071 19363
rect 18981 19329 19015 19363
rect 1685 19261 1719 19295
rect 1961 19261 1995 19295
rect 2973 19261 3007 19295
rect 4820 19261 4854 19295
rect 5080 19261 5114 19295
rect 8861 19261 8895 19295
rect 10517 19261 10551 19295
rect 11805 19261 11839 19295
rect 14013 19261 14047 19295
rect 15025 19261 15059 19295
rect 16497 19261 16531 19295
rect 17233 19261 17267 19295
rect 18061 19261 18095 19295
rect 18797 19261 18831 19295
rect 19901 19261 19935 19295
rect 20453 19261 20487 19295
rect 20729 19261 20763 19295
rect 4261 19193 4295 19227
rect 7288 19193 7322 19227
rect 9128 19193 9162 19227
rect 10793 19193 10827 19227
rect 11713 19193 11747 19227
rect 12817 19193 12851 19227
rect 15117 19193 15151 19227
rect 16773 19193 16807 19227
rect 17509 19193 17543 19227
rect 2513 19125 2547 19159
rect 2881 19125 2915 19159
rect 3801 19125 3835 19159
rect 4169 19125 4203 19159
rect 6193 19125 6227 19159
rect 11345 19125 11379 19159
rect 12909 19125 12943 19159
rect 13645 19125 13679 19159
rect 14105 19125 14139 19159
rect 15853 19125 15887 19159
rect 15945 19125 15979 19159
rect 18245 19125 18279 19159
rect 20085 19125 20119 19159
rect 2973 18921 3007 18955
rect 6193 18921 6227 18955
rect 9689 18921 9723 18955
rect 12817 18921 12851 18955
rect 14749 18921 14783 18955
rect 1961 18853 1995 18887
rect 3341 18853 3375 18887
rect 7021 18853 7055 18887
rect 10057 18853 10091 18887
rect 13338 18853 13372 18887
rect 18153 18853 18187 18887
rect 20361 18853 20395 18887
rect 1685 18785 1719 18819
rect 2421 18785 2455 18819
rect 4077 18785 4111 18819
rect 4344 18785 4378 18819
rect 6101 18785 6135 18819
rect 6745 18785 6779 18819
rect 7748 18785 7782 18819
rect 10701 18785 10735 18819
rect 11704 18785 11738 18819
rect 16681 18785 16715 18819
rect 17325 18785 17359 18819
rect 17877 18785 17911 18819
rect 18613 18785 18647 18819
rect 18889 18785 18923 18819
rect 19073 18785 19107 18819
rect 19349 18785 19383 18819
rect 20085 18785 20119 18819
rect 3433 18717 3467 18751
rect 3617 18717 3651 18751
rect 6285 18717 6319 18751
rect 7481 18717 7515 18751
rect 9137 18717 9171 18751
rect 10149 18717 10183 18751
rect 10241 18717 10275 18751
rect 10977 18717 11011 18751
rect 11437 18717 11471 18751
rect 13093 18717 13127 18751
rect 16773 18717 16807 18751
rect 16957 18717 16991 18751
rect 19257 18717 19291 18751
rect 19625 18717 19659 18751
rect 16313 18649 16347 18683
rect 2605 18581 2639 18615
rect 5457 18581 5491 18615
rect 5733 18581 5767 18615
rect 8861 18581 8895 18615
rect 14473 18581 14507 18615
rect 16221 18581 16255 18615
rect 17509 18581 17543 18615
rect 1961 18377 1995 18411
rect 7021 18377 7055 18411
rect 7481 18377 7515 18411
rect 8493 18377 8527 18411
rect 9505 18377 9539 18411
rect 12081 18377 12115 18411
rect 12449 18377 12483 18411
rect 13461 18377 13495 18411
rect 15117 18377 15151 18411
rect 16129 18377 16163 18411
rect 17601 18309 17635 18343
rect 2421 18241 2455 18275
rect 4537 18241 4571 18275
rect 4721 18241 4755 18275
rect 8033 18241 8067 18275
rect 8953 18241 8987 18275
rect 9045 18241 9079 18275
rect 10057 18241 10091 18275
rect 13001 18241 13035 18275
rect 14013 18241 14047 18275
rect 15577 18241 15611 18275
rect 15761 18241 15795 18275
rect 16589 18241 16623 18275
rect 16773 18241 16807 18275
rect 19533 18241 19567 18275
rect 20729 18241 20763 18275
rect 1777 18173 1811 18207
rect 4997 18173 5031 18207
rect 5089 18173 5123 18207
rect 5356 18173 5390 18207
rect 6837 18173 6871 18207
rect 9873 18173 9907 18207
rect 10701 18173 10735 18207
rect 10968 18173 11002 18207
rect 12817 18173 12851 18207
rect 13829 18173 13863 18207
rect 14565 18173 14599 18207
rect 17417 18173 17451 18207
rect 18521 18173 18555 18207
rect 18797 18173 18831 18207
rect 19349 18173 19383 18207
rect 20453 18173 20487 18207
rect 2688 18105 2722 18139
rect 7849 18105 7883 18139
rect 8861 18105 8895 18139
rect 12909 18105 12943 18139
rect 13921 18105 13955 18139
rect 15485 18105 15519 18139
rect 20545 18105 20579 18139
rect 3801 18037 3835 18071
rect 4077 18037 4111 18071
rect 4445 18037 4479 18071
rect 4997 18037 5031 18071
rect 6469 18037 6503 18071
rect 7941 18037 7975 18071
rect 9965 18037 9999 18071
rect 14749 18037 14783 18071
rect 16497 18037 16531 18071
rect 18429 18037 18463 18071
rect 20085 18037 20119 18071
rect 1869 17833 1903 17867
rect 2421 17833 2455 17867
rect 2881 17833 2915 17867
rect 4077 17833 4111 17867
rect 4537 17833 4571 17867
rect 5089 17833 5123 17867
rect 6837 17833 6871 17867
rect 7481 17833 7515 17867
rect 8585 17833 8619 17867
rect 8953 17833 8987 17867
rect 9689 17833 9723 17867
rect 11069 17833 11103 17867
rect 13093 17833 13127 17867
rect 17417 17833 17451 17867
rect 17877 17833 17911 17867
rect 19257 17833 19291 17867
rect 19809 17833 19843 17867
rect 4445 17765 4479 17799
rect 7941 17765 7975 17799
rect 13921 17765 13955 17799
rect 17785 17765 17819 17799
rect 20177 17765 20211 17799
rect 1777 17697 1811 17731
rect 2789 17697 2823 17731
rect 3433 17697 3467 17731
rect 5457 17697 5491 17731
rect 7849 17697 7883 17731
rect 10057 17697 10091 17731
rect 11161 17697 11195 17731
rect 12173 17697 12207 17731
rect 12909 17697 12943 17731
rect 13829 17697 13863 17731
rect 14473 17697 14507 17731
rect 16017 17697 16051 17731
rect 19165 17697 19199 17731
rect 2053 17629 2087 17663
rect 2973 17629 3007 17663
rect 4721 17629 4755 17663
rect 5549 17629 5583 17663
rect 5641 17629 5675 17663
rect 6929 17629 6963 17663
rect 7113 17629 7147 17663
rect 8125 17629 8159 17663
rect 9045 17629 9079 17663
rect 9137 17629 9171 17663
rect 10149 17629 10183 17663
rect 10241 17629 10275 17663
rect 11345 17629 11379 17663
rect 12265 17629 12299 17663
rect 12357 17629 12391 17663
rect 14105 17629 14139 17663
rect 15301 17629 15335 17663
rect 15761 17629 15795 17663
rect 17969 17629 18003 17663
rect 19349 17629 19383 17663
rect 20269 17629 20303 17663
rect 20453 17629 20487 17663
rect 1409 17561 1443 17595
rect 14657 17561 14691 17595
rect 3617 17493 3651 17527
rect 6469 17493 6503 17527
rect 10701 17493 10735 17527
rect 11805 17493 11839 17527
rect 13461 17493 13495 17527
rect 17141 17493 17175 17527
rect 18797 17493 18831 17527
rect 3525 17289 3559 17323
rect 4261 17289 4295 17323
rect 5641 17289 5675 17323
rect 8309 17289 8343 17323
rect 9413 17289 9447 17323
rect 10425 17289 10459 17323
rect 11621 17289 11655 17323
rect 12449 17289 12483 17323
rect 16865 17289 16899 17323
rect 19073 17289 19107 17323
rect 20269 17289 20303 17323
rect 4813 17153 4847 17187
rect 1409 17085 1443 17119
rect 2145 17085 2179 17119
rect 9045 17221 9079 17255
rect 15209 17221 15243 17255
rect 18061 17221 18095 17255
rect 6193 17153 6227 17187
rect 6377 17153 6411 17187
rect 6929 17153 6963 17187
rect 9965 17153 9999 17187
rect 10977 17153 11011 17187
rect 12909 17153 12943 17187
rect 13093 17153 13127 17187
rect 18705 17153 18739 17187
rect 19625 17153 19659 17187
rect 20913 17153 20947 17187
rect 21833 17153 21867 17187
rect 6101 17085 6135 17119
rect 8861 17085 8895 17119
rect 11437 17085 11471 17119
rect 13829 17085 13863 17119
rect 14096 17085 14130 17119
rect 15485 17085 15519 17119
rect 17417 17085 17451 17119
rect 18521 17085 18555 17119
rect 19533 17085 19567 17119
rect 20637 17085 20671 17119
rect 1685 17017 1719 17051
rect 2412 17017 2446 17051
rect 4629 17017 4663 17051
rect 5549 17017 5583 17051
rect 7196 17017 7230 17051
rect 9873 17017 9907 17051
rect 10793 17017 10827 17051
rect 15730 17017 15764 17051
rect 3801 16949 3835 16983
rect 4721 16949 4755 16983
rect 5273 16949 5307 16983
rect 5733 16949 5767 16983
rect 9781 16949 9815 16983
rect 10885 16949 10919 16983
rect 12817 16949 12851 16983
rect 17601 16949 17635 16983
rect 18429 16949 18463 16983
rect 19441 16949 19475 16983
rect 20729 16949 20763 16983
rect 1593 16745 1627 16779
rect 2053 16745 2087 16779
rect 2605 16745 2639 16779
rect 4077 16745 4111 16779
rect 4445 16745 4479 16779
rect 6929 16745 6963 16779
rect 7389 16745 7423 16779
rect 9321 16745 9355 16779
rect 10149 16745 10183 16779
rect 12357 16745 12391 16779
rect 15301 16745 15335 16779
rect 15761 16745 15795 16779
rect 16313 16745 16347 16779
rect 17325 16745 17359 16779
rect 18337 16745 18371 16779
rect 19441 16745 19475 16779
rect 19809 16745 19843 16779
rect 1961 16677 1995 16711
rect 8208 16677 8242 16711
rect 13268 16677 13302 16711
rect 17693 16677 17727 16711
rect 18705 16677 18739 16711
rect 2973 16609 3007 16643
rect 4537 16609 4571 16643
rect 5540 16609 5574 16643
rect 7297 16609 7331 16643
rect 9965 16609 9999 16643
rect 10517 16609 10551 16643
rect 10784 16609 10818 16643
rect 12173 16609 12207 16643
rect 14657 16609 14691 16643
rect 15669 16609 15703 16643
rect 16681 16609 16715 16643
rect 17785 16609 17819 16643
rect 18797 16609 18831 16643
rect 19901 16609 19935 16643
rect 2237 16541 2271 16575
rect 3065 16541 3099 16575
rect 3249 16541 3283 16575
rect 4721 16541 4755 16575
rect 5273 16541 5307 16575
rect 7481 16541 7515 16575
rect 7941 16541 7975 16575
rect 13001 16541 13035 16575
rect 15945 16541 15979 16575
rect 16773 16541 16807 16575
rect 16865 16541 16899 16575
rect 17877 16541 17911 16575
rect 18889 16541 18923 16575
rect 19993 16541 20027 16575
rect 6653 16405 6687 16439
rect 11897 16405 11931 16439
rect 14381 16405 14415 16439
rect 14841 16405 14875 16439
rect 1685 16201 1719 16235
rect 2789 16201 2823 16235
rect 6009 16201 6043 16235
rect 8217 16201 8251 16235
rect 9505 16201 9539 16235
rect 12449 16201 12483 16235
rect 14565 16201 14599 16235
rect 15577 16201 15611 16235
rect 16589 16201 16623 16235
rect 20085 16201 20119 16235
rect 3801 16133 3835 16167
rect 6377 16133 6411 16167
rect 8493 16133 8527 16167
rect 19073 16133 19107 16167
rect 3341 16065 3375 16099
rect 4353 16065 4387 16099
rect 5365 16065 5399 16099
rect 9137 16065 9171 16099
rect 10057 16065 10091 16099
rect 13001 16065 13035 16099
rect 13921 16065 13955 16099
rect 14105 16065 14139 16099
rect 15209 16065 15243 16099
rect 16221 16065 16255 16099
rect 17141 16065 17175 16099
rect 18521 16065 18555 16099
rect 18705 16065 18739 16099
rect 18981 16065 19015 16099
rect 19625 16065 19659 16099
rect 20545 16065 20579 16099
rect 20637 16065 20671 16099
rect 1501 15997 1535 16031
rect 2053 15997 2087 16031
rect 2329 15997 2363 16031
rect 4169 15997 4203 16031
rect 5825 15997 5859 16031
rect 6561 15997 6595 16031
rect 6837 15997 6871 16031
rect 10517 15997 10551 16031
rect 13829 15997 13863 16031
rect 14933 15997 14967 16031
rect 3157 15929 3191 15963
rect 7104 15929 7138 15963
rect 8953 15929 8987 15963
rect 10784 15929 10818 15963
rect 12909 15929 12943 15963
rect 20453 15997 20487 16031
rect 19533 15929 19567 15963
rect 3249 15861 3283 15895
rect 4261 15861 4295 15895
rect 4813 15861 4847 15895
rect 5181 15861 5215 15895
rect 5273 15861 5307 15895
rect 8861 15861 8895 15895
rect 9873 15861 9907 15895
rect 9965 15861 9999 15895
rect 11897 15861 11931 15895
rect 12817 15861 12851 15895
rect 13461 15861 13495 15895
rect 15025 15861 15059 15895
rect 15945 15861 15979 15895
rect 16037 15861 16071 15895
rect 16957 15861 16991 15895
rect 17049 15861 17083 15895
rect 18061 15861 18095 15895
rect 18429 15861 18463 15895
rect 18981 15861 19015 15895
rect 19441 15861 19475 15895
rect 1593 15657 1627 15691
rect 1961 15657 1995 15691
rect 2329 15657 2363 15691
rect 3433 15657 3467 15691
rect 4721 15657 4755 15691
rect 5365 15657 5399 15691
rect 6561 15657 6595 15691
rect 7573 15657 7607 15691
rect 8033 15657 8067 15691
rect 8585 15657 8619 15691
rect 14841 15657 14875 15691
rect 15301 15657 15335 15691
rect 16313 15657 16347 15691
rect 18337 15657 18371 15691
rect 19349 15657 19383 15691
rect 6929 15589 6963 15623
rect 8953 15589 8987 15623
rect 9045 15589 9079 15623
rect 11520 15589 11554 15623
rect 18705 15589 18739 15623
rect 19717 15589 19751 15623
rect 1409 15521 1443 15555
rect 3341 15521 3375 15555
rect 4629 15521 4663 15555
rect 5733 15521 5767 15555
rect 5825 15521 5859 15555
rect 7941 15521 7975 15555
rect 10425 15521 10459 15555
rect 11253 15521 11287 15555
rect 12725 15521 12759 15555
rect 13176 15521 13210 15555
rect 14657 15521 14691 15555
rect 15669 15521 15703 15555
rect 16681 15521 16715 15555
rect 17693 15521 17727 15555
rect 17785 15521 17819 15555
rect 18797 15521 18831 15555
rect 2421 15453 2455 15487
rect 2605 15453 2639 15487
rect 3617 15453 3651 15487
rect 4813 15453 4847 15487
rect 5917 15453 5951 15487
rect 7021 15453 7055 15487
rect 7205 15453 7239 15487
rect 8217 15453 8251 15487
rect 9229 15453 9263 15487
rect 10517 15453 10551 15487
rect 10701 15453 10735 15487
rect 12909 15453 12943 15487
rect 15761 15453 15795 15487
rect 15945 15453 15979 15487
rect 16773 15453 16807 15487
rect 16957 15453 16991 15487
rect 17877 15453 17911 15487
rect 18981 15453 19015 15487
rect 19809 15453 19843 15487
rect 19993 15453 20027 15487
rect 2973 15385 3007 15419
rect 12633 15385 12667 15419
rect 12725 15385 12759 15419
rect 16129 15385 16163 15419
rect 4261 15317 4295 15351
rect 10057 15317 10091 15351
rect 14289 15317 14323 15351
rect 17325 15317 17359 15351
rect 6837 15113 6871 15147
rect 11805 15113 11839 15147
rect 12449 15113 12483 15147
rect 13829 15113 13863 15147
rect 17601 15113 17635 15147
rect 8033 15045 8067 15079
rect 8309 15045 8343 15079
rect 3433 14977 3467 15011
rect 7389 14977 7423 15011
rect 1777 14909 1811 14943
rect 3700 14909 3734 14943
rect 5089 14909 5123 14943
rect 7849 14909 7883 14943
rect 2044 14841 2078 14875
rect 5356 14841 5390 14875
rect 8769 14977 8803 15011
rect 10425 14977 10459 15011
rect 13001 14977 13035 15011
rect 18613 14977 18647 15011
rect 19717 14977 19751 15011
rect 20637 14977 20671 15011
rect 8585 14909 8619 14943
rect 12265 14909 12299 14943
rect 13645 14909 13679 14943
rect 14197 14909 14231 14943
rect 16221 14909 16255 14943
rect 18521 14909 18555 14943
rect 19441 14909 19475 14943
rect 9036 14841 9070 14875
rect 10692 14841 10726 14875
rect 14464 14841 14498 14875
rect 16488 14841 16522 14875
rect 18429 14841 18463 14875
rect 20453 14841 20487 14875
rect 3157 14773 3191 14807
rect 4813 14773 4847 14807
rect 6469 14773 6503 14807
rect 7205 14773 7239 14807
rect 7297 14773 7331 14807
rect 8309 14773 8343 14807
rect 8401 14773 8435 14807
rect 10149 14773 10183 14807
rect 12081 14773 12115 14807
rect 12817 14773 12851 14807
rect 12909 14773 12943 14807
rect 15577 14773 15611 14807
rect 18061 14773 18095 14807
rect 19073 14773 19107 14807
rect 19533 14773 19567 14807
rect 20085 14773 20119 14807
rect 20545 14773 20579 14807
rect 2881 14569 2915 14603
rect 3249 14569 3283 14603
rect 4077 14569 4111 14603
rect 4537 14569 4571 14603
rect 7941 14569 7975 14603
rect 9965 14569 9999 14603
rect 12357 14569 12391 14603
rect 16405 14569 16439 14603
rect 16865 14569 16899 14603
rect 18429 14569 18463 14603
rect 18705 14569 18739 14603
rect 19717 14569 19751 14603
rect 2329 14501 2363 14535
rect 2697 14501 2731 14535
rect 3341 14501 3375 14535
rect 5365 14501 5399 14535
rect 6162 14501 6196 14535
rect 10425 14501 10459 14535
rect 12449 14501 12483 14535
rect 15577 14501 15611 14535
rect 1409 14433 1443 14467
rect 2237 14433 2271 14467
rect 2421 14365 2455 14399
rect 1869 14297 1903 14331
rect 4445 14433 4479 14467
rect 5089 14433 5123 14467
rect 8953 14433 8987 14467
rect 10333 14433 10367 14467
rect 11345 14433 11379 14467
rect 13369 14433 13403 14467
rect 14381 14433 14415 14467
rect 14473 14433 14507 14467
rect 15301 14433 15335 14467
rect 3525 14365 3559 14399
rect 4721 14365 4755 14399
rect 5917 14365 5951 14399
rect 8033 14365 8067 14399
rect 8125 14365 8159 14399
rect 9045 14365 9079 14399
rect 9137 14365 9171 14399
rect 10517 14365 10551 14399
rect 11437 14365 11471 14399
rect 11529 14365 11563 14399
rect 12541 14365 12575 14399
rect 13461 14365 13495 14399
rect 13553 14365 13587 14399
rect 14565 14365 14599 14399
rect 16497 14365 16531 14399
rect 16589 14365 16623 14399
rect 8585 14297 8619 14331
rect 16037 14297 16071 14331
rect 17316 14501 17350 14535
rect 20177 14501 20211 14535
rect 17049 14433 17083 14467
rect 19073 14433 19107 14467
rect 20085 14433 20119 14467
rect 19165 14365 19199 14399
rect 19257 14365 19291 14399
rect 20269 14365 20303 14399
rect 20913 14365 20947 14399
rect 2697 14229 2731 14263
rect 7297 14229 7331 14263
rect 7573 14229 7607 14263
rect 10977 14229 11011 14263
rect 11989 14229 12023 14263
rect 13001 14229 13035 14263
rect 14013 14229 14047 14263
rect 16865 14229 16899 14263
rect 1593 14025 1627 14059
rect 5365 14025 5399 14059
rect 5641 14025 5675 14059
rect 9229 14025 9263 14059
rect 9781 14025 9815 14059
rect 10149 14025 10183 14059
rect 11161 14025 11195 14059
rect 14105 14025 14139 14059
rect 14749 14025 14783 14059
rect 16773 14025 16807 14059
rect 19717 14025 19751 14059
rect 20913 14025 20947 14059
rect 16497 13957 16531 13991
rect 2421 13889 2455 13923
rect 2605 13889 2639 13923
rect 3433 13889 3467 13923
rect 3617 13889 3651 13923
rect 6193 13889 6227 13923
rect 7389 13889 7423 13923
rect 7849 13889 7883 13923
rect 10609 13889 10643 13923
rect 10793 13889 10827 13923
rect 11713 13889 11747 13923
rect 17417 13889 17451 13923
rect 20177 13889 20211 13923
rect 20269 13889 20303 13923
rect 1409 13821 1443 13855
rect 3985 13821 4019 13855
rect 4241 13821 4275 13855
rect 7297 13821 7331 13855
rect 8116 13821 8150 13855
rect 9597 13821 9631 13855
rect 11621 13821 11655 13855
rect 12725 13821 12759 13855
rect 14565 13821 14599 13855
rect 15117 13821 15151 13855
rect 15384 13821 15418 13855
rect 18061 13821 18095 13855
rect 18328 13821 18362 13855
rect 20729 13821 20763 13855
rect 3341 13753 3375 13787
rect 6009 13753 6043 13787
rect 7205 13753 7239 13787
rect 10517 13753 10551 13787
rect 12992 13753 13026 13787
rect 20085 13753 20119 13787
rect 1961 13685 1995 13719
rect 2329 13685 2363 13719
rect 2973 13685 3007 13719
rect 6101 13685 6135 13719
rect 6837 13685 6871 13719
rect 11529 13685 11563 13719
rect 17141 13685 17175 13719
rect 17233 13685 17267 13719
rect 19441 13685 19475 13719
rect 3709 13481 3743 13515
rect 4169 13481 4203 13515
rect 4537 13481 4571 13515
rect 5181 13481 5215 13515
rect 5549 13481 5583 13515
rect 6837 13481 6871 13515
rect 8217 13481 8251 13515
rect 10057 13481 10091 13515
rect 10701 13481 10735 13515
rect 11161 13481 11195 13515
rect 11713 13481 11747 13515
rect 12081 13481 12115 13515
rect 12173 13481 12207 13515
rect 15301 13481 15335 13515
rect 15761 13481 15795 13515
rect 16405 13481 16439 13515
rect 16773 13481 16807 13515
rect 17417 13481 17451 13515
rect 17785 13481 17819 13515
rect 7297 13413 7331 13447
rect 10609 13413 10643 13447
rect 18613 13413 18647 13447
rect 19349 13413 19383 13447
rect 19809 13413 19843 13447
rect 1593 13345 1627 13379
rect 2596 13345 2630 13379
rect 4629 13345 4663 13379
rect 6101 13345 6135 13379
rect 7205 13345 7239 13379
rect 8861 13345 8895 13379
rect 10149 13345 10183 13379
rect 1869 13277 1903 13311
rect 2329 13277 2363 13311
rect 4721 13277 4755 13311
rect 5641 13277 5675 13311
rect 5733 13277 5767 13311
rect 7389 13277 7423 13311
rect 8309 13277 8343 13311
rect 8493 13277 8527 13311
rect 10333 13277 10367 13311
rect 11069 13345 11103 13379
rect 12909 13345 12943 13379
rect 13001 13345 13035 13379
rect 13553 13345 13587 13379
rect 13820 13345 13854 13379
rect 15669 13345 15703 13379
rect 16865 13345 16899 13379
rect 17877 13345 17911 13379
rect 18705 13345 18739 13379
rect 11253 13277 11287 13311
rect 12265 13277 12299 13311
rect 15945 13277 15979 13311
rect 16957 13277 16991 13311
rect 17969 13277 18003 13311
rect 18889 13277 18923 13311
rect 19901 13277 19935 13311
rect 19993 13277 20027 13311
rect 12725 13209 12759 13243
rect 6285 13141 6319 13175
rect 6745 13141 6779 13175
rect 7849 13141 7883 13175
rect 9045 13141 9079 13175
rect 9689 13141 9723 13175
rect 10609 13141 10643 13175
rect 13185 13141 13219 13175
rect 14933 13141 14967 13175
rect 18245 13141 18279 13175
rect 19441 13141 19475 13175
rect 1593 12937 1627 12971
rect 4261 12937 4295 12971
rect 5457 12937 5491 12971
rect 6469 12937 6503 12971
rect 7205 12937 7239 12971
rect 9965 12937 9999 12971
rect 14381 12937 14415 12971
rect 16221 12937 16255 12971
rect 17877 12937 17911 12971
rect 3985 12869 4019 12903
rect 8677 12869 8711 12903
rect 14105 12869 14139 12903
rect 2053 12801 2087 12835
rect 2237 12801 2271 12835
rect 4813 12801 4847 12835
rect 6009 12801 6043 12835
rect 6837 12801 6871 12835
rect 9505 12801 9539 12835
rect 10517 12801 10551 12835
rect 11529 12801 11563 12835
rect 14933 12801 14967 12835
rect 16773 12801 16807 12835
rect 17877 12801 17911 12835
rect 18797 12801 18831 12835
rect 18981 12801 19015 12835
rect 19901 12801 19935 12835
rect 20913 12801 20947 12835
rect 2605 12733 2639 12767
rect 4721 12733 4755 12767
rect 6653 12733 6687 12767
rect 7297 12733 7331 12767
rect 7564 12733 7598 12767
rect 9321 12733 9355 12767
rect 10425 12733 10459 12767
rect 11437 12733 11471 12767
rect 12725 12733 12759 12767
rect 14749 12733 14783 12767
rect 14841 12733 14875 12767
rect 15577 12733 15611 12767
rect 15669 12733 15703 12767
rect 17233 12733 17267 12767
rect 19717 12733 19751 12767
rect 19809 12733 19843 12767
rect 20729 12733 20763 12767
rect 2872 12665 2906 12699
rect 4629 12665 4663 12699
rect 5825 12665 5859 12699
rect 9413 12665 9447 12699
rect 12992 12665 13026 12699
rect 16681 12665 16715 12699
rect 17509 12665 17543 12699
rect 1961 12597 1995 12631
rect 5917 12597 5951 12631
rect 8953 12597 8987 12631
rect 10333 12597 10367 12631
rect 10977 12597 11011 12631
rect 11345 12597 11379 12631
rect 15393 12597 15427 12631
rect 15853 12597 15887 12631
rect 16589 12597 16623 12631
rect 18337 12597 18371 12631
rect 18705 12597 18739 12631
rect 19349 12597 19383 12631
rect 20361 12597 20395 12631
rect 20821 12597 20855 12631
rect 1593 12393 1627 12427
rect 2973 12393 3007 12427
rect 4261 12393 4295 12427
rect 6101 12393 6135 12427
rect 7389 12393 7423 12427
rect 8217 12393 8251 12427
rect 8861 12393 8895 12427
rect 11529 12393 11563 12427
rect 11897 12393 11931 12427
rect 11989 12393 12023 12427
rect 12725 12393 12759 12427
rect 13093 12393 13127 12427
rect 13737 12393 13771 12427
rect 17877 12393 17911 12427
rect 19809 12393 19843 12427
rect 20177 12393 20211 12427
rect 20913 12393 20947 12427
rect 7757 12325 7791 12359
rect 1409 12257 1443 12291
rect 2329 12257 2363 12291
rect 3341 12257 3375 12291
rect 3893 12257 3927 12291
rect 4077 12257 4111 12291
rect 4721 12257 4755 12291
rect 4988 12257 5022 12291
rect 6745 12257 6779 12291
rect 2421 12189 2455 12223
rect 2605 12189 2639 12223
rect 3433 12189 3467 12223
rect 3525 12189 3559 12223
rect 6837 12189 6871 12223
rect 6929 12189 6963 12223
rect 7849 12189 7883 12223
rect 8033 12189 8067 12223
rect 8769 12325 8803 12359
rect 15853 12325 15887 12359
rect 16764 12325 16798 12359
rect 18420 12325 18454 12359
rect 9873 12257 9907 12291
rect 10129 12257 10163 12291
rect 14105 12257 14139 12291
rect 14749 12257 14783 12291
rect 17969 12257 18003 12291
rect 18153 12257 18187 12291
rect 8953 12189 8987 12223
rect 11345 12189 11379 12223
rect 12081 12189 12115 12223
rect 13185 12189 13219 12223
rect 13369 12189 13403 12223
rect 14197 12189 14231 12223
rect 14289 12189 14323 12223
rect 15945 12189 15979 12223
rect 16037 12189 16071 12223
rect 16497 12189 16531 12223
rect 6377 12121 6411 12155
rect 8217 12121 8251 12155
rect 11253 12121 11287 12155
rect 15485 12121 15519 12155
rect 1961 12053 1995 12087
rect 3893 12053 3927 12087
rect 8401 12053 8435 12087
rect 11345 12053 11379 12087
rect 20269 12189 20303 12223
rect 20361 12189 20395 12223
rect 17969 12053 18003 12087
rect 19533 12053 19567 12087
rect 4997 11849 5031 11883
rect 5549 11849 5583 11883
rect 6837 11849 6871 11883
rect 7849 11849 7883 11883
rect 8861 11849 8895 11883
rect 14105 11849 14139 11883
rect 15761 11849 15795 11883
rect 18797 11849 18831 11883
rect 21005 11849 21039 11883
rect 4721 11781 4755 11815
rect 11989 11781 12023 11815
rect 13829 11781 13863 11815
rect 2881 11713 2915 11747
rect 6101 11713 6135 11747
rect 7389 11713 7423 11747
rect 8493 11713 8527 11747
rect 9413 11713 9447 11747
rect 10241 11713 10275 11747
rect 18337 11713 18371 11747
rect 19349 11713 19383 11747
rect 20361 11713 20395 11747
rect 1501 11645 1535 11679
rect 3341 11645 3375 11679
rect 3597 11645 3631 11679
rect 4813 11645 4847 11679
rect 5457 11645 5491 11679
rect 5917 11645 5951 11679
rect 8217 11645 8251 11679
rect 8309 11645 8343 11679
rect 9229 11645 9263 11679
rect 10057 11645 10091 11679
rect 10609 11645 10643 11679
rect 12449 11645 12483 11679
rect 14289 11645 14323 11679
rect 14381 11645 14415 11679
rect 16313 11645 16347 11679
rect 16580 11645 16614 11679
rect 18061 11645 18095 11679
rect 19257 11645 19291 11679
rect 20177 11645 20211 11679
rect 20821 11645 20855 11679
rect 1777 11577 1811 11611
rect 6009 11577 6043 11611
rect 7297 11577 7331 11611
rect 10876 11577 10910 11611
rect 12694 11577 12728 11611
rect 14648 11577 14682 11611
rect 2237 11509 2271 11543
rect 2605 11509 2639 11543
rect 2697 11509 2731 11543
rect 7205 11509 7239 11543
rect 9321 11509 9355 11543
rect 9689 11509 9723 11543
rect 10149 11509 10183 11543
rect 17693 11509 17727 11543
rect 19165 11509 19199 11543
rect 19809 11509 19843 11543
rect 20269 11509 20303 11543
rect 1409 11305 1443 11339
rect 3249 11305 3283 11339
rect 3525 11305 3559 11339
rect 4077 11305 4111 11339
rect 5273 11305 5307 11339
rect 7205 11305 7239 11339
rect 7389 11305 7423 11339
rect 8861 11305 8895 11339
rect 11989 11305 12023 11339
rect 15669 11305 15703 11339
rect 15761 11305 15795 11339
rect 16589 11305 16623 11339
rect 18061 11305 18095 11339
rect 18797 11305 18831 11339
rect 20913 11305 20947 11339
rect 6092 11237 6126 11271
rect 1869 11169 1903 11203
rect 2136 11169 2170 11203
rect 4445 11169 4479 11203
rect 5089 11169 5123 11203
rect 8953 11237 8987 11271
rect 9137 11237 9171 11271
rect 10517 11237 10551 11271
rect 17049 11237 17083 11271
rect 17509 11237 17543 11271
rect 19432 11237 19466 11271
rect 7481 11169 7515 11203
rect 7748 11169 7782 11203
rect 4537 11101 4571 11135
rect 4629 11101 4663 11135
rect 5825 11101 5859 11135
rect 7389 11101 7423 11135
rect 9965 11169 9999 11203
rect 12716 11169 12750 11203
rect 14473 11169 14507 11203
rect 14565 11169 14599 11203
rect 16957 11169 16991 11203
rect 12449 11101 12483 11135
rect 14749 11101 14783 11135
rect 15945 11101 15979 11135
rect 17141 11101 17175 11135
rect 17969 11169 18003 11203
rect 18613 11169 18647 11203
rect 18245 11101 18279 11135
rect 19165 11101 19199 11135
rect 8953 11033 8987 11067
rect 13829 11033 13863 11067
rect 15301 11033 15335 11067
rect 17509 11033 17543 11067
rect 20545 11033 20579 11067
rect 10149 10965 10183 10999
rect 14105 10965 14139 10999
rect 17601 10965 17635 10999
rect 3249 10761 3283 10795
rect 3709 10761 3743 10795
rect 4445 10761 4479 10795
rect 8861 10761 8895 10795
rect 12173 10761 12207 10795
rect 16957 10761 16991 10795
rect 21005 10761 21039 10795
rect 7665 10693 7699 10727
rect 9321 10693 9355 10727
rect 11069 10693 11103 10727
rect 13461 10693 13495 10727
rect 14749 10693 14783 10727
rect 15945 10693 15979 10727
rect 5089 10625 5123 10659
rect 5917 10625 5951 10659
rect 6009 10625 6043 10659
rect 7481 10625 7515 10659
rect 1869 10557 1903 10591
rect 3525 10557 3559 10591
rect 4905 10557 4939 10591
rect 2136 10489 2170 10523
rect 4813 10489 4847 10523
rect 5825 10489 5859 10523
rect 7297 10489 7331 10523
rect 8401 10625 8435 10659
rect 11713 10625 11747 10659
rect 13093 10625 13127 10659
rect 13921 10625 13955 10659
rect 14013 10625 14047 10659
rect 15393 10625 15427 10659
rect 16589 10625 16623 10659
rect 17509 10625 17543 10659
rect 20361 10625 20395 10659
rect 9045 10557 9079 10591
rect 9137 10557 9171 10591
rect 9689 10557 9723 10591
rect 11529 10557 11563 10591
rect 11621 10557 11655 10591
rect 11989 10557 12023 10591
rect 13829 10557 13863 10591
rect 15117 10557 15151 10591
rect 16405 10557 16439 10591
rect 17325 10557 17359 10591
rect 18153 10557 18187 10591
rect 18420 10557 18454 10591
rect 20821 10557 20855 10591
rect 9956 10489 9990 10523
rect 12909 10489 12943 10523
rect 1409 10421 1443 10455
rect 5457 10421 5491 10455
rect 6837 10421 6871 10455
rect 7205 10421 7239 10455
rect 7665 10421 7699 10455
rect 7849 10421 7883 10455
rect 8217 10421 8251 10455
rect 8309 10421 8343 10455
rect 11161 10421 11195 10455
rect 12449 10421 12483 10455
rect 12817 10421 12851 10455
rect 15209 10421 15243 10455
rect 16313 10421 16347 10455
rect 17417 10421 17451 10455
rect 19533 10421 19567 10455
rect 19809 10421 19843 10455
rect 20177 10421 20211 10455
rect 20269 10421 20303 10455
rect 1685 10217 1719 10251
rect 3249 10217 3283 10251
rect 6929 10217 6963 10251
rect 8217 10217 8251 10251
rect 9229 10217 9263 10251
rect 11437 10217 11471 10251
rect 11897 10217 11931 10251
rect 13829 10217 13863 10251
rect 14841 10217 14875 10251
rect 20453 10217 20487 10251
rect 2421 10149 2455 10183
rect 4322 10149 4356 10183
rect 7021 10149 7055 10183
rect 12909 10149 12943 10183
rect 18613 10149 18647 10183
rect 18981 10149 19015 10183
rect 1501 10081 1535 10115
rect 2513 10081 2547 10115
rect 3065 10081 3099 10115
rect 4077 10081 4111 10115
rect 6101 10081 6135 10115
rect 8125 10081 8159 10115
rect 8953 10081 8987 10115
rect 9045 10081 9079 10115
rect 9689 10081 9723 10115
rect 9945 10081 9979 10115
rect 11805 10081 11839 10115
rect 12817 10081 12851 10115
rect 13921 10081 13955 10115
rect 14657 10081 14691 10115
rect 15568 10081 15602 10115
rect 17693 10081 17727 10115
rect 17785 10081 17819 10115
rect 18347 10081 18381 10115
rect 19340 10081 19374 10115
rect 2605 10013 2639 10047
rect 6193 10013 6227 10047
rect 6285 10013 6319 10047
rect 7113 10013 7147 10047
rect 8401 10013 8435 10047
rect 12081 10013 12115 10047
rect 13093 10013 13127 10047
rect 13369 10013 13403 10047
rect 14013 10013 14047 10047
rect 15301 10013 15335 10047
rect 17141 10013 17175 10047
rect 17877 10013 17911 10047
rect 18981 10013 19015 10047
rect 19073 10013 19107 10047
rect 20913 10013 20947 10047
rect 2053 9877 2087 9911
rect 5457 9877 5491 9911
rect 5733 9877 5767 9911
rect 6561 9877 6595 9911
rect 7573 9877 7607 9911
rect 7757 9877 7791 9911
rect 8769 9877 8803 9911
rect 11069 9877 11103 9911
rect 12449 9877 12483 9911
rect 13369 9877 13403 9911
rect 13461 9877 13495 9911
rect 16681 9877 16715 9911
rect 17325 9877 17359 9911
rect 3157 9673 3191 9707
rect 9229 9673 9263 9707
rect 17601 9673 17635 9707
rect 18061 9673 18095 9707
rect 1777 9605 1811 9639
rect 4169 9605 4203 9639
rect 6377 9605 6411 9639
rect 6837 9605 6871 9639
rect 11345 9605 11379 9639
rect 14381 9605 14415 9639
rect 17141 9605 17175 9639
rect 17325 9605 17359 9639
rect 19073 9605 19107 9639
rect 20085 9605 20119 9639
rect 2697 9537 2731 9571
rect 3709 9537 3743 9571
rect 4721 9537 4755 9571
rect 5733 9537 5767 9571
rect 7389 9537 7423 9571
rect 10149 9537 10183 9571
rect 11069 9537 11103 9571
rect 11897 9537 11931 9571
rect 14933 9537 14967 9571
rect 18613 9537 18647 9571
rect 19717 9537 19751 9571
rect 19993 9537 20027 9571
rect 20637 9537 20671 9571
rect 1593 9469 1627 9503
rect 4629 9469 4663 9503
rect 6193 9469 6227 9503
rect 7849 9469 7883 9503
rect 9873 9469 9907 9503
rect 12449 9469 12483 9503
rect 14281 9469 14315 9503
rect 15761 9469 15795 9503
rect 17325 9469 17359 9503
rect 17417 9469 17451 9503
rect 18429 9469 18463 9503
rect 19441 9469 19475 9503
rect 2605 9401 2639 9435
rect 4537 9401 4571 9435
rect 7297 9401 7331 9435
rect 8116 9401 8150 9435
rect 10977 9401 11011 9435
rect 11713 9401 11747 9435
rect 11805 9401 11839 9435
rect 12716 9401 12750 9435
rect 14749 9401 14783 9435
rect 16028 9401 16062 9435
rect 18521 9401 18555 9435
rect 20453 9469 20487 9503
rect 2145 9333 2179 9367
rect 2513 9333 2547 9367
rect 3525 9333 3559 9367
rect 3617 9333 3651 9367
rect 5181 9333 5215 9367
rect 5549 9333 5583 9367
rect 5641 9333 5675 9367
rect 7205 9333 7239 9367
rect 9505 9333 9539 9367
rect 9965 9333 9999 9367
rect 10517 9333 10551 9367
rect 10885 9333 10919 9367
rect 13829 9333 13863 9367
rect 14105 9333 14139 9367
rect 14841 9333 14875 9367
rect 19533 9333 19567 9367
rect 19993 9333 20027 9367
rect 20545 9333 20579 9367
rect 1961 9129 1995 9163
rect 2421 9129 2455 9163
rect 4077 9129 4111 9163
rect 7021 9129 7055 9163
rect 8769 9129 8803 9163
rect 9229 9129 9263 9163
rect 10057 9129 10091 9163
rect 13001 9129 13035 9163
rect 13553 9129 13587 9163
rect 14841 9129 14875 9163
rect 15301 9129 15335 9163
rect 16313 9129 16347 9163
rect 17233 9129 17267 9163
rect 2329 9061 2363 9095
rect 3341 9061 3375 9095
rect 13093 9061 13127 9095
rect 1409 8993 1443 9027
rect 4445 8993 4479 9027
rect 5089 8993 5123 9027
rect 5356 8993 5390 9027
rect 6837 8993 6871 9027
rect 7389 8993 7423 9027
rect 7656 8993 7690 9027
rect 9045 8993 9079 9027
rect 9413 8993 9447 9027
rect 10149 8993 10183 9027
rect 10609 8993 10643 9027
rect 11244 8993 11278 9027
rect 2605 8925 2639 8959
rect 3433 8925 3467 8959
rect 3525 8925 3559 8959
rect 4537 8925 4571 8959
rect 4629 8925 4663 8959
rect 1593 8857 1627 8891
rect 10241 8925 10275 8959
rect 10977 8925 11011 8959
rect 13185 8925 13219 8959
rect 14013 9061 14047 9095
rect 14657 8993 14691 9027
rect 15669 8993 15703 9027
rect 15761 8993 15795 9027
rect 16681 8993 16715 9027
rect 16773 8993 16807 9027
rect 14105 8925 14139 8959
rect 14289 8925 14323 8959
rect 15025 8925 15059 8959
rect 15853 8925 15887 8959
rect 16865 8925 16899 8959
rect 18153 9129 18187 9163
rect 19717 9129 19751 9163
rect 20913 9129 20947 9163
rect 17693 8993 17727 9027
rect 17785 8993 17819 9027
rect 20269 9061 20303 9095
rect 18337 8993 18371 9027
rect 18604 8993 18638 9027
rect 19993 8993 20027 9027
rect 17969 8925 18003 8959
rect 18153 8925 18187 8959
rect 17233 8857 17267 8891
rect 2973 8789 3007 8823
rect 6469 8789 6503 8823
rect 9413 8789 9447 8823
rect 9689 8789 9723 8823
rect 10793 8789 10827 8823
rect 12357 8789 12391 8823
rect 12633 8789 12667 8823
rect 13553 8789 13587 8823
rect 13645 8789 13679 8823
rect 15025 8789 15059 8823
rect 17325 8789 17359 8823
rect 2421 8585 2455 8619
rect 3617 8585 3651 8619
rect 5365 8585 5399 8619
rect 5733 8585 5767 8619
rect 6561 8585 6595 8619
rect 8401 8585 8435 8619
rect 1869 8449 1903 8483
rect 2053 8449 2087 8483
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 3985 8449 4019 8483
rect 6193 8449 6227 8483
rect 6377 8449 6411 8483
rect 6561 8449 6595 8483
rect 6837 8449 6871 8483
rect 3433 8381 3467 8415
rect 9321 8585 9355 8619
rect 10517 8585 10551 8619
rect 18889 8585 18923 8619
rect 19073 8585 19107 8619
rect 20085 8585 20119 8619
rect 9137 8449 9171 8483
rect 15761 8517 15795 8551
rect 18061 8517 18095 8551
rect 10149 8449 10183 8483
rect 11069 8449 11103 8483
rect 13001 8449 13035 8483
rect 14013 8449 14047 8483
rect 14933 8449 14967 8483
rect 15117 8449 15151 8483
rect 18613 8449 18647 8483
rect 18889 8449 18923 8483
rect 11805 8381 11839 8415
rect 13829 8381 13863 8415
rect 15577 8381 15611 8415
rect 16129 8381 16163 8415
rect 16396 8381 16430 8415
rect 18521 8381 18555 8415
rect 1777 8313 1811 8347
rect 2789 8313 2823 8347
rect 4230 8313 4264 8347
rect 7104 8313 7138 8347
rect 8401 8313 8435 8347
rect 8861 8313 8895 8347
rect 9321 8313 9355 8347
rect 9873 8313 9907 8347
rect 10977 8313 11011 8347
rect 12909 8313 12943 8347
rect 14841 8313 14875 8347
rect 18429 8313 18463 8347
rect 18889 8313 18923 8347
rect 19625 8449 19659 8483
rect 20637 8449 20671 8483
rect 20545 8381 20579 8415
rect 19533 8313 19567 8347
rect 1409 8245 1443 8279
rect 6101 8245 6135 8279
rect 8217 8245 8251 8279
rect 8493 8245 8527 8279
rect 8953 8245 8987 8279
rect 9505 8245 9539 8279
rect 9965 8245 9999 8279
rect 10885 8245 10919 8279
rect 11989 8245 12023 8279
rect 12449 8245 12483 8279
rect 12817 8245 12851 8279
rect 13461 8245 13495 8279
rect 13921 8245 13955 8279
rect 14473 8245 14507 8279
rect 17509 8245 17543 8279
rect 18981 8245 19015 8279
rect 19441 8245 19475 8279
rect 20453 8245 20487 8279
rect 2145 8041 2179 8075
rect 4077 8041 4111 8075
rect 4537 8041 4571 8075
rect 5089 8041 5123 8075
rect 5549 8041 5583 8075
rect 6929 8041 6963 8075
rect 7389 8041 7423 8075
rect 14933 8041 14967 8075
rect 15025 8041 15059 8075
rect 15301 8041 15335 8075
rect 18613 8041 18647 8075
rect 19809 8041 19843 8075
rect 21833 8041 21867 8075
rect 10876 7973 10910 8007
rect 12633 7973 12667 8007
rect 12725 7973 12759 8007
rect 1593 7905 1627 7939
rect 1869 7905 1903 7939
rect 2145 7905 2179 7939
rect 2596 7905 2630 7939
rect 4445 7905 4479 7939
rect 5457 7905 5491 7939
rect 6285 7905 6319 7939
rect 6377 7905 6411 7939
rect 7297 7905 7331 7939
rect 7941 7905 7975 7939
rect 8208 7905 8242 7939
rect 9965 7905 9999 7939
rect 10609 7905 10643 7939
rect 13461 7905 13495 7939
rect 13820 7905 13854 7939
rect 2329 7837 2363 7871
rect 4629 7837 4663 7871
rect 5641 7837 5675 7871
rect 7573 7837 7607 7871
rect 12909 7837 12943 7871
rect 13185 7837 13219 7871
rect 13553 7837 13587 7871
rect 3709 7769 3743 7803
rect 6101 7769 6135 7803
rect 9321 7769 9355 7803
rect 15669 7905 15703 7939
rect 16497 7905 16531 7939
rect 16589 7905 16623 7939
rect 17141 7905 17175 7939
rect 17397 7905 17431 7939
rect 18981 7905 19015 7939
rect 19073 7905 19107 7939
rect 20177 7905 20211 7939
rect 15761 7837 15795 7871
rect 15853 7837 15887 7871
rect 19257 7837 19291 7871
rect 20269 7837 20303 7871
rect 20361 7837 20395 7871
rect 15025 7769 15059 7803
rect 19717 7769 19751 7803
rect 6561 7701 6595 7735
rect 10149 7701 10183 7735
rect 11989 7701 12023 7735
rect 12265 7701 12299 7735
rect 13185 7701 13219 7735
rect 13277 7701 13311 7735
rect 16313 7701 16347 7735
rect 16773 7701 16807 7735
rect 18521 7701 18555 7735
rect 3157 7497 3191 7531
rect 5181 7497 5215 7531
rect 5457 7497 5491 7531
rect 8861 7497 8895 7531
rect 16405 7497 16439 7531
rect 17601 7497 17635 7531
rect 18889 7497 18923 7531
rect 20085 7497 20119 7531
rect 8493 7429 8527 7463
rect 14105 7429 14139 7463
rect 6009 7361 6043 7395
rect 9413 7361 9447 7395
rect 10517 7361 10551 7395
rect 11437 7361 11471 7395
rect 14657 7361 14691 7395
rect 15853 7361 15887 7395
rect 16037 7361 16071 7395
rect 16957 7361 16991 7395
rect 18613 7361 18647 7395
rect 1777 7293 1811 7327
rect 2044 7293 2078 7327
rect 3801 7293 3835 7327
rect 5825 7293 5859 7327
rect 7113 7293 7147 7327
rect 9321 7293 9355 7327
rect 12449 7293 12483 7327
rect 12716 7293 12750 7327
rect 14013 7293 14047 7327
rect 14473 7293 14507 7327
rect 17417 7293 17451 7327
rect 18429 7293 18463 7327
rect 4046 7225 4080 7259
rect 7380 7225 7414 7259
rect 10333 7225 10367 7259
rect 11253 7225 11287 7259
rect 11897 7225 11931 7259
rect 14565 7225 14599 7259
rect 16865 7225 16899 7259
rect 19717 7361 19751 7395
rect 20637 7361 20671 7395
rect 5917 7157 5951 7191
rect 9229 7157 9263 7191
rect 9873 7157 9907 7191
rect 10241 7157 10275 7191
rect 10885 7157 10919 7191
rect 11345 7157 11379 7191
rect 13829 7157 13863 7191
rect 14013 7157 14047 7191
rect 15393 7157 15427 7191
rect 15761 7157 15795 7191
rect 16773 7157 16807 7191
rect 18061 7157 18095 7191
rect 18521 7157 18555 7191
rect 18889 7157 18923 7191
rect 18981 7293 19015 7327
rect 19533 7293 19567 7327
rect 18981 7157 19015 7191
rect 19073 7157 19107 7191
rect 19441 7157 19475 7191
rect 20453 7157 20487 7191
rect 20545 7157 20579 7191
rect 2513 6953 2547 6987
rect 3617 6953 3651 6987
rect 8953 6953 8987 6987
rect 10241 6953 10275 6987
rect 10333 6953 10367 6987
rect 11253 6953 11287 6987
rect 11345 6953 11379 6987
rect 11897 6953 11931 6987
rect 13277 6953 13311 6987
rect 13921 6953 13955 6987
rect 15669 6953 15703 6987
rect 16497 6953 16531 6987
rect 17233 6953 17267 6987
rect 17877 6953 17911 6987
rect 18337 6953 18371 6987
rect 2605 6885 2639 6919
rect 4445 6885 4479 6919
rect 5641 6885 5675 6919
rect 7665 6885 7699 6919
rect 8217 6885 8251 6919
rect 12265 6885 12299 6919
rect 18245 6885 18279 6919
rect 1593 6817 1627 6851
rect 3433 6817 3467 6851
rect 6469 6817 6503 6851
rect 2697 6749 2731 6783
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 5733 6749 5767 6783
rect 5825 6749 5859 6783
rect 6561 6749 6595 6783
rect 6745 6749 6779 6783
rect 7757 6749 7791 6783
rect 7941 6749 7975 6783
rect 8493 6817 8527 6851
rect 9045 6817 9079 6851
rect 14289 6817 14323 6851
rect 16313 6817 16347 6851
rect 19432 6817 19466 6851
rect 9229 6749 9263 6783
rect 10425 6749 10459 6783
rect 10793 6749 10827 6783
rect 11529 6749 11563 6783
rect 12357 6749 12391 6783
rect 12541 6749 12575 6783
rect 13369 6749 13403 6783
rect 13461 6749 13495 6783
rect 14381 6749 14415 6783
rect 14473 6749 14507 6783
rect 15761 6749 15795 6783
rect 15945 6749 15979 6783
rect 17325 6749 17359 6783
rect 17509 6749 17543 6783
rect 18521 6749 18555 6783
rect 19073 6749 19107 6783
rect 19165 6749 19199 6783
rect 20913 6749 20947 6783
rect 1777 6681 1811 6715
rect 4077 6681 4111 6715
rect 7297 6681 7331 6715
rect 8217 6681 8251 6715
rect 9873 6681 9907 6715
rect 12909 6681 12943 6715
rect 15301 6681 15335 6715
rect 20545 6681 20579 6715
rect 2145 6613 2179 6647
rect 5273 6613 5307 6647
rect 6101 6613 6135 6647
rect 7113 6613 7147 6647
rect 8309 6613 8343 6647
rect 8585 6613 8619 6647
rect 10793 6613 10827 6647
rect 10885 6613 10919 6647
rect 16865 6613 16899 6647
rect 19073 6613 19107 6647
rect 1593 6409 1627 6443
rect 3617 6409 3651 6443
rect 8769 6409 8803 6443
rect 14657 6409 14691 6443
rect 16865 6409 16899 6443
rect 16957 6409 16991 6443
rect 19257 6409 19291 6443
rect 20729 6409 20763 6443
rect 3341 6341 3375 6375
rect 4905 6341 4939 6375
rect 5181 6341 5215 6375
rect 5273 6341 5307 6375
rect 7481 6341 7515 6375
rect 7573 6341 7607 6375
rect 14013 6341 14047 6375
rect 16405 6341 16439 6375
rect 4169 6273 4203 6307
rect 1409 6205 1443 6239
rect 1961 6205 1995 6239
rect 4721 6205 4755 6239
rect 5825 6273 5859 6307
rect 6285 6273 6319 6307
rect 8401 6273 8435 6307
rect 9413 6273 9447 6307
rect 9597 6273 9631 6307
rect 15025 6273 15059 6307
rect 5641 6205 5675 6239
rect 5733 6205 5767 6239
rect 7021 6205 7055 6239
rect 7481 6205 7515 6239
rect 8217 6205 8251 6239
rect 9229 6205 9263 6239
rect 2228 6137 2262 6171
rect 4077 6137 4111 6171
rect 5181 6137 5215 6171
rect 8125 6137 8159 6171
rect 9781 6205 9815 6239
rect 11805 6205 11839 6239
rect 12633 6205 12667 6239
rect 14473 6205 14507 6239
rect 17417 6273 17451 6307
rect 17601 6273 17635 6307
rect 18521 6273 18555 6307
rect 18613 6273 18647 6307
rect 19349 6273 19383 6307
rect 19257 6205 19291 6239
rect 10048 6137 10082 6171
rect 12900 6137 12934 6171
rect 15292 6137 15326 6171
rect 16865 6137 16899 6171
rect 18429 6137 18463 6171
rect 19616 6137 19650 6171
rect 3985 6069 4019 6103
rect 7205 6069 7239 6103
rect 7757 6069 7791 6103
rect 9137 6069 9171 6103
rect 9597 6069 9631 6103
rect 11161 6069 11195 6103
rect 11989 6069 12023 6103
rect 17325 6069 17359 6103
rect 18061 6069 18095 6103
rect 1777 5865 1811 5899
rect 5457 5865 5491 5899
rect 7021 5865 7055 5899
rect 7205 5865 7239 5899
rect 8217 5865 8251 5899
rect 14473 5865 14507 5899
rect 14749 5865 14783 5899
rect 15853 5865 15887 5899
rect 18521 5865 18555 5899
rect 19349 5865 19383 5899
rect 20361 5865 20395 5899
rect 2504 5797 2538 5831
rect 5733 5797 5767 5831
rect 4344 5729 4378 5763
rect 6561 5729 6595 5763
rect 6653 5729 6687 5763
rect 2237 5661 2271 5695
rect 4077 5661 4111 5695
rect 6837 5661 6871 5695
rect 7573 5797 7607 5831
rect 8125 5797 8159 5831
rect 8585 5797 8619 5831
rect 8677 5797 8711 5831
rect 9956 5797 9990 5831
rect 11805 5797 11839 5831
rect 13360 5797 13394 5831
rect 18613 5797 18647 5831
rect 7665 5661 7699 5695
rect 7849 5661 7883 5695
rect 9689 5729 9723 5763
rect 11713 5729 11747 5763
rect 12541 5729 12575 5763
rect 16681 5729 16715 5763
rect 16948 5729 16982 5763
rect 19165 5729 19199 5763
rect 19717 5729 19751 5763
rect 19809 5729 19843 5763
rect 8769 5661 8803 5695
rect 11989 5661 12023 5695
rect 13093 5661 13127 5695
rect 15945 5661 15979 5695
rect 16037 5661 16071 5695
rect 18705 5661 18739 5695
rect 19993 5661 20027 5695
rect 8125 5593 8159 5627
rect 15485 5593 15519 5627
rect 18153 5593 18187 5627
rect 3617 5525 3651 5559
rect 6193 5525 6227 5559
rect 7021 5525 7055 5559
rect 11069 5525 11103 5559
rect 11345 5525 11379 5559
rect 12725 5525 12759 5559
rect 18061 5525 18095 5559
rect 3341 5321 3375 5355
rect 5733 5321 5767 5355
rect 8217 5321 8251 5355
rect 10333 5321 10367 5355
rect 14749 5321 14783 5355
rect 17141 5321 17175 5355
rect 20177 5321 20211 5355
rect 6653 5253 6687 5287
rect 1593 5185 1627 5219
rect 2697 5185 2731 5219
rect 3985 5185 4019 5219
rect 4997 5185 5031 5219
rect 6377 5185 6411 5219
rect 1409 5117 1443 5151
rect 4813 5117 4847 5151
rect 6101 5117 6135 5151
rect 10609 5253 10643 5287
rect 13369 5253 13403 5287
rect 13461 5253 13495 5287
rect 17601 5253 17635 5287
rect 11437 5185 11471 5219
rect 11529 5185 11563 5219
rect 13093 5185 13127 5219
rect 6837 5117 6871 5151
rect 8769 5117 8803 5151
rect 9036 5117 9070 5151
rect 10333 5117 10367 5151
rect 10425 5117 10459 5151
rect 12909 5117 12943 5151
rect 3709 5049 3743 5083
rect 6653 5049 6687 5083
rect 7082 5049 7116 5083
rect 11345 5049 11379 5083
rect 14197 5185 14231 5219
rect 15209 5185 15243 5219
rect 15393 5185 15427 5219
rect 15761 5185 15795 5219
rect 18797 5185 18831 5219
rect 20637 5185 20671 5219
rect 14013 5117 14047 5151
rect 16028 5117 16062 5151
rect 17417 5117 17451 5151
rect 18061 5117 18095 5151
rect 20453 5117 20487 5151
rect 14105 5049 14139 5083
rect 15117 5049 15151 5083
rect 18337 5049 18371 5083
rect 19064 5049 19098 5083
rect 2145 4981 2179 5015
rect 2513 4981 2547 5015
rect 2605 4981 2639 5015
rect 3801 4981 3835 5015
rect 4353 4981 4387 5015
rect 4721 4981 4755 5015
rect 6193 4981 6227 5015
rect 10149 4981 10183 5015
rect 10977 4981 11011 5015
rect 12449 4981 12483 5015
rect 12817 4981 12851 5015
rect 13461 4981 13495 5015
rect 13645 4981 13679 5015
rect 2881 4777 2915 4811
rect 3617 4777 3651 4811
rect 4077 4777 4111 4811
rect 4537 4777 4571 4811
rect 7021 4777 7055 4811
rect 7297 4777 7331 4811
rect 7665 4777 7699 4811
rect 7757 4777 7791 4811
rect 8309 4777 8343 4811
rect 8677 4777 8711 4811
rect 10241 4777 10275 4811
rect 10425 4777 10459 4811
rect 10885 4777 10919 4811
rect 11805 4777 11839 4811
rect 12909 4777 12943 4811
rect 13829 4777 13863 4811
rect 15301 4777 15335 4811
rect 16129 4777 16163 4811
rect 1768 4641 1802 4675
rect 3433 4641 3467 4675
rect 4445 4641 4479 4675
rect 5089 4641 5123 4675
rect 5897 4641 5931 4675
rect 8769 4641 8803 4675
rect 9873 4641 9907 4675
rect 1501 4573 1535 4607
rect 4629 4573 4663 4607
rect 5641 4573 5675 4607
rect 7849 4573 7883 4607
rect 8861 4573 8895 4607
rect 12265 4709 12299 4743
rect 10793 4641 10827 4675
rect 11069 4573 11103 4607
rect 11897 4573 11931 4607
rect 11989 4573 12023 4607
rect 17408 4709 17442 4743
rect 12817 4641 12851 4675
rect 13921 4641 13955 4675
rect 14657 4641 14691 4675
rect 15669 4641 15703 4675
rect 16129 4641 16163 4675
rect 16313 4641 16347 4675
rect 17141 4641 17175 4675
rect 19441 4641 19475 4675
rect 20085 4641 20119 4675
rect 13001 4573 13035 4607
rect 14013 4573 14047 4607
rect 15761 4573 15795 4607
rect 15945 4573 15979 4607
rect 16589 4573 16623 4607
rect 19533 4573 19567 4607
rect 19717 4573 19751 4607
rect 20361 4573 20395 4607
rect 20913 4573 20947 4607
rect 13461 4505 13495 4539
rect 5273 4437 5307 4471
rect 10057 4437 10091 4471
rect 10241 4437 10275 4471
rect 11437 4437 11471 4471
rect 12265 4437 12299 4471
rect 12449 4437 12483 4471
rect 14841 4437 14875 4471
rect 18521 4437 18555 4471
rect 19073 4437 19107 4471
rect 3709 4233 3743 4267
rect 2513 4097 2547 4131
rect 3433 4097 3467 4131
rect 6101 4233 6135 4267
rect 14473 4233 14507 4267
rect 14749 4233 14783 4267
rect 19717 4233 19751 4267
rect 4537 4097 4571 4131
rect 5457 4097 5491 4131
rect 16773 4165 16807 4199
rect 7297 4097 7331 4131
rect 7481 4097 7515 4131
rect 8585 4097 8619 4131
rect 11621 4097 11655 4131
rect 11713 4097 11747 4131
rect 13093 4097 13127 4131
rect 15209 4097 15243 4131
rect 15301 4097 15335 4131
rect 16405 4097 16439 4131
rect 17417 4097 17451 4131
rect 18061 4097 18095 4131
rect 20269 4097 20303 4131
rect 1409 4029 1443 4063
rect 3709 4029 3743 4063
rect 4261 4029 4295 4063
rect 5273 4029 5307 4063
rect 5365 4029 5399 4063
rect 6101 4029 6135 4063
rect 6193 4029 6227 4063
rect 7205 4029 7239 4063
rect 8033 4029 8067 4063
rect 10241 4029 10275 4063
rect 10517 4029 10551 4063
rect 12541 4029 12575 4063
rect 16129 4029 16163 4063
rect 20085 4029 20119 4063
rect 20729 4029 20763 4063
rect 2237 3961 2271 3995
rect 3249 3961 3283 3995
rect 8852 3961 8886 3995
rect 11529 3961 11563 3995
rect 13360 3961 13394 3995
rect 17233 3961 17267 3995
rect 18328 3961 18362 3995
rect 20177 3961 20211 3995
rect 1869 3893 1903 3927
rect 2329 3893 2363 3927
rect 2881 3893 2915 3927
rect 3341 3893 3375 3927
rect 3893 3893 3927 3927
rect 4353 3893 4387 3927
rect 4905 3893 4939 3927
rect 6377 3893 6411 3927
rect 6837 3893 6871 3927
rect 8217 3893 8251 3927
rect 9965 3893 9999 3927
rect 11161 3893 11195 3927
rect 12725 3893 12759 3927
rect 15117 3893 15151 3927
rect 15761 3893 15795 3927
rect 16221 3893 16255 3927
rect 17141 3893 17175 3927
rect 19441 3893 19475 3927
rect 20913 3893 20947 3927
rect 4169 3689 4203 3723
rect 4261 3689 4295 3723
rect 4813 3689 4847 3723
rect 5825 3689 5859 3723
rect 9689 3689 9723 3723
rect 10057 3689 10091 3723
rect 12265 3689 12299 3723
rect 12449 3689 12483 3723
rect 12817 3689 12851 3723
rect 13461 3689 13495 3723
rect 13921 3689 13955 3723
rect 18429 3689 18463 3723
rect 18521 3689 18555 3723
rect 19165 3689 19199 3723
rect 19533 3689 19567 3723
rect 2228 3553 2262 3587
rect 1501 3485 1535 3519
rect 1961 3485 1995 3519
rect 3341 3417 3375 3451
rect 5917 3621 5951 3655
rect 8125 3621 8159 3655
rect 5365 3553 5399 3587
rect 7021 3553 7055 3587
rect 8033 3553 8067 3587
rect 8861 3553 8895 3587
rect 9137 3553 9171 3587
rect 11060 3553 11094 3587
rect 4905 3485 4939 3519
rect 5089 3485 5123 3519
rect 6009 3485 6043 3519
rect 7113 3485 7147 3519
rect 7297 3485 7331 3519
rect 8309 3485 8343 3519
rect 10149 3485 10183 3519
rect 10241 3485 10275 3519
rect 10793 3485 10827 3519
rect 5457 3417 5491 3451
rect 12909 3621 12943 3655
rect 19625 3621 19659 3655
rect 13829 3553 13863 3587
rect 14473 3553 14507 3587
rect 14749 3553 14783 3587
rect 15301 3553 15335 3587
rect 15853 3553 15887 3587
rect 16120 3553 16154 3587
rect 17509 3553 17543 3587
rect 20177 3553 20211 3587
rect 13001 3485 13035 3519
rect 14105 3485 14139 3519
rect 18705 3485 18739 3519
rect 19809 3485 19843 3519
rect 20913 3485 20947 3519
rect 4169 3349 4203 3383
rect 4445 3349 4479 3383
rect 6653 3349 6687 3383
rect 7665 3349 7699 3383
rect 12173 3349 12207 3383
rect 12265 3349 12299 3383
rect 15485 3349 15519 3383
rect 17233 3349 17267 3383
rect 17693 3349 17727 3383
rect 18061 3349 18095 3383
rect 20361 3349 20395 3383
rect 1685 3145 1719 3179
rect 2697 3145 2731 3179
rect 5273 3145 5307 3179
rect 5733 3145 5767 3179
rect 8217 3145 8251 3179
rect 9873 3145 9907 3179
rect 13737 3145 13771 3179
rect 14657 3145 14691 3179
rect 14841 3145 14875 3179
rect 16405 3145 16439 3179
rect 18245 3145 18279 3179
rect 19441 3145 19475 3179
rect 12081 3077 12115 3111
rect 12541 3077 12575 3111
rect 13829 3077 13863 3111
rect 15669 3077 15703 3111
rect 16037 3077 16071 3111
rect 2329 3009 2363 3043
rect 3341 3009 3375 3043
rect 6285 3009 6319 3043
rect 2053 2941 2087 2975
rect 3893 2941 3927 2975
rect 6837 2941 6871 2975
rect 8493 2941 8527 2975
rect 8760 2941 8794 2975
rect 10149 2941 10183 2975
rect 10701 2941 10735 2975
rect 10968 2941 11002 2975
rect 4160 2873 4194 2907
rect 6101 2873 6135 2907
rect 7104 2873 7138 2907
rect 13093 3009 13127 3043
rect 13277 3009 13311 3043
rect 14289 3009 14323 3043
rect 14473 3009 14507 3043
rect 15301 3009 15335 3043
rect 15485 3009 15519 3043
rect 17049 3009 17083 3043
rect 18889 3009 18923 3043
rect 19993 3009 20027 3043
rect 13001 2941 13035 2975
rect 14197 2941 14231 2975
rect 15209 2941 15243 2975
rect 15853 2941 15887 2975
rect 16773 2941 16807 2975
rect 16865 2941 16899 2975
rect 17417 2941 17451 2975
rect 19901 2941 19935 2975
rect 20453 2941 20487 2975
rect 18613 2873 18647 2907
rect 19809 2873 19843 2907
rect 20729 2873 20763 2907
rect 2145 2805 2179 2839
rect 3065 2805 3099 2839
rect 3157 2805 3191 2839
rect 6193 2805 6227 2839
rect 10333 2805 10367 2839
rect 12541 2805 12575 2839
rect 12633 2805 12667 2839
rect 17601 2805 17635 2839
rect 18705 2805 18739 2839
rect 1961 2601 1995 2635
rect 2329 2601 2363 2635
rect 2973 2601 3007 2635
rect 3341 2601 3375 2635
rect 5457 2601 5491 2635
rect 5825 2601 5859 2635
rect 6929 2601 6963 2635
rect 7297 2601 7331 2635
rect 10149 2601 10183 2635
rect 11253 2601 11287 2635
rect 14381 2601 14415 2635
rect 16221 2601 16255 2635
rect 16681 2601 16715 2635
rect 18337 2601 18371 2635
rect 18797 2601 18831 2635
rect 19349 2601 19383 2635
rect 19717 2601 19751 2635
rect 2421 2533 2455 2567
rect 4322 2533 4356 2567
rect 6193 2533 6227 2567
rect 8309 2533 8343 2567
rect 11161 2533 11195 2567
rect 12081 2533 12115 2567
rect 12909 2533 12943 2567
rect 15761 2533 15795 2567
rect 17601 2533 17635 2567
rect 19809 2533 19843 2567
rect 20637 2533 20671 2567
rect 4077 2465 4111 2499
rect 7389 2465 7423 2499
rect 8401 2465 8435 2499
rect 9137 2465 9171 2499
rect 11805 2465 11839 2499
rect 12633 2465 12667 2499
rect 13737 2465 13771 2499
rect 14749 2465 14783 2499
rect 14841 2465 14875 2499
rect 15485 2465 15519 2499
rect 16589 2465 16623 2499
rect 18705 2465 18739 2499
rect 20361 2465 20395 2499
rect 2605 2397 2639 2431
rect 3433 2397 3467 2431
rect 3617 2397 3651 2431
rect 6285 2397 6319 2431
rect 6377 2397 6411 2431
rect 7573 2397 7607 2431
rect 8585 2397 8619 2431
rect 10241 2397 10275 2431
rect 10333 2397 10367 2431
rect 11437 2397 11471 2431
rect 13829 2397 13863 2431
rect 14013 2397 14047 2431
rect 15025 2397 15059 2431
rect 15209 2397 15243 2431
rect 16773 2397 16807 2431
rect 17693 2397 17727 2431
rect 17877 2397 17911 2431
rect 18981 2397 19015 2431
rect 19901 2397 19935 2431
rect 7941 2329 7975 2363
rect 9781 2329 9815 2363
rect 13369 2329 13403 2363
rect 9321 2261 9355 2295
rect 10793 2261 10827 2295
rect 15209 2261 15243 2295
rect 17233 2261 17267 2295
<< metal1 >>
rect 3878 21224 3884 21276
rect 3936 21264 3942 21276
rect 8294 21264 8300 21276
rect 3936 21236 8300 21264
rect 3936 21224 3942 21236
rect 8294 21224 8300 21236
rect 8352 21224 8358 21276
rect 4062 20952 4068 21004
rect 4120 20992 4126 21004
rect 5994 20992 6000 21004
rect 4120 20964 6000 20992
rect 4120 20952 4126 20964
rect 5994 20952 6000 20964
rect 6052 20952 6058 21004
rect 3786 20612 3792 20664
rect 3844 20652 3850 20664
rect 11606 20652 11612 20664
rect 3844 20624 11612 20652
rect 3844 20612 3850 20624
rect 11606 20612 11612 20624
rect 11664 20612 11670 20664
rect 15286 20612 15292 20664
rect 15344 20652 15350 20664
rect 19518 20652 19524 20664
rect 15344 20624 19524 20652
rect 15344 20612 15350 20624
rect 19518 20612 19524 20624
rect 19576 20612 19582 20664
rect 8754 20544 8760 20596
rect 8812 20584 8818 20596
rect 19334 20584 19340 20596
rect 8812 20556 19340 20584
rect 8812 20544 8818 20556
rect 19334 20544 19340 20556
rect 19392 20544 19398 20596
rect 4982 20408 4988 20460
rect 5040 20448 5046 20460
rect 12250 20448 12256 20460
rect 5040 20420 12256 20448
rect 5040 20408 5046 20420
rect 12250 20408 12256 20420
rect 12308 20408 12314 20460
rect 566 20272 572 20324
rect 624 20312 630 20324
rect 5350 20312 5356 20324
rect 624 20284 5356 20312
rect 624 20272 630 20284
rect 5350 20272 5356 20284
rect 5408 20272 5414 20324
rect 7558 20272 7564 20324
rect 7616 20312 7622 20324
rect 15102 20312 15108 20324
rect 7616 20284 15108 20312
rect 7616 20272 7622 20284
rect 15102 20272 15108 20284
rect 15160 20272 15166 20324
rect 5368 20244 5396 20272
rect 8478 20244 8484 20256
rect 5368 20216 8484 20244
rect 8478 20204 8484 20216
rect 8536 20204 8542 20256
rect 8662 20204 8668 20256
rect 8720 20244 8726 20256
rect 9306 20244 9312 20256
rect 8720 20216 9312 20244
rect 8720 20204 8726 20216
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 13998 20204 14004 20256
rect 14056 20244 14062 20256
rect 15010 20244 15016 20256
rect 14056 20216 15016 20244
rect 14056 20204 14062 20216
rect 15010 20204 15016 20216
rect 15068 20204 15074 20256
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 7558 20040 7564 20052
rect 2424 20012 7564 20040
rect 1946 19972 1952 19984
rect 1907 19944 1952 19972
rect 1946 19932 1952 19944
rect 2004 19932 2010 19984
rect 1673 19907 1731 19913
rect 1673 19873 1685 19907
rect 1719 19904 1731 19907
rect 2314 19904 2320 19916
rect 1719 19876 2320 19904
rect 1719 19873 1731 19876
rect 1673 19867 1731 19873
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 2424 19913 2452 20012
rect 7558 20000 7564 20012
rect 7616 20000 7622 20052
rect 7650 20000 7656 20052
rect 7708 20040 7714 20052
rect 8941 20043 8999 20049
rect 8941 20040 8953 20043
rect 7708 20012 8953 20040
rect 7708 20000 7714 20012
rect 8941 20009 8953 20012
rect 8987 20009 8999 20043
rect 8941 20003 8999 20009
rect 11149 20043 11207 20049
rect 11149 20009 11161 20043
rect 11195 20040 11207 20043
rect 12710 20040 12716 20052
rect 11195 20012 12716 20040
rect 11195 20009 11207 20012
rect 11149 20003 11207 20009
rect 12710 20000 12716 20012
rect 12768 20000 12774 20052
rect 13541 20043 13599 20049
rect 13541 20009 13553 20043
rect 13587 20040 13599 20043
rect 13814 20040 13820 20052
rect 13587 20012 13820 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 13814 20000 13820 20012
rect 13872 20000 13878 20052
rect 16393 20043 16451 20049
rect 16393 20009 16405 20043
rect 16439 20040 16451 20043
rect 19058 20040 19064 20052
rect 16439 20012 19064 20040
rect 16439 20009 16451 20012
rect 16393 20003 16451 20009
rect 19058 20000 19064 20012
rect 19116 20000 19122 20052
rect 21818 20040 21824 20052
rect 19352 20012 21824 20040
rect 6365 19975 6423 19981
rect 6365 19972 6377 19975
rect 3436 19944 6377 19972
rect 3436 19913 3464 19944
rect 6365 19941 6377 19944
rect 6411 19941 6423 19975
rect 8018 19972 8024 19984
rect 6365 19935 6423 19941
rect 6932 19944 8024 19972
rect 2409 19907 2467 19913
rect 2409 19873 2421 19907
rect 2455 19873 2467 19907
rect 2409 19867 2467 19873
rect 3421 19907 3479 19913
rect 3421 19873 3433 19907
rect 3467 19873 3479 19907
rect 3421 19867 3479 19873
rect 3510 19864 3516 19916
rect 3568 19904 3574 19916
rect 4433 19907 4491 19913
rect 4433 19904 4445 19907
rect 3568 19876 4445 19904
rect 3568 19864 3574 19876
rect 4433 19873 4445 19876
rect 4479 19873 4491 19907
rect 4890 19904 4896 19916
rect 4433 19867 4491 19873
rect 4540 19876 4896 19904
rect 2685 19839 2743 19845
rect 2685 19805 2697 19839
rect 2731 19836 2743 19839
rect 2774 19836 2780 19848
rect 2731 19808 2780 19836
rect 2731 19805 2743 19808
rect 2685 19799 2743 19805
rect 2774 19796 2780 19808
rect 2832 19796 2838 19848
rect 4540 19845 4568 19876
rect 4890 19864 4896 19876
rect 4948 19864 4954 19916
rect 5350 19864 5356 19916
rect 5408 19904 5414 19916
rect 5445 19907 5503 19913
rect 5445 19904 5457 19907
rect 5408 19876 5457 19904
rect 5408 19864 5414 19876
rect 5445 19873 5457 19876
rect 5491 19873 5503 19907
rect 6086 19904 6092 19916
rect 6047 19876 6092 19904
rect 5445 19867 5503 19873
rect 6086 19864 6092 19876
rect 6144 19864 6150 19916
rect 4525 19839 4583 19845
rect 4525 19836 4537 19839
rect 3528 19808 4537 19836
rect 1670 19728 1676 19780
rect 1728 19768 1734 19780
rect 3528 19768 3556 19808
rect 4525 19805 4537 19808
rect 4571 19805 4583 19839
rect 4525 19799 4583 19805
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19805 4767 19839
rect 4709 19799 4767 19805
rect 1728 19740 3556 19768
rect 3605 19771 3663 19777
rect 1728 19728 1734 19740
rect 3605 19737 3617 19771
rect 3651 19768 3663 19771
rect 3786 19768 3792 19780
rect 3651 19740 3792 19768
rect 3651 19737 3663 19740
rect 3605 19731 3663 19737
rect 3786 19728 3792 19740
rect 3844 19728 3850 19780
rect 4724 19768 4752 19799
rect 5258 19796 5264 19848
rect 5316 19836 5322 19848
rect 5537 19839 5595 19845
rect 5537 19836 5549 19839
rect 5316 19808 5549 19836
rect 5316 19796 5322 19808
rect 5537 19805 5549 19808
rect 5583 19805 5595 19839
rect 5537 19799 5595 19805
rect 5721 19839 5779 19845
rect 5721 19805 5733 19839
rect 5767 19836 5779 19839
rect 5767 19808 6408 19836
rect 5767 19805 5779 19808
rect 5721 19799 5779 19805
rect 5166 19768 5172 19780
rect 4724 19740 5172 19768
rect 5166 19728 5172 19740
rect 5224 19728 5230 19780
rect 5350 19728 5356 19780
rect 5408 19768 5414 19780
rect 5736 19768 5764 19799
rect 5408 19740 5764 19768
rect 5408 19728 5414 19740
rect 4062 19700 4068 19712
rect 4023 19672 4068 19700
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 5077 19703 5135 19709
rect 5077 19669 5089 19703
rect 5123 19700 5135 19703
rect 6178 19700 6184 19712
rect 5123 19672 6184 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 6178 19660 6184 19672
rect 6236 19660 6242 19712
rect 6380 19700 6408 19808
rect 6638 19796 6644 19848
rect 6696 19836 6702 19848
rect 6932 19845 6960 19944
rect 8018 19932 8024 19944
rect 8076 19932 8082 19984
rect 8404 19944 9168 19972
rect 8404 19916 8432 19944
rect 7184 19907 7242 19913
rect 7184 19873 7196 19907
rect 7230 19904 7242 19907
rect 8386 19904 8392 19916
rect 7230 19876 8392 19904
rect 7230 19873 7242 19876
rect 7184 19867 7242 19873
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 6917 19839 6975 19845
rect 6917 19836 6929 19839
rect 6696 19808 6929 19836
rect 6696 19796 6702 19808
rect 6917 19805 6929 19808
rect 6963 19805 6975 19839
rect 9030 19836 9036 19848
rect 8991 19808 9036 19836
rect 6917 19799 6975 19805
rect 9030 19796 9036 19808
rect 9088 19796 9094 19848
rect 9140 19845 9168 19944
rect 9858 19932 9864 19984
rect 9916 19972 9922 19984
rect 11977 19975 12035 19981
rect 9916 19944 11008 19972
rect 9916 19932 9922 19944
rect 9490 19864 9496 19916
rect 9548 19904 9554 19916
rect 10980 19913 11008 19944
rect 11977 19941 11989 19975
rect 12023 19972 12035 19975
rect 12158 19972 12164 19984
rect 12023 19944 12164 19972
rect 12023 19941 12035 19944
rect 11977 19935 12035 19941
rect 12158 19932 12164 19944
rect 12216 19932 12222 19984
rect 12250 19932 12256 19984
rect 12308 19972 12314 19984
rect 14737 19975 14795 19981
rect 14737 19972 14749 19975
rect 12308 19944 14749 19972
rect 12308 19932 12314 19944
rect 14737 19941 14749 19944
rect 14783 19941 14795 19975
rect 15470 19972 15476 19984
rect 14737 19935 14795 19941
rect 15120 19944 15476 19972
rect 15120 19916 15148 19944
rect 15470 19932 15476 19944
rect 15528 19972 15534 19984
rect 16574 19972 16580 19984
rect 15528 19944 16580 19972
rect 15528 19932 15534 19944
rect 16574 19932 16580 19944
rect 16632 19972 16638 19984
rect 17037 19975 17095 19981
rect 16632 19944 16804 19972
rect 16632 19932 16638 19944
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 9548 19876 10149 19904
rect 9548 19864 9554 19876
rect 10137 19873 10149 19876
rect 10183 19873 10195 19907
rect 10137 19867 10195 19873
rect 10965 19907 11023 19913
rect 10965 19873 10977 19907
rect 11011 19873 11023 19907
rect 10965 19867 11023 19873
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19904 11943 19907
rect 12434 19904 12440 19916
rect 11931 19876 12440 19904
rect 11931 19873 11943 19876
rect 11885 19867 11943 19873
rect 12434 19864 12440 19876
rect 12492 19864 12498 19916
rect 12618 19904 12624 19916
rect 12579 19876 12624 19904
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 12897 19907 12955 19913
rect 12897 19873 12909 19907
rect 12943 19904 12955 19907
rect 13357 19907 13415 19913
rect 13357 19904 13369 19907
rect 12943 19876 13369 19904
rect 12943 19873 12955 19876
rect 12897 19867 12955 19873
rect 13357 19873 13369 19876
rect 13403 19873 13415 19907
rect 13906 19904 13912 19916
rect 13867 19876 13912 19904
rect 13357 19867 13415 19873
rect 13906 19864 13912 19876
rect 13964 19864 13970 19916
rect 14458 19904 14464 19916
rect 14419 19876 14464 19904
rect 14458 19864 14464 19876
rect 14516 19864 14522 19916
rect 15013 19907 15071 19913
rect 15013 19873 15025 19907
rect 15059 19904 15071 19907
rect 15102 19904 15108 19916
rect 15059 19876 15108 19904
rect 15059 19873 15071 19876
rect 15013 19867 15071 19873
rect 15102 19864 15108 19876
rect 15160 19864 15166 19916
rect 15654 19904 15660 19916
rect 15615 19876 15660 19904
rect 15654 19864 15660 19876
rect 15712 19864 15718 19916
rect 16776 19913 16804 19944
rect 17037 19941 17049 19975
rect 17083 19972 17095 19975
rect 19150 19972 19156 19984
rect 17083 19944 19012 19972
rect 19111 19944 19156 19972
rect 17083 19941 17095 19944
rect 17037 19935 17095 19941
rect 16209 19907 16267 19913
rect 16209 19873 16221 19907
rect 16255 19873 16267 19907
rect 16209 19867 16267 19873
rect 16761 19907 16819 19913
rect 16761 19873 16773 19907
rect 16807 19873 16819 19907
rect 16761 19867 16819 19873
rect 9125 19839 9183 19845
rect 9125 19805 9137 19839
rect 9171 19805 9183 19839
rect 10226 19836 10232 19848
rect 10187 19808 10232 19836
rect 9125 19799 9183 19805
rect 10226 19796 10232 19808
rect 10284 19796 10290 19848
rect 10318 19796 10324 19848
rect 10376 19836 10382 19848
rect 10376 19808 10421 19836
rect 10376 19796 10382 19808
rect 12066 19796 12072 19848
rect 12124 19836 12130 19848
rect 15838 19836 15844 19848
rect 12124 19808 12169 19836
rect 15799 19808 15844 19836
rect 12124 19796 12130 19808
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 16224 19836 16252 19867
rect 17218 19864 17224 19916
rect 17276 19904 17282 19916
rect 17497 19907 17555 19913
rect 17497 19904 17509 19907
rect 17276 19876 17509 19904
rect 17276 19864 17282 19876
rect 17497 19873 17509 19876
rect 17543 19873 17555 19907
rect 18325 19907 18383 19913
rect 18325 19904 18337 19907
rect 17497 19867 17555 19873
rect 17604 19876 18337 19904
rect 17236 19836 17264 19864
rect 16224 19808 17264 19836
rect 8938 19728 8944 19780
rect 8996 19768 9002 19780
rect 9769 19771 9827 19777
rect 9769 19768 9781 19771
rect 8996 19740 9781 19768
rect 8996 19728 9002 19740
rect 9769 19737 9781 19740
rect 9815 19737 9827 19771
rect 9769 19731 9827 19737
rect 13446 19728 13452 19780
rect 13504 19768 13510 19780
rect 14093 19771 14151 19777
rect 14093 19768 14105 19771
rect 13504 19740 14105 19768
rect 13504 19728 13510 19740
rect 14093 19737 14105 19740
rect 14139 19737 14151 19771
rect 14093 19731 14151 19737
rect 15197 19771 15255 19777
rect 15197 19737 15209 19771
rect 15243 19768 15255 19771
rect 15286 19768 15292 19780
rect 15243 19740 15292 19768
rect 15243 19737 15255 19740
rect 15197 19731 15255 19737
rect 15286 19728 15292 19740
rect 15344 19728 15350 19780
rect 8297 19703 8355 19709
rect 8297 19700 8309 19703
rect 6380 19672 8309 19700
rect 8297 19669 8309 19672
rect 8343 19669 8355 19703
rect 8297 19663 8355 19669
rect 8573 19703 8631 19709
rect 8573 19669 8585 19703
rect 8619 19700 8631 19703
rect 9674 19700 9680 19712
rect 8619 19672 9680 19700
rect 8619 19669 8631 19672
rect 8573 19663 8631 19669
rect 9674 19660 9680 19672
rect 9732 19660 9738 19712
rect 11517 19703 11575 19709
rect 11517 19669 11529 19703
rect 11563 19700 11575 19703
rect 12802 19700 12808 19712
rect 11563 19672 12808 19700
rect 11563 19669 11575 19672
rect 11517 19663 11575 19669
rect 12802 19660 12808 19672
rect 12860 19660 12866 19712
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 16224 19700 16252 19808
rect 17494 19728 17500 19780
rect 17552 19768 17558 19780
rect 17604 19768 17632 19876
rect 18325 19873 18337 19876
rect 18371 19873 18383 19907
rect 18325 19867 18383 19873
rect 18782 19864 18788 19916
rect 18840 19904 18846 19916
rect 18877 19907 18935 19913
rect 18877 19904 18889 19907
rect 18840 19876 18889 19904
rect 18840 19864 18846 19876
rect 18877 19873 18889 19876
rect 18923 19873 18935 19907
rect 18984 19904 19012 19944
rect 19150 19932 19156 19944
rect 19208 19932 19214 19984
rect 19352 19904 19380 20012
rect 21818 20000 21824 20012
rect 21876 20000 21882 20052
rect 20622 19972 20628 19984
rect 20583 19944 20628 19972
rect 20622 19932 20628 19944
rect 20680 19932 20686 19984
rect 18984 19876 19380 19904
rect 19613 19907 19671 19913
rect 18877 19867 18935 19873
rect 19613 19873 19625 19907
rect 19659 19904 19671 19907
rect 19702 19904 19708 19916
rect 19659 19876 19708 19904
rect 19659 19873 19671 19876
rect 19613 19867 19671 19873
rect 19702 19864 19708 19876
rect 19760 19864 19766 19916
rect 20346 19904 20352 19916
rect 20307 19876 20352 19904
rect 20346 19864 20352 19876
rect 20404 19864 20410 19916
rect 17773 19839 17831 19845
rect 17773 19805 17785 19839
rect 17819 19805 17831 19839
rect 17773 19799 17831 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 22186 19836 22192 19848
rect 19935 19808 22192 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 17552 19740 17632 19768
rect 17788 19768 17816 19799
rect 22186 19796 22192 19808
rect 22244 19796 22250 19848
rect 21450 19768 21456 19780
rect 17788 19740 21456 19768
rect 17552 19728 17558 19740
rect 21450 19728 21456 19740
rect 21508 19728 21514 19780
rect 13872 19672 16252 19700
rect 18509 19703 18567 19709
rect 13872 19660 13878 19672
rect 18509 19669 18521 19703
rect 18555 19700 18567 19703
rect 18874 19700 18880 19712
rect 18555 19672 18880 19700
rect 18555 19669 18567 19672
rect 18509 19663 18567 19669
rect 18874 19660 18880 19672
rect 18932 19660 18938 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 4062 19456 4068 19508
rect 4120 19496 4126 19508
rect 6822 19496 6828 19508
rect 4120 19468 6828 19496
rect 4120 19456 4126 19468
rect 6822 19456 6828 19468
rect 6880 19456 6886 19508
rect 8386 19496 8392 19508
rect 8347 19468 8392 19496
rect 8386 19456 8392 19468
rect 8444 19456 8450 19508
rect 8754 19456 8760 19508
rect 8812 19496 8818 19508
rect 10229 19499 10287 19505
rect 10229 19496 10241 19499
rect 8812 19468 10241 19496
rect 8812 19456 8818 19468
rect 10229 19465 10241 19468
rect 10275 19496 10287 19499
rect 10318 19496 10324 19508
rect 10275 19468 10324 19496
rect 10275 19465 10287 19468
rect 10229 19459 10287 19465
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 15473 19499 15531 19505
rect 12492 19468 12537 19496
rect 12492 19456 12498 19468
rect 15473 19465 15485 19499
rect 15519 19496 15531 19499
rect 15654 19496 15660 19508
rect 15519 19468 15660 19496
rect 15519 19465 15531 19468
rect 15473 19459 15531 19465
rect 15654 19456 15660 19468
rect 15712 19456 15718 19508
rect 16574 19456 16580 19508
rect 16632 19496 16638 19508
rect 19150 19496 19156 19508
rect 16632 19468 19156 19496
rect 16632 19456 16638 19468
rect 19150 19456 19156 19468
rect 19208 19456 19214 19508
rect 14645 19431 14703 19437
rect 3160 19400 4384 19428
rect 3160 19369 3188 19400
rect 3145 19363 3203 19369
rect 3145 19329 3157 19363
rect 3191 19329 3203 19363
rect 3145 19323 3203 19329
rect 3510 19320 3516 19372
rect 3568 19360 3574 19372
rect 4246 19360 4252 19372
rect 3568 19332 4252 19360
rect 3568 19320 3574 19332
rect 4246 19320 4252 19332
rect 4304 19320 4310 19372
rect 4356 19369 4384 19400
rect 14645 19397 14657 19431
rect 14691 19428 14703 19431
rect 16206 19428 16212 19440
rect 14691 19400 16212 19428
rect 14691 19397 14703 19400
rect 14645 19391 14703 19397
rect 16206 19388 16212 19400
rect 16264 19388 16270 19440
rect 4341 19363 4399 19369
rect 4341 19329 4353 19363
rect 4387 19360 4399 19363
rect 4387 19332 4936 19360
rect 4387 19329 4399 19332
rect 4341 19323 4399 19329
rect 1670 19292 1676 19304
rect 1631 19264 1676 19292
rect 1670 19252 1676 19264
rect 1728 19252 1734 19304
rect 1854 19252 1860 19304
rect 1912 19292 1918 19304
rect 1949 19295 2007 19301
rect 1949 19292 1961 19295
rect 1912 19264 1961 19292
rect 1912 19252 1918 19264
rect 1949 19261 1961 19264
rect 1995 19261 2007 19295
rect 1949 19255 2007 19261
rect 2038 19252 2044 19304
rect 2096 19292 2102 19304
rect 2961 19295 3019 19301
rect 2961 19292 2973 19295
rect 2096 19264 2973 19292
rect 2096 19252 2102 19264
rect 2961 19261 2973 19264
rect 3007 19292 3019 19295
rect 4062 19292 4068 19304
rect 3007 19264 4068 19292
rect 3007 19261 3019 19264
rect 2961 19255 3019 19261
rect 4062 19252 4068 19264
rect 4120 19252 4126 19304
rect 4154 19252 4160 19304
rect 4212 19292 4218 19304
rect 4808 19295 4866 19301
rect 4808 19292 4820 19295
rect 4212 19264 4820 19292
rect 4212 19252 4218 19264
rect 4808 19261 4820 19264
rect 4854 19261 4866 19295
rect 4808 19255 4866 19261
rect 1302 19184 1308 19236
rect 1360 19224 1366 19236
rect 4249 19227 4307 19233
rect 4249 19224 4261 19227
rect 1360 19196 4261 19224
rect 1360 19184 1366 19196
rect 4249 19193 4261 19196
rect 4295 19224 4307 19227
rect 4338 19224 4344 19236
rect 4295 19196 4344 19224
rect 4295 19193 4307 19196
rect 4249 19187 4307 19193
rect 4338 19184 4344 19196
rect 4396 19184 4402 19236
rect 4908 19224 4936 19332
rect 6638 19320 6644 19372
rect 6696 19360 6702 19372
rect 7009 19363 7067 19369
rect 7009 19360 7021 19363
rect 6696 19332 7021 19360
rect 6696 19320 6702 19332
rect 7009 19329 7021 19332
rect 7055 19329 7067 19363
rect 7009 19323 7067 19329
rect 8018 19320 8024 19372
rect 8076 19360 8082 19372
rect 8076 19332 8340 19360
rect 8076 19320 8082 19332
rect 5068 19295 5126 19301
rect 5068 19261 5080 19295
rect 5114 19292 5126 19295
rect 5350 19292 5356 19304
rect 5114 19264 5356 19292
rect 5114 19261 5126 19264
rect 5068 19255 5126 19261
rect 5350 19252 5356 19264
rect 5408 19252 5414 19304
rect 8312 19292 8340 19332
rect 10134 19320 10140 19372
rect 10192 19360 10198 19372
rect 10318 19360 10324 19372
rect 10192 19332 10324 19360
rect 10192 19320 10198 19332
rect 10318 19320 10324 19332
rect 10376 19320 10382 19372
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19360 12035 19363
rect 12066 19360 12072 19372
rect 12023 19332 12072 19360
rect 12023 19329 12035 19332
rect 11977 19323 12035 19329
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 13081 19363 13139 19369
rect 13081 19329 13093 19363
rect 13127 19360 13139 19363
rect 13630 19360 13636 19372
rect 13127 19332 13636 19360
rect 13127 19329 13139 19332
rect 13081 19323 13139 19329
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 14277 19363 14335 19369
rect 14277 19329 14289 19363
rect 14323 19360 14335 19363
rect 15102 19360 15108 19372
rect 14323 19332 15108 19360
rect 14323 19329 14335 19332
rect 14277 19323 14335 19329
rect 15102 19320 15108 19332
rect 15160 19360 15166 19372
rect 15197 19363 15255 19369
rect 15197 19360 15209 19363
rect 15160 19332 15209 19360
rect 15160 19320 15166 19332
rect 15197 19329 15209 19332
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 15930 19320 15936 19372
rect 15988 19360 15994 19372
rect 16025 19363 16083 19369
rect 16025 19360 16037 19363
rect 15988 19332 16037 19360
rect 15988 19320 15994 19332
rect 16025 19329 16037 19332
rect 16071 19329 16083 19363
rect 18598 19360 18604 19372
rect 16025 19323 16083 19329
rect 17880 19332 18604 19360
rect 8849 19295 8907 19301
rect 8849 19292 8861 19295
rect 8312 19264 8861 19292
rect 8849 19261 8861 19264
rect 8895 19261 8907 19295
rect 9398 19292 9404 19304
rect 8849 19255 8907 19261
rect 9048 19264 9404 19292
rect 7276 19227 7334 19233
rect 4908 19196 6224 19224
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2774 19156 2780 19168
rect 2547 19128 2780 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2774 19116 2780 19128
rect 2832 19116 2838 19168
rect 2869 19159 2927 19165
rect 2869 19125 2881 19159
rect 2915 19156 2927 19159
rect 2958 19156 2964 19168
rect 2915 19128 2964 19156
rect 2915 19125 2927 19128
rect 2869 19119 2927 19125
rect 2958 19116 2964 19128
rect 3016 19156 3022 19168
rect 3510 19156 3516 19168
rect 3016 19128 3516 19156
rect 3016 19116 3022 19128
rect 3510 19116 3516 19128
rect 3568 19116 3574 19168
rect 3786 19156 3792 19168
rect 3747 19128 3792 19156
rect 3786 19116 3792 19128
rect 3844 19116 3850 19168
rect 4157 19159 4215 19165
rect 4157 19125 4169 19159
rect 4203 19156 4215 19159
rect 4890 19156 4896 19168
rect 4203 19128 4896 19156
rect 4203 19125 4215 19128
rect 4157 19119 4215 19125
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 5166 19116 5172 19168
rect 5224 19156 5230 19168
rect 5350 19156 5356 19168
rect 5224 19128 5356 19156
rect 5224 19116 5230 19128
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 6196 19165 6224 19196
rect 7276 19193 7288 19227
rect 7322 19224 7334 19227
rect 7742 19224 7748 19236
rect 7322 19196 7748 19224
rect 7322 19193 7334 19196
rect 7276 19187 7334 19193
rect 7742 19184 7748 19196
rect 7800 19184 7806 19236
rect 8110 19184 8116 19236
rect 8168 19224 8174 19236
rect 9048 19224 9076 19264
rect 9398 19252 9404 19264
rect 9456 19252 9462 19304
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 10505 19295 10563 19301
rect 10505 19292 10517 19295
rect 9732 19264 10517 19292
rect 9732 19252 9738 19264
rect 10505 19261 10517 19264
rect 10551 19261 10563 19295
rect 10505 19255 10563 19261
rect 11793 19295 11851 19301
rect 11793 19261 11805 19295
rect 11839 19292 11851 19295
rect 12526 19292 12532 19304
rect 11839 19264 12532 19292
rect 11839 19261 11851 19264
rect 11793 19255 11851 19261
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 14001 19295 14059 19301
rect 14001 19261 14013 19295
rect 14047 19292 14059 19295
rect 14918 19292 14924 19304
rect 14047 19264 14924 19292
rect 14047 19261 14059 19264
rect 14001 19255 14059 19261
rect 14918 19252 14924 19264
rect 14976 19252 14982 19304
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 16485 19295 16543 19301
rect 15059 19264 16436 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 8168 19196 9076 19224
rect 9116 19227 9174 19233
rect 8168 19184 8174 19196
rect 9116 19193 9128 19227
rect 9162 19224 9174 19227
rect 9214 19224 9220 19236
rect 9162 19196 9220 19224
rect 9162 19193 9174 19196
rect 9116 19187 9174 19193
rect 9214 19184 9220 19196
rect 9272 19184 9278 19236
rect 9950 19184 9956 19236
rect 10008 19224 10014 19236
rect 10781 19227 10839 19233
rect 10781 19224 10793 19227
rect 10008 19196 10793 19224
rect 10008 19184 10014 19196
rect 10781 19193 10793 19196
rect 10827 19193 10839 19227
rect 10781 19187 10839 19193
rect 11701 19227 11759 19233
rect 11701 19193 11713 19227
rect 11747 19224 11759 19227
rect 12805 19227 12863 19233
rect 11747 19196 12112 19224
rect 11747 19193 11759 19196
rect 11701 19187 11759 19193
rect 6181 19159 6239 19165
rect 6181 19125 6193 19159
rect 6227 19156 6239 19159
rect 6270 19156 6276 19168
rect 6227 19128 6276 19156
rect 6227 19125 6239 19128
rect 6181 19119 6239 19125
rect 6270 19116 6276 19128
rect 6328 19116 6334 19168
rect 6454 19116 6460 19168
rect 6512 19156 6518 19168
rect 10042 19156 10048 19168
rect 6512 19128 10048 19156
rect 6512 19116 6518 19128
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 11333 19159 11391 19165
rect 11333 19125 11345 19159
rect 11379 19156 11391 19159
rect 11790 19156 11796 19168
rect 11379 19128 11796 19156
rect 11379 19125 11391 19128
rect 11333 19119 11391 19125
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 12084 19156 12112 19196
rect 12805 19193 12817 19227
rect 12851 19224 12863 19227
rect 14274 19224 14280 19236
rect 12851 19196 14280 19224
rect 12851 19193 12863 19196
rect 12805 19187 12863 19193
rect 14274 19184 14280 19196
rect 14332 19184 14338 19236
rect 15105 19227 15163 19233
rect 15105 19193 15117 19227
rect 15151 19224 15163 19227
rect 16114 19224 16120 19236
rect 15151 19196 16120 19224
rect 15151 19193 15163 19196
rect 15105 19187 15163 19193
rect 16114 19184 16120 19196
rect 16172 19184 16178 19236
rect 16408 19224 16436 19264
rect 16485 19261 16497 19295
rect 16531 19292 16543 19295
rect 16574 19292 16580 19304
rect 16531 19264 16580 19292
rect 16531 19261 16543 19264
rect 16485 19255 16543 19261
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 17218 19292 17224 19304
rect 17179 19264 17224 19292
rect 17218 19252 17224 19264
rect 17276 19252 17282 19304
rect 17880 19292 17908 19332
rect 18598 19320 18604 19332
rect 18656 19320 18662 19372
rect 18966 19360 18972 19372
rect 18927 19332 18972 19360
rect 18966 19320 18972 19332
rect 19024 19320 19030 19372
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 19392 19332 20484 19360
rect 19392 19320 19398 19332
rect 17420 19264 17908 19292
rect 16666 19224 16672 19236
rect 16408 19196 16672 19224
rect 16666 19184 16672 19196
rect 16724 19184 16730 19236
rect 16761 19227 16819 19233
rect 16761 19193 16773 19227
rect 16807 19224 16819 19227
rect 17420 19224 17448 19264
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 18012 19264 18061 19292
rect 18012 19252 18018 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18138 19252 18144 19304
rect 18196 19292 18202 19304
rect 18785 19295 18843 19301
rect 18196 19264 18736 19292
rect 18196 19252 18202 19264
rect 16807 19196 17448 19224
rect 17497 19227 17555 19233
rect 16807 19193 16819 19196
rect 16761 19187 16819 19193
rect 17497 19193 17509 19227
rect 17543 19224 17555 19227
rect 18506 19224 18512 19236
rect 17543 19196 18512 19224
rect 17543 19193 17555 19196
rect 17497 19187 17555 19193
rect 18506 19184 18512 19196
rect 18564 19184 18570 19236
rect 18708 19224 18736 19264
rect 18785 19261 18797 19295
rect 18831 19292 18843 19295
rect 19794 19292 19800 19304
rect 18831 19264 19800 19292
rect 18831 19261 18843 19264
rect 18785 19255 18843 19261
rect 19794 19252 19800 19264
rect 19852 19252 19858 19304
rect 20456 19301 20484 19332
rect 19889 19295 19947 19301
rect 19889 19261 19901 19295
rect 19935 19261 19947 19295
rect 19889 19255 19947 19261
rect 20441 19295 20499 19301
rect 20441 19261 20453 19295
rect 20487 19261 20499 19295
rect 20441 19255 20499 19261
rect 20717 19295 20775 19301
rect 20717 19261 20729 19295
rect 20763 19292 20775 19295
rect 20806 19292 20812 19304
rect 20763 19264 20812 19292
rect 20763 19261 20775 19264
rect 20717 19255 20775 19261
rect 19518 19224 19524 19236
rect 18708 19196 19524 19224
rect 19518 19184 19524 19196
rect 19576 19184 19582 19236
rect 12710 19156 12716 19168
rect 12084 19128 12716 19156
rect 12710 19116 12716 19128
rect 12768 19116 12774 19168
rect 12897 19159 12955 19165
rect 12897 19125 12909 19159
rect 12943 19156 12955 19159
rect 13446 19156 13452 19168
rect 12943 19128 13452 19156
rect 12943 19125 12955 19128
rect 12897 19119 12955 19125
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 13538 19116 13544 19168
rect 13596 19156 13602 19168
rect 13633 19159 13691 19165
rect 13633 19156 13645 19159
rect 13596 19128 13645 19156
rect 13596 19116 13602 19128
rect 13633 19125 13645 19128
rect 13679 19125 13691 19159
rect 14090 19156 14096 19168
rect 14051 19128 14096 19156
rect 13633 19119 13691 19125
rect 14090 19116 14096 19128
rect 14148 19116 14154 19168
rect 15010 19116 15016 19168
rect 15068 19156 15074 19168
rect 15841 19159 15899 19165
rect 15841 19156 15853 19159
rect 15068 19128 15853 19156
rect 15068 19116 15074 19128
rect 15841 19125 15853 19128
rect 15887 19125 15899 19159
rect 15841 19119 15899 19125
rect 15930 19116 15936 19168
rect 15988 19156 15994 19168
rect 15988 19128 16033 19156
rect 15988 19116 15994 19128
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 17770 19156 17776 19168
rect 16448 19128 17776 19156
rect 16448 19116 16454 19128
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18966 19156 18972 19168
rect 18279 19128 18972 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18966 19116 18972 19128
rect 19024 19116 19030 19168
rect 19426 19116 19432 19168
rect 19484 19156 19490 19168
rect 19904 19156 19932 19255
rect 20806 19252 20812 19264
rect 20864 19252 20870 19304
rect 19484 19128 19932 19156
rect 20073 19159 20131 19165
rect 19484 19116 19490 19128
rect 20073 19125 20085 19159
rect 20119 19156 20131 19159
rect 20162 19156 20168 19168
rect 20119 19128 20168 19156
rect 20119 19125 20131 19128
rect 20073 19119 20131 19125
rect 20162 19116 20168 19128
rect 20220 19116 20226 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 2961 18955 3019 18961
rect 2961 18921 2973 18955
rect 3007 18952 3019 18955
rect 4706 18952 4712 18964
rect 3007 18924 4712 18952
rect 3007 18921 3019 18924
rect 2961 18915 3019 18921
rect 4706 18912 4712 18924
rect 4764 18912 4770 18964
rect 4798 18912 4804 18964
rect 4856 18952 4862 18964
rect 5810 18952 5816 18964
rect 4856 18924 5816 18952
rect 4856 18912 4862 18924
rect 5810 18912 5816 18924
rect 5868 18912 5874 18964
rect 6178 18952 6184 18964
rect 6139 18924 6184 18952
rect 6178 18912 6184 18924
rect 6236 18912 6242 18964
rect 9677 18955 9735 18961
rect 6288 18924 8984 18952
rect 1946 18884 1952 18896
rect 1907 18856 1952 18884
rect 1946 18844 1952 18856
rect 2004 18844 2010 18896
rect 3329 18887 3387 18893
rect 3329 18853 3341 18887
rect 3375 18884 3387 18887
rect 5074 18884 5080 18896
rect 3375 18856 5080 18884
rect 3375 18853 3387 18856
rect 3329 18847 3387 18853
rect 5074 18844 5080 18856
rect 5132 18844 5138 18896
rect 5718 18844 5724 18896
rect 5776 18884 5782 18896
rect 6288 18884 6316 18924
rect 5776 18856 6316 18884
rect 7009 18887 7067 18893
rect 5776 18844 5782 18856
rect 7009 18853 7021 18887
rect 7055 18884 7067 18887
rect 8846 18884 8852 18896
rect 7055 18856 8852 18884
rect 7055 18853 7067 18856
rect 7009 18847 7067 18853
rect 8846 18844 8852 18856
rect 8904 18844 8910 18896
rect 1673 18819 1731 18825
rect 1673 18785 1685 18819
rect 1719 18785 1731 18819
rect 1673 18779 1731 18785
rect 1688 18680 1716 18779
rect 2314 18776 2320 18828
rect 2372 18816 2378 18828
rect 2409 18819 2467 18825
rect 2409 18816 2421 18819
rect 2372 18788 2421 18816
rect 2372 18776 2378 18788
rect 2409 18785 2421 18788
rect 2455 18785 2467 18819
rect 4065 18819 4123 18825
rect 4065 18816 4077 18819
rect 2409 18779 2467 18785
rect 3252 18788 4077 18816
rect 2222 18708 2228 18760
rect 2280 18748 2286 18760
rect 3252 18748 3280 18788
rect 4065 18785 4077 18788
rect 4111 18816 4123 18819
rect 4154 18816 4160 18828
rect 4111 18788 4160 18816
rect 4111 18785 4123 18788
rect 4065 18779 4123 18785
rect 4154 18776 4160 18788
rect 4212 18776 4218 18828
rect 4332 18819 4390 18825
rect 4332 18785 4344 18819
rect 4378 18816 4390 18819
rect 4798 18816 4804 18828
rect 4378 18788 4804 18816
rect 4378 18785 4390 18788
rect 4332 18779 4390 18785
rect 4798 18776 4804 18788
rect 4856 18776 4862 18828
rect 6086 18816 6092 18828
rect 6047 18788 6092 18816
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 6733 18819 6791 18825
rect 6733 18785 6745 18819
rect 6779 18816 6791 18819
rect 7374 18816 7380 18828
rect 6779 18788 7380 18816
rect 6779 18785 6791 18788
rect 6733 18779 6791 18785
rect 7374 18776 7380 18788
rect 7432 18776 7438 18828
rect 7736 18819 7794 18825
rect 7736 18785 7748 18819
rect 7782 18816 7794 18819
rect 8754 18816 8760 18828
rect 7782 18788 8760 18816
rect 7782 18785 7794 18788
rect 7736 18779 7794 18785
rect 8754 18776 8760 18788
rect 8812 18776 8818 18828
rect 8956 18816 8984 18924
rect 9677 18921 9689 18955
rect 9723 18952 9735 18955
rect 10226 18952 10232 18964
rect 9723 18924 10232 18952
rect 9723 18921 9735 18924
rect 9677 18915 9735 18921
rect 10226 18912 10232 18924
rect 10284 18912 10290 18964
rect 12805 18955 12863 18961
rect 12805 18921 12817 18955
rect 12851 18921 12863 18955
rect 12805 18915 12863 18921
rect 9398 18844 9404 18896
rect 9456 18884 9462 18896
rect 10042 18884 10048 18896
rect 9456 18856 9904 18884
rect 10003 18856 10048 18884
rect 9456 18844 9462 18856
rect 9674 18816 9680 18828
rect 8956 18788 9680 18816
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 9876 18816 9904 18856
rect 10042 18844 10048 18856
rect 10100 18844 10106 18896
rect 12820 18884 12848 18915
rect 14274 18912 14280 18964
rect 14332 18952 14338 18964
rect 14737 18955 14795 18961
rect 14737 18952 14749 18955
rect 14332 18924 14749 18952
rect 14332 18912 14338 18924
rect 14737 18921 14749 18924
rect 14783 18921 14795 18955
rect 14737 18915 14795 18921
rect 15286 18912 15292 18964
rect 15344 18952 15350 18964
rect 15470 18952 15476 18964
rect 15344 18924 15476 18952
rect 15344 18912 15350 18924
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 16206 18912 16212 18964
rect 16264 18952 16270 18964
rect 19978 18952 19984 18964
rect 16264 18924 19984 18952
rect 16264 18912 16270 18924
rect 19978 18912 19984 18924
rect 20036 18912 20042 18964
rect 12986 18884 12992 18896
rect 12820 18856 12992 18884
rect 12986 18844 12992 18856
rect 13044 18884 13050 18896
rect 13326 18887 13384 18893
rect 13326 18884 13338 18887
rect 13044 18856 13338 18884
rect 13044 18844 13050 18856
rect 13326 18853 13338 18856
rect 13372 18853 13384 18887
rect 13326 18847 13384 18853
rect 14090 18844 14096 18896
rect 14148 18884 14154 18896
rect 17126 18884 17132 18896
rect 14148 18856 17132 18884
rect 14148 18844 14154 18856
rect 17126 18844 17132 18856
rect 17184 18844 17190 18896
rect 18138 18844 18144 18896
rect 18196 18884 18202 18896
rect 18196 18856 18241 18884
rect 18524 18856 19196 18884
rect 18196 18844 18202 18856
rect 10594 18816 10600 18828
rect 9876 18788 10600 18816
rect 10594 18776 10600 18788
rect 10652 18776 10658 18828
rect 10689 18819 10747 18825
rect 10689 18785 10701 18819
rect 10735 18816 10747 18819
rect 11514 18816 11520 18828
rect 10735 18788 11520 18816
rect 10735 18785 10747 18788
rect 10689 18779 10747 18785
rect 11514 18776 11520 18788
rect 11572 18776 11578 18828
rect 11692 18819 11750 18825
rect 11692 18785 11704 18819
rect 11738 18816 11750 18819
rect 12066 18816 12072 18828
rect 11738 18788 12072 18816
rect 11738 18785 11750 18788
rect 11692 18779 11750 18785
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 12250 18776 12256 18828
rect 12308 18816 12314 18828
rect 16669 18819 16727 18825
rect 16669 18816 16681 18819
rect 12308 18788 16681 18816
rect 12308 18776 12314 18788
rect 16669 18785 16681 18788
rect 16715 18785 16727 18819
rect 16669 18779 16727 18785
rect 17218 18776 17224 18828
rect 17276 18816 17282 18828
rect 17313 18819 17371 18825
rect 17313 18816 17325 18819
rect 17276 18788 17325 18816
rect 17276 18776 17282 18788
rect 17313 18785 17325 18788
rect 17359 18785 17371 18819
rect 17313 18779 17371 18785
rect 17770 18776 17776 18828
rect 17828 18816 17834 18828
rect 17865 18819 17923 18825
rect 17865 18816 17877 18819
rect 17828 18788 17877 18816
rect 17828 18776 17834 18788
rect 17865 18785 17877 18788
rect 17911 18816 17923 18819
rect 18524 18816 18552 18856
rect 17911 18788 18552 18816
rect 18601 18819 18659 18825
rect 17911 18785 17923 18788
rect 17865 18779 17923 18785
rect 18601 18785 18613 18819
rect 18647 18816 18659 18819
rect 18690 18816 18696 18828
rect 18647 18788 18696 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 18690 18776 18696 18788
rect 18748 18776 18754 18828
rect 18877 18819 18935 18825
rect 18877 18785 18889 18819
rect 18923 18816 18935 18819
rect 19061 18819 19119 18825
rect 19061 18816 19073 18819
rect 18923 18788 19073 18816
rect 18923 18785 18935 18788
rect 18877 18779 18935 18785
rect 19061 18785 19073 18788
rect 19107 18785 19119 18819
rect 19061 18779 19119 18785
rect 3418 18748 3424 18760
rect 2280 18720 3280 18748
rect 3379 18720 3424 18748
rect 2280 18708 2286 18720
rect 3418 18708 3424 18720
rect 3476 18708 3482 18760
rect 3605 18751 3663 18757
rect 3605 18717 3617 18751
rect 3651 18717 3663 18751
rect 3605 18711 3663 18717
rect 3510 18680 3516 18692
rect 1688 18652 3516 18680
rect 3510 18640 3516 18652
rect 3568 18640 3574 18692
rect 2593 18615 2651 18621
rect 2593 18581 2605 18615
rect 2639 18612 2651 18615
rect 2774 18612 2780 18624
rect 2639 18584 2780 18612
rect 2639 18581 2651 18584
rect 2593 18575 2651 18581
rect 2774 18572 2780 18584
rect 2832 18572 2838 18624
rect 3620 18612 3648 18711
rect 5166 18708 5172 18760
rect 5224 18748 5230 18760
rect 6270 18748 6276 18760
rect 5224 18720 6276 18748
rect 5224 18708 5230 18720
rect 6270 18708 6276 18720
rect 6328 18708 6334 18760
rect 6638 18708 6644 18760
rect 6696 18748 6702 18760
rect 7469 18751 7527 18757
rect 7469 18748 7481 18751
rect 6696 18720 7481 18748
rect 6696 18708 6702 18720
rect 7469 18717 7481 18720
rect 7515 18717 7527 18751
rect 9122 18748 9128 18760
rect 9083 18720 9128 18748
rect 7469 18711 7527 18717
rect 9122 18708 9128 18720
rect 9180 18708 9186 18760
rect 10042 18748 10048 18760
rect 9232 18720 10048 18748
rect 8478 18640 8484 18692
rect 8536 18680 8542 18692
rect 9232 18680 9260 18720
rect 10042 18708 10048 18720
rect 10100 18748 10106 18760
rect 10137 18751 10195 18757
rect 10137 18748 10149 18751
rect 10100 18720 10149 18748
rect 10100 18708 10106 18720
rect 10137 18717 10149 18720
rect 10183 18717 10195 18751
rect 10137 18711 10195 18717
rect 10229 18751 10287 18757
rect 10229 18717 10241 18751
rect 10275 18717 10287 18751
rect 10229 18711 10287 18717
rect 10965 18751 11023 18757
rect 10965 18717 10977 18751
rect 11011 18748 11023 18751
rect 11146 18748 11152 18760
rect 11011 18720 11152 18748
rect 11011 18717 11023 18720
rect 10965 18711 11023 18717
rect 10244 18680 10272 18711
rect 11146 18708 11152 18720
rect 11204 18708 11210 18760
rect 11425 18751 11483 18757
rect 11425 18717 11437 18751
rect 11471 18717 11483 18751
rect 11425 18711 11483 18717
rect 8536 18652 9260 18680
rect 9416 18652 10272 18680
rect 8536 18640 8542 18652
rect 5350 18612 5356 18624
rect 3620 18584 5356 18612
rect 5350 18572 5356 18584
rect 5408 18612 5414 18624
rect 5445 18615 5503 18621
rect 5445 18612 5457 18615
rect 5408 18584 5457 18612
rect 5408 18572 5414 18584
rect 5445 18581 5457 18584
rect 5491 18581 5503 18615
rect 5718 18612 5724 18624
rect 5679 18584 5724 18612
rect 5445 18575 5503 18581
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 5902 18572 5908 18624
rect 5960 18612 5966 18624
rect 7282 18612 7288 18624
rect 5960 18584 7288 18612
rect 5960 18572 5966 18584
rect 7282 18572 7288 18584
rect 7340 18572 7346 18624
rect 7742 18572 7748 18624
rect 7800 18612 7806 18624
rect 8849 18615 8907 18621
rect 8849 18612 8861 18615
rect 7800 18584 8861 18612
rect 7800 18572 7806 18584
rect 8849 18581 8861 18584
rect 8895 18581 8907 18615
rect 8849 18575 8907 18581
rect 9214 18572 9220 18624
rect 9272 18612 9278 18624
rect 9416 18612 9444 18652
rect 10594 18640 10600 18692
rect 10652 18680 10658 18692
rect 11440 18680 11468 18711
rect 12894 18708 12900 18760
rect 12952 18748 12958 18760
rect 13081 18751 13139 18757
rect 13081 18748 13093 18751
rect 12952 18720 13093 18748
rect 12952 18708 12958 18720
rect 13081 18717 13093 18720
rect 13127 18717 13139 18751
rect 16761 18751 16819 18757
rect 16761 18748 16773 18751
rect 13081 18711 13139 18717
rect 16224 18720 16773 18748
rect 10652 18652 11468 18680
rect 10652 18640 10658 18652
rect 16224 18624 16252 18720
rect 16761 18717 16773 18720
rect 16807 18717 16819 18751
rect 16761 18711 16819 18717
rect 16945 18751 17003 18757
rect 16945 18717 16957 18751
rect 16991 18748 17003 18751
rect 16991 18720 19104 18748
rect 16991 18717 17003 18720
rect 16945 18711 17003 18717
rect 16301 18683 16359 18689
rect 16301 18649 16313 18683
rect 16347 18680 16359 18683
rect 16347 18652 19012 18680
rect 16347 18649 16359 18652
rect 16301 18643 16359 18649
rect 18984 18624 19012 18652
rect 9272 18584 9444 18612
rect 9272 18572 9278 18584
rect 9582 18572 9588 18624
rect 9640 18612 9646 18624
rect 13814 18612 13820 18624
rect 9640 18584 13820 18612
rect 9640 18572 9646 18584
rect 13814 18572 13820 18584
rect 13872 18572 13878 18624
rect 14090 18572 14096 18624
rect 14148 18612 14154 18624
rect 14461 18615 14519 18621
rect 14461 18612 14473 18615
rect 14148 18584 14473 18612
rect 14148 18572 14154 18584
rect 14461 18581 14473 18584
rect 14507 18581 14519 18615
rect 16206 18612 16212 18624
rect 16167 18584 16212 18612
rect 14461 18575 14519 18581
rect 16206 18572 16212 18584
rect 16264 18572 16270 18624
rect 17497 18615 17555 18621
rect 17497 18581 17509 18615
rect 17543 18612 17555 18615
rect 17954 18612 17960 18624
rect 17543 18584 17960 18612
rect 17543 18581 17555 18584
rect 17497 18575 17555 18581
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 18966 18572 18972 18624
rect 19024 18572 19030 18624
rect 19076 18612 19104 18720
rect 19168 18680 19196 18856
rect 19242 18844 19248 18896
rect 19300 18884 19306 18896
rect 20349 18887 20407 18893
rect 20349 18884 20361 18887
rect 19300 18856 20361 18884
rect 19300 18844 19306 18856
rect 20349 18853 20361 18856
rect 20395 18853 20407 18887
rect 20349 18847 20407 18853
rect 19334 18816 19340 18828
rect 19295 18788 19340 18816
rect 19334 18776 19340 18788
rect 19392 18776 19398 18828
rect 19702 18776 19708 18828
rect 19760 18816 19766 18828
rect 20073 18819 20131 18825
rect 20073 18816 20085 18819
rect 19760 18788 20085 18816
rect 19760 18776 19766 18788
rect 20073 18785 20085 18788
rect 20119 18785 20131 18819
rect 20073 18779 20131 18785
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 19613 18751 19671 18757
rect 19300 18720 19345 18748
rect 19300 18708 19306 18720
rect 19613 18717 19625 18751
rect 19659 18748 19671 18751
rect 22554 18748 22560 18760
rect 19659 18720 22560 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 22554 18708 22560 18720
rect 22612 18708 22618 18760
rect 20346 18680 20352 18692
rect 19168 18652 20352 18680
rect 20346 18640 20352 18652
rect 20404 18640 20410 18692
rect 20898 18612 20904 18624
rect 19076 18584 20904 18612
rect 20898 18572 20904 18584
rect 20956 18572 20962 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 5718 18408 5724 18420
rect 4540 18380 5724 18408
rect 4430 18340 4436 18352
rect 3436 18312 4436 18340
rect 2222 18232 2228 18284
rect 2280 18272 2286 18284
rect 2409 18275 2467 18281
rect 2409 18272 2421 18275
rect 2280 18244 2421 18272
rect 2280 18232 2286 18244
rect 2409 18241 2421 18244
rect 2455 18241 2467 18275
rect 2409 18235 2467 18241
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18204 1823 18207
rect 3436 18204 3464 18312
rect 4430 18300 4436 18312
rect 4488 18300 4494 18352
rect 3510 18232 3516 18284
rect 3568 18272 3574 18284
rect 4540 18281 4568 18380
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 5994 18368 6000 18420
rect 6052 18408 6058 18420
rect 7009 18411 7067 18417
rect 7009 18408 7021 18411
rect 6052 18380 7021 18408
rect 6052 18368 6058 18380
rect 7009 18377 7021 18380
rect 7055 18377 7067 18411
rect 7009 18371 7067 18377
rect 7469 18411 7527 18417
rect 7469 18377 7481 18411
rect 7515 18408 7527 18411
rect 7650 18408 7656 18420
rect 7515 18380 7656 18408
rect 7515 18377 7527 18380
rect 7469 18371 7527 18377
rect 7650 18368 7656 18380
rect 7708 18368 7714 18420
rect 8481 18411 8539 18417
rect 8481 18377 8493 18411
rect 8527 18408 8539 18411
rect 9030 18408 9036 18420
rect 8527 18380 9036 18408
rect 8527 18377 8539 18380
rect 8481 18371 8539 18377
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 9490 18408 9496 18420
rect 9451 18380 9496 18408
rect 9490 18368 9496 18380
rect 9548 18368 9554 18420
rect 9582 18368 9588 18420
rect 9640 18368 9646 18420
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 10042 18408 10048 18420
rect 9732 18380 10048 18408
rect 9732 18368 9738 18380
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 12066 18408 12072 18420
rect 12027 18380 12072 18408
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 12437 18411 12495 18417
rect 12437 18377 12449 18411
rect 12483 18408 12495 18411
rect 12618 18408 12624 18420
rect 12483 18380 12624 18408
rect 12483 18377 12495 18380
rect 12437 18371 12495 18377
rect 12618 18368 12624 18380
rect 12676 18368 12682 18420
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 13449 18411 13507 18417
rect 13449 18408 13461 18411
rect 12768 18380 13461 18408
rect 12768 18368 12774 18380
rect 13449 18377 13461 18380
rect 13495 18377 13507 18411
rect 13449 18371 13507 18377
rect 15105 18411 15163 18417
rect 15105 18377 15117 18411
rect 15151 18408 15163 18411
rect 15930 18408 15936 18420
rect 15151 18380 15936 18408
rect 15151 18377 15163 18380
rect 15105 18371 15163 18377
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 16114 18408 16120 18420
rect 16075 18380 16120 18408
rect 16114 18368 16120 18380
rect 16172 18368 16178 18420
rect 18690 18408 18696 18420
rect 17328 18380 18696 18408
rect 9600 18340 9628 18368
rect 8036 18312 9076 18340
rect 4525 18275 4583 18281
rect 3568 18244 4476 18272
rect 3568 18232 3574 18244
rect 1811 18176 3464 18204
rect 1811 18173 1823 18176
rect 1765 18167 1823 18173
rect 3786 18164 3792 18216
rect 3844 18204 3850 18216
rect 4338 18204 4344 18216
rect 3844 18176 4344 18204
rect 3844 18164 3850 18176
rect 4338 18164 4344 18176
rect 4396 18164 4402 18216
rect 4448 18204 4476 18244
rect 4525 18241 4537 18275
rect 4571 18241 4583 18275
rect 4706 18272 4712 18284
rect 4667 18244 4712 18272
rect 4525 18235 4583 18241
rect 4706 18232 4712 18244
rect 4764 18232 4770 18284
rect 6288 18244 6868 18272
rect 5350 18213 5356 18216
rect 4985 18207 5043 18213
rect 4448 18176 4936 18204
rect 2676 18139 2734 18145
rect 2676 18105 2688 18139
rect 2722 18136 2734 18139
rect 2958 18136 2964 18148
rect 2722 18108 2964 18136
rect 2722 18105 2734 18108
rect 2676 18099 2734 18105
rect 2958 18096 2964 18108
rect 3016 18096 3022 18148
rect 4522 18136 4528 18148
rect 3804 18108 4528 18136
rect 3804 18077 3832 18108
rect 4522 18096 4528 18108
rect 4580 18136 4586 18148
rect 4798 18136 4804 18148
rect 4580 18108 4804 18136
rect 4580 18096 4586 18108
rect 4798 18096 4804 18108
rect 4856 18096 4862 18148
rect 4908 18136 4936 18176
rect 4985 18173 4997 18207
rect 5031 18204 5043 18207
rect 5077 18207 5135 18213
rect 5077 18204 5089 18207
rect 5031 18176 5089 18204
rect 5031 18173 5043 18176
rect 4985 18167 5043 18173
rect 5077 18173 5089 18176
rect 5123 18173 5135 18207
rect 5344 18204 5356 18213
rect 5311 18176 5356 18204
rect 5077 18167 5135 18173
rect 5344 18167 5356 18176
rect 5350 18164 5356 18167
rect 5408 18164 5414 18216
rect 6288 18136 6316 18244
rect 6840 18213 6868 18244
rect 7742 18232 7748 18284
rect 7800 18272 7806 18284
rect 8036 18281 8064 18312
rect 8021 18275 8079 18281
rect 8021 18272 8033 18275
rect 7800 18244 8033 18272
rect 7800 18232 7806 18244
rect 8021 18241 8033 18244
rect 8067 18241 8079 18275
rect 8938 18272 8944 18284
rect 8899 18244 8944 18272
rect 8021 18235 8079 18241
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 9048 18281 9076 18312
rect 9140 18312 9628 18340
rect 12360 18312 13676 18340
rect 9033 18275 9091 18281
rect 9033 18241 9045 18275
rect 9079 18241 9091 18275
rect 9033 18235 9091 18241
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18204 6883 18207
rect 9140 18204 9168 18312
rect 9214 18232 9220 18284
rect 9272 18272 9278 18284
rect 10045 18275 10103 18281
rect 10045 18272 10057 18275
rect 9272 18244 10057 18272
rect 9272 18232 9278 18244
rect 9600 18216 9628 18244
rect 10045 18241 10057 18244
rect 10091 18241 10103 18275
rect 10045 18235 10103 18241
rect 6871 18176 9168 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 9582 18164 9588 18216
rect 9640 18164 9646 18216
rect 9766 18164 9772 18216
rect 9824 18204 9830 18216
rect 9861 18207 9919 18213
rect 9861 18204 9873 18207
rect 9824 18176 9873 18204
rect 9824 18164 9830 18176
rect 9861 18173 9873 18176
rect 9907 18204 9919 18207
rect 10318 18204 10324 18216
rect 9907 18176 10324 18204
rect 9907 18173 9919 18176
rect 9861 18167 9919 18173
rect 10318 18164 10324 18176
rect 10376 18164 10382 18216
rect 10594 18164 10600 18216
rect 10652 18204 10658 18216
rect 10689 18207 10747 18213
rect 10689 18204 10701 18207
rect 10652 18176 10701 18204
rect 10652 18164 10658 18176
rect 10689 18173 10701 18176
rect 10735 18173 10747 18207
rect 10689 18167 10747 18173
rect 10956 18207 11014 18213
rect 10956 18173 10968 18207
rect 11002 18204 11014 18207
rect 12360 18204 12388 18312
rect 13648 18284 13676 18312
rect 13906 18300 13912 18352
rect 13964 18340 13970 18352
rect 13964 18312 16620 18340
rect 13964 18300 13970 18312
rect 12986 18272 12992 18284
rect 12947 18244 12992 18272
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 13630 18232 13636 18284
rect 13688 18272 13694 18284
rect 14001 18275 14059 18281
rect 14001 18272 14013 18275
rect 13688 18244 14013 18272
rect 13688 18232 13694 18244
rect 14001 18241 14013 18244
rect 14047 18241 14059 18275
rect 14001 18235 14059 18241
rect 15470 18232 15476 18284
rect 15528 18272 15534 18284
rect 15565 18275 15623 18281
rect 15565 18272 15577 18275
rect 15528 18244 15577 18272
rect 15528 18232 15534 18244
rect 15565 18241 15577 18244
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18272 15807 18275
rect 15930 18272 15936 18284
rect 15795 18244 15936 18272
rect 15795 18241 15807 18244
rect 15749 18235 15807 18241
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 16592 18281 16620 18312
rect 16577 18275 16635 18281
rect 16577 18241 16589 18275
rect 16623 18241 16635 18275
rect 16758 18272 16764 18284
rect 16719 18244 16764 18272
rect 16577 18235 16635 18241
rect 16758 18232 16764 18244
rect 16816 18232 16822 18284
rect 11002 18176 12388 18204
rect 11002 18173 11014 18176
rect 10956 18167 11014 18173
rect 12710 18164 12716 18216
rect 12768 18204 12774 18216
rect 12805 18207 12863 18213
rect 12805 18204 12817 18207
rect 12768 18176 12817 18204
rect 12768 18164 12774 18176
rect 12805 18173 12817 18176
rect 12851 18173 12863 18207
rect 13814 18204 13820 18216
rect 13775 18176 13820 18204
rect 12805 18167 12863 18173
rect 13814 18164 13820 18176
rect 13872 18164 13878 18216
rect 14553 18207 14611 18213
rect 14553 18173 14565 18207
rect 14599 18204 14611 18207
rect 17328 18204 17356 18380
rect 18690 18368 18696 18380
rect 18748 18368 18754 18420
rect 17589 18343 17647 18349
rect 17589 18309 17601 18343
rect 17635 18340 17647 18343
rect 18506 18340 18512 18352
rect 17635 18312 18512 18340
rect 17635 18309 17647 18312
rect 17589 18303 17647 18309
rect 18506 18300 18512 18312
rect 18564 18300 18570 18352
rect 19521 18275 19579 18281
rect 19521 18272 19533 18275
rect 17420 18244 19533 18272
rect 17420 18213 17448 18244
rect 19521 18241 19533 18244
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 20717 18275 20775 18281
rect 20717 18241 20729 18275
rect 20763 18272 20775 18275
rect 20898 18272 20904 18284
rect 20763 18244 20904 18272
rect 20763 18241 20775 18244
rect 20717 18235 20775 18241
rect 20898 18232 20904 18244
rect 20956 18232 20962 18284
rect 14599 18176 17356 18204
rect 17405 18207 17463 18213
rect 14599 18173 14611 18176
rect 14553 18167 14611 18173
rect 17405 18173 17417 18207
rect 17451 18173 17463 18207
rect 17405 18167 17463 18173
rect 18414 18164 18420 18216
rect 18472 18204 18478 18216
rect 18509 18207 18567 18213
rect 18509 18204 18521 18207
rect 18472 18176 18521 18204
rect 18472 18164 18478 18176
rect 18509 18173 18521 18176
rect 18555 18173 18567 18207
rect 18509 18167 18567 18173
rect 18598 18164 18604 18216
rect 18656 18204 18662 18216
rect 18785 18207 18843 18213
rect 18785 18204 18797 18207
rect 18656 18176 18797 18204
rect 18656 18164 18662 18176
rect 18785 18173 18797 18176
rect 18831 18173 18843 18207
rect 19334 18204 19340 18216
rect 19295 18176 19340 18204
rect 18785 18167 18843 18173
rect 19334 18164 19340 18176
rect 19392 18164 19398 18216
rect 19610 18164 19616 18216
rect 19668 18204 19674 18216
rect 20441 18207 20499 18213
rect 20441 18204 20453 18207
rect 19668 18176 20453 18204
rect 19668 18164 19674 18176
rect 20441 18173 20453 18176
rect 20487 18173 20499 18207
rect 20441 18167 20499 18173
rect 4908 18108 6316 18136
rect 7837 18139 7895 18145
rect 7837 18105 7849 18139
rect 7883 18136 7895 18139
rect 8570 18136 8576 18148
rect 7883 18108 8576 18136
rect 7883 18105 7895 18108
rect 7837 18099 7895 18105
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 8849 18139 8907 18145
rect 8849 18105 8861 18139
rect 8895 18136 8907 18139
rect 9674 18136 9680 18148
rect 8895 18108 9680 18136
rect 8895 18105 8907 18108
rect 8849 18099 8907 18105
rect 9674 18096 9680 18108
rect 9732 18096 9738 18148
rect 10134 18096 10140 18148
rect 10192 18136 10198 18148
rect 11238 18136 11244 18148
rect 10192 18108 11244 18136
rect 10192 18096 10198 18108
rect 11238 18096 11244 18108
rect 11296 18096 11302 18148
rect 11790 18096 11796 18148
rect 11848 18136 11854 18148
rect 12897 18139 12955 18145
rect 12897 18136 12909 18139
rect 11848 18108 12909 18136
rect 11848 18096 11854 18108
rect 12897 18105 12909 18108
rect 12943 18105 12955 18139
rect 12897 18099 12955 18105
rect 13170 18096 13176 18148
rect 13228 18136 13234 18148
rect 13909 18139 13967 18145
rect 13909 18136 13921 18139
rect 13228 18108 13921 18136
rect 13228 18096 13234 18108
rect 13909 18105 13921 18108
rect 13955 18105 13967 18139
rect 15473 18139 15531 18145
rect 13909 18099 13967 18105
rect 14200 18108 15424 18136
rect 3789 18071 3847 18077
rect 3789 18037 3801 18071
rect 3835 18037 3847 18071
rect 3789 18031 3847 18037
rect 4065 18071 4123 18077
rect 4065 18037 4077 18071
rect 4111 18068 4123 18071
rect 4338 18068 4344 18080
rect 4111 18040 4344 18068
rect 4111 18037 4123 18040
rect 4065 18031 4123 18037
rect 4338 18028 4344 18040
rect 4396 18028 4402 18080
rect 4430 18028 4436 18080
rect 4488 18068 4494 18080
rect 4985 18071 5043 18077
rect 4488 18040 4533 18068
rect 4488 18028 4494 18040
rect 4985 18037 4997 18071
rect 5031 18068 5043 18071
rect 5350 18068 5356 18080
rect 5031 18040 5356 18068
rect 5031 18037 5043 18040
rect 4985 18031 5043 18037
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 6454 18068 6460 18080
rect 6415 18040 6460 18068
rect 6454 18028 6460 18040
rect 6512 18028 6518 18080
rect 7929 18071 7987 18077
rect 7929 18037 7941 18071
rect 7975 18068 7987 18071
rect 9766 18068 9772 18080
rect 7975 18040 9772 18068
rect 7975 18037 7987 18040
rect 7929 18031 7987 18037
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 9953 18071 10011 18077
rect 9953 18037 9965 18071
rect 9999 18068 10011 18071
rect 10042 18068 10048 18080
rect 9999 18040 10048 18068
rect 9999 18037 10011 18040
rect 9953 18031 10011 18037
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 12526 18028 12532 18080
rect 12584 18068 12590 18080
rect 14200 18068 14228 18108
rect 12584 18040 14228 18068
rect 12584 18028 12590 18040
rect 14366 18028 14372 18080
rect 14424 18068 14430 18080
rect 14737 18071 14795 18077
rect 14737 18068 14749 18071
rect 14424 18040 14749 18068
rect 14424 18028 14430 18040
rect 14737 18037 14749 18040
rect 14783 18037 14795 18071
rect 15396 18068 15424 18108
rect 15473 18105 15485 18139
rect 15519 18136 15531 18139
rect 16298 18136 16304 18148
rect 15519 18108 16304 18136
rect 15519 18105 15531 18108
rect 15473 18099 15531 18105
rect 16298 18096 16304 18108
rect 16356 18096 16362 18148
rect 19702 18136 19708 18148
rect 16408 18108 19708 18136
rect 16408 18068 16436 18108
rect 19702 18096 19708 18108
rect 19760 18096 19766 18148
rect 19794 18096 19800 18148
rect 19852 18136 19858 18148
rect 20533 18139 20591 18145
rect 20533 18136 20545 18139
rect 19852 18108 20545 18136
rect 19852 18096 19858 18108
rect 20533 18105 20545 18108
rect 20579 18105 20591 18139
rect 20533 18099 20591 18105
rect 15396 18040 16436 18068
rect 16485 18071 16543 18077
rect 14737 18031 14795 18037
rect 16485 18037 16497 18071
rect 16531 18068 16543 18071
rect 16942 18068 16948 18080
rect 16531 18040 16948 18068
rect 16531 18037 16543 18040
rect 16485 18031 16543 18037
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 18414 18068 18420 18080
rect 18375 18040 18420 18068
rect 18414 18028 18420 18040
rect 18472 18028 18478 18080
rect 20070 18068 20076 18080
rect 20031 18040 20076 18068
rect 20070 18028 20076 18040
rect 20128 18028 20134 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 198 17824 204 17876
rect 256 17864 262 17876
rect 1854 17864 1860 17876
rect 256 17836 1860 17864
rect 256 17824 262 17836
rect 1854 17824 1860 17836
rect 1912 17824 1918 17876
rect 2409 17867 2467 17873
rect 2409 17833 2421 17867
rect 2455 17833 2467 17867
rect 2866 17864 2872 17876
rect 2827 17836 2872 17864
rect 2409 17827 2467 17833
rect 2424 17796 2452 17827
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 3234 17864 3240 17876
rect 3108 17836 3240 17864
rect 3108 17824 3114 17836
rect 3234 17824 3240 17836
rect 3292 17824 3298 17876
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 3476 17836 4077 17864
rect 3476 17824 3482 17836
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 4338 17824 4344 17876
rect 4396 17864 4402 17876
rect 4525 17867 4583 17873
rect 4525 17864 4537 17867
rect 4396 17836 4537 17864
rect 4396 17824 4402 17836
rect 4525 17833 4537 17836
rect 4571 17833 4583 17867
rect 5074 17864 5080 17876
rect 5035 17836 5080 17864
rect 4525 17827 4583 17833
rect 5074 17824 5080 17836
rect 5132 17824 5138 17876
rect 6822 17864 6828 17876
rect 6783 17836 6828 17864
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7098 17864 7104 17876
rect 6972 17836 7104 17864
rect 6972 17824 6978 17836
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 7469 17867 7527 17873
rect 7469 17864 7481 17867
rect 7432 17836 7481 17864
rect 7432 17824 7438 17836
rect 7469 17833 7481 17836
rect 7515 17833 7527 17867
rect 8570 17864 8576 17876
rect 8531 17836 8576 17864
rect 7469 17827 7527 17833
rect 8570 17824 8576 17836
rect 8628 17824 8634 17876
rect 8941 17867 8999 17873
rect 8941 17833 8953 17867
rect 8987 17864 8999 17867
rect 9122 17864 9128 17876
rect 8987 17836 9128 17864
rect 8987 17833 8999 17836
rect 8941 17827 8999 17833
rect 9122 17824 9128 17836
rect 9180 17824 9186 17876
rect 9674 17864 9680 17876
rect 9635 17836 9680 17864
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 10042 17824 10048 17876
rect 10100 17864 10106 17876
rect 11057 17867 11115 17873
rect 11057 17864 11069 17867
rect 10100 17836 11069 17864
rect 10100 17824 10106 17836
rect 11057 17833 11069 17836
rect 11103 17833 11115 17867
rect 13078 17864 13084 17876
rect 11057 17827 11115 17833
rect 11808 17836 12388 17864
rect 13039 17836 13084 17864
rect 4433 17799 4491 17805
rect 4433 17796 4445 17799
rect 2424 17768 4445 17796
rect 4433 17765 4445 17768
rect 4479 17765 4491 17799
rect 7929 17799 7987 17805
rect 7929 17796 7941 17799
rect 4433 17759 4491 17765
rect 5184 17768 5672 17796
rect 934 17688 940 17740
rect 992 17728 998 17740
rect 1762 17728 1768 17740
rect 992 17700 1768 17728
rect 992 17688 998 17700
rect 1762 17688 1768 17700
rect 1820 17688 1826 17740
rect 2590 17688 2596 17740
rect 2648 17728 2654 17740
rect 2777 17731 2835 17737
rect 2777 17728 2789 17731
rect 2648 17700 2789 17728
rect 2648 17688 2654 17700
rect 2777 17697 2789 17700
rect 2823 17697 2835 17731
rect 3418 17728 3424 17740
rect 3379 17700 3424 17728
rect 2777 17691 2835 17697
rect 3418 17688 3424 17700
rect 3476 17688 3482 17740
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17660 2099 17663
rect 2498 17660 2504 17672
rect 2087 17632 2504 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 2498 17620 2504 17632
rect 2556 17620 2562 17672
rect 2958 17660 2964 17672
rect 2919 17632 2964 17660
rect 2958 17620 2964 17632
rect 3016 17620 3022 17672
rect 4522 17620 4528 17672
rect 4580 17660 4586 17672
rect 4709 17663 4767 17669
rect 4709 17660 4721 17663
rect 4580 17632 4721 17660
rect 4580 17620 4586 17632
rect 4709 17629 4721 17632
rect 4755 17660 4767 17663
rect 5184 17660 5212 17768
rect 5442 17728 5448 17740
rect 5403 17700 5448 17728
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 5534 17660 5540 17672
rect 4755 17632 5212 17660
rect 5495 17632 5540 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 5534 17620 5540 17632
rect 5592 17620 5598 17672
rect 5644 17669 5672 17768
rect 7024 17768 7941 17796
rect 6822 17688 6828 17740
rect 6880 17728 6886 17740
rect 7024 17728 7052 17768
rect 7929 17765 7941 17768
rect 7975 17765 7987 17799
rect 11808 17796 11836 17836
rect 7929 17759 7987 17765
rect 8036 17768 11836 17796
rect 6880 17700 7052 17728
rect 6880 17688 6886 17700
rect 7190 17688 7196 17740
rect 7248 17728 7254 17740
rect 7837 17731 7895 17737
rect 7837 17728 7849 17731
rect 7248 17700 7849 17728
rect 7248 17688 7254 17700
rect 7837 17697 7849 17700
rect 7883 17697 7895 17731
rect 7837 17691 7895 17697
rect 5629 17663 5687 17669
rect 5629 17629 5641 17663
rect 5675 17629 5687 17663
rect 6917 17663 6975 17669
rect 6917 17660 6929 17663
rect 5629 17623 5687 17629
rect 5736 17632 6929 17660
rect 1397 17595 1455 17601
rect 1397 17561 1409 17595
rect 1443 17592 1455 17595
rect 5736 17592 5764 17632
rect 6917 17629 6929 17632
rect 6963 17629 6975 17663
rect 7098 17660 7104 17672
rect 7059 17632 7104 17660
rect 6917 17623 6975 17629
rect 7098 17620 7104 17632
rect 7156 17620 7162 17672
rect 1443 17564 5764 17592
rect 1443 17561 1455 17564
rect 1397 17555 1455 17561
rect 6086 17552 6092 17604
rect 6144 17592 6150 17604
rect 8036 17592 8064 17768
rect 11882 17756 11888 17808
rect 11940 17796 11946 17808
rect 12360 17796 12388 17836
rect 13078 17824 13084 17836
rect 13136 17824 13142 17876
rect 15930 17824 15936 17876
rect 15988 17824 15994 17876
rect 16666 17824 16672 17876
rect 16724 17864 16730 17876
rect 17405 17867 17463 17873
rect 17405 17864 17417 17867
rect 16724 17836 17417 17864
rect 16724 17824 16730 17836
rect 17405 17833 17417 17836
rect 17451 17833 17463 17867
rect 17405 17827 17463 17833
rect 17494 17824 17500 17876
rect 17552 17864 17558 17876
rect 17865 17867 17923 17873
rect 17865 17864 17877 17867
rect 17552 17836 17877 17864
rect 17552 17824 17558 17836
rect 17865 17833 17877 17836
rect 17911 17833 17923 17867
rect 17865 17827 17923 17833
rect 19245 17867 19303 17873
rect 19245 17833 19257 17867
rect 19291 17864 19303 17867
rect 19797 17867 19855 17873
rect 19797 17864 19809 17867
rect 19291 17836 19809 17864
rect 19291 17833 19303 17836
rect 19245 17827 19303 17833
rect 19797 17833 19809 17836
rect 19843 17833 19855 17867
rect 21450 17864 21456 17876
rect 19797 17827 19855 17833
rect 20088 17836 21456 17864
rect 13909 17799 13967 17805
rect 13909 17796 13921 17799
rect 11940 17768 12296 17796
rect 12360 17768 13921 17796
rect 11940 17756 11946 17768
rect 8386 17688 8392 17740
rect 8444 17728 8450 17740
rect 8662 17728 8668 17740
rect 8444 17700 8668 17728
rect 8444 17688 8450 17700
rect 8662 17688 8668 17700
rect 8720 17688 8726 17740
rect 8754 17688 8760 17740
rect 8812 17728 8818 17740
rect 8812 17700 9168 17728
rect 8812 17688 8818 17700
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17660 8171 17663
rect 8294 17660 8300 17672
rect 8159 17632 8300 17660
rect 8159 17629 8171 17632
rect 8113 17623 8171 17629
rect 8294 17620 8300 17632
rect 8352 17620 8358 17672
rect 9030 17660 9036 17672
rect 8991 17632 9036 17660
rect 9030 17620 9036 17632
rect 9088 17620 9094 17672
rect 9140 17669 9168 17700
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9456 17700 10057 17728
rect 9456 17688 9462 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10962 17728 10968 17740
rect 10045 17691 10103 17697
rect 10244 17700 10968 17728
rect 9125 17663 9183 17669
rect 9125 17629 9137 17663
rect 9171 17629 9183 17663
rect 10134 17660 10140 17672
rect 10095 17632 10140 17660
rect 9125 17623 9183 17629
rect 6144 17564 8064 17592
rect 9140 17592 9168 17623
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 10244 17669 10272 17700
rect 10962 17688 10968 17700
rect 11020 17688 11026 17740
rect 11149 17731 11207 17737
rect 11149 17697 11161 17731
rect 11195 17728 11207 17731
rect 11238 17728 11244 17740
rect 11195 17700 11244 17728
rect 11195 17697 11207 17700
rect 11149 17691 11207 17697
rect 11238 17688 11244 17700
rect 11296 17688 11302 17740
rect 12066 17688 12072 17740
rect 12124 17728 12130 17740
rect 12161 17731 12219 17737
rect 12161 17728 12173 17731
rect 12124 17700 12173 17728
rect 12124 17688 12130 17700
rect 12161 17697 12173 17700
rect 12207 17697 12219 17731
rect 12268 17728 12296 17768
rect 13909 17765 13921 17768
rect 13955 17765 13967 17799
rect 13909 17759 13967 17765
rect 12268 17700 12388 17728
rect 12161 17691 12219 17697
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17629 10287 17663
rect 10229 17623 10287 17629
rect 11333 17663 11391 17669
rect 11333 17629 11345 17663
rect 11379 17660 11391 17663
rect 11882 17660 11888 17672
rect 11379 17632 11888 17660
rect 11379 17629 11391 17632
rect 11333 17623 11391 17629
rect 10244 17592 10272 17623
rect 11882 17620 11888 17632
rect 11940 17620 11946 17672
rect 12250 17660 12256 17672
rect 12211 17632 12256 17660
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 12360 17669 12388 17700
rect 12526 17688 12532 17740
rect 12584 17728 12590 17740
rect 12897 17731 12955 17737
rect 12897 17728 12909 17731
rect 12584 17700 12909 17728
rect 12584 17688 12590 17700
rect 12897 17697 12909 17700
rect 12943 17697 12955 17731
rect 12897 17691 12955 17697
rect 13078 17688 13084 17740
rect 13136 17728 13142 17740
rect 13817 17731 13875 17737
rect 13817 17728 13829 17731
rect 13136 17700 13829 17728
rect 13136 17688 13142 17700
rect 13817 17697 13829 17700
rect 13863 17697 13875 17731
rect 13817 17691 13875 17697
rect 14461 17731 14519 17737
rect 14461 17697 14473 17731
rect 14507 17728 14519 17731
rect 14642 17728 14648 17740
rect 14507 17700 14648 17728
rect 14507 17697 14519 17700
rect 14461 17691 14519 17697
rect 14642 17688 14648 17700
rect 14700 17688 14706 17740
rect 15194 17688 15200 17740
rect 15252 17728 15258 17740
rect 15948 17728 15976 17824
rect 17773 17799 17831 17805
rect 17773 17765 17785 17799
rect 17819 17796 17831 17799
rect 20088 17796 20116 17836
rect 21450 17824 21456 17836
rect 21508 17824 21514 17876
rect 17819 17768 20116 17796
rect 20165 17799 20223 17805
rect 17819 17765 17831 17768
rect 17773 17759 17831 17765
rect 20165 17765 20177 17799
rect 20211 17796 20223 17799
rect 20254 17796 20260 17808
rect 20211 17768 20260 17796
rect 20211 17765 20223 17768
rect 20165 17759 20223 17765
rect 20254 17756 20260 17768
rect 20312 17756 20318 17808
rect 16005 17731 16063 17737
rect 16005 17728 16017 17731
rect 15252 17700 16017 17728
rect 15252 17688 15258 17700
rect 16005 17697 16017 17700
rect 16051 17728 16063 17731
rect 16574 17728 16580 17740
rect 16051 17700 16580 17728
rect 16051 17697 16063 17700
rect 16005 17691 16063 17697
rect 16574 17688 16580 17700
rect 16632 17688 16638 17740
rect 19150 17728 19156 17740
rect 19111 17700 19156 17728
rect 19150 17688 19156 17700
rect 19208 17688 19214 17740
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17629 12403 17663
rect 14090 17660 14096 17672
rect 14051 17632 14096 17660
rect 12345 17623 12403 17629
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17660 15347 17663
rect 15470 17660 15476 17672
rect 15335 17632 15476 17660
rect 15335 17629 15347 17632
rect 15289 17623 15347 17629
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 15749 17663 15807 17669
rect 15749 17629 15761 17663
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 17957 17663 18015 17669
rect 17957 17629 17969 17663
rect 18003 17629 18015 17663
rect 17957 17623 18015 17629
rect 14645 17595 14703 17601
rect 14645 17592 14657 17595
rect 9140 17564 10272 17592
rect 10336 17564 14657 17592
rect 6144 17552 6150 17564
rect 3142 17484 3148 17536
rect 3200 17524 3206 17536
rect 3605 17527 3663 17533
rect 3605 17524 3617 17527
rect 3200 17496 3617 17524
rect 3200 17484 3206 17496
rect 3605 17493 3617 17496
rect 3651 17493 3663 17527
rect 3605 17487 3663 17493
rect 6457 17527 6515 17533
rect 6457 17493 6469 17527
rect 6503 17524 6515 17527
rect 7098 17524 7104 17536
rect 6503 17496 7104 17524
rect 6503 17493 6515 17496
rect 6457 17487 6515 17493
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 7834 17484 7840 17536
rect 7892 17524 7898 17536
rect 10336 17524 10364 17564
rect 14645 17561 14657 17564
rect 14691 17561 14703 17595
rect 14645 17555 14703 17561
rect 7892 17496 10364 17524
rect 10689 17527 10747 17533
rect 7892 17484 7898 17496
rect 10689 17493 10701 17527
rect 10735 17524 10747 17527
rect 11606 17524 11612 17536
rect 10735 17496 11612 17524
rect 10735 17493 10747 17496
rect 10689 17487 10747 17493
rect 11606 17484 11612 17496
rect 11664 17484 11670 17536
rect 11793 17527 11851 17533
rect 11793 17493 11805 17527
rect 11839 17524 11851 17527
rect 13170 17524 13176 17536
rect 11839 17496 13176 17524
rect 11839 17493 11851 17496
rect 11793 17487 11851 17493
rect 13170 17484 13176 17496
rect 13228 17484 13234 17536
rect 13449 17527 13507 17533
rect 13449 17493 13461 17527
rect 13495 17524 13507 17527
rect 15654 17524 15660 17536
rect 13495 17496 15660 17524
rect 13495 17493 13507 17496
rect 13449 17487 13507 17493
rect 15654 17484 15660 17496
rect 15712 17484 15718 17536
rect 15764 17524 15792 17623
rect 16758 17552 16764 17604
rect 16816 17592 16822 17604
rect 17402 17592 17408 17604
rect 16816 17564 17408 17592
rect 16816 17552 16822 17564
rect 17402 17552 17408 17564
rect 17460 17592 17466 17604
rect 17972 17592 18000 17623
rect 19242 17620 19248 17672
rect 19300 17660 19306 17672
rect 19337 17663 19395 17669
rect 19337 17660 19349 17663
rect 19300 17632 19349 17660
rect 19300 17620 19306 17632
rect 19337 17629 19349 17632
rect 19383 17629 19395 17663
rect 19337 17623 19395 17629
rect 19886 17620 19892 17672
rect 19944 17660 19950 17672
rect 20257 17663 20315 17669
rect 20257 17660 20269 17663
rect 19944 17632 20269 17660
rect 19944 17620 19950 17632
rect 20257 17629 20269 17632
rect 20303 17629 20315 17663
rect 20438 17660 20444 17672
rect 20351 17632 20444 17660
rect 20257 17623 20315 17629
rect 20438 17620 20444 17632
rect 20496 17660 20502 17672
rect 20898 17660 20904 17672
rect 20496 17632 20904 17660
rect 20496 17620 20502 17632
rect 20898 17620 20904 17632
rect 20956 17620 20962 17672
rect 17460 17564 18000 17592
rect 17460 17552 17466 17564
rect 18598 17552 18604 17604
rect 18656 17592 18662 17604
rect 21726 17592 21732 17604
rect 18656 17564 21732 17592
rect 18656 17552 18662 17564
rect 21726 17552 21732 17564
rect 21784 17552 21790 17604
rect 15930 17524 15936 17536
rect 15764 17496 15936 17524
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 16482 17484 16488 17536
rect 16540 17524 16546 17536
rect 17129 17527 17187 17533
rect 17129 17524 17141 17527
rect 16540 17496 17141 17524
rect 16540 17484 16546 17496
rect 17129 17493 17141 17496
rect 17175 17493 17187 17527
rect 17129 17487 17187 17493
rect 18785 17527 18843 17533
rect 18785 17493 18797 17527
rect 18831 17524 18843 17527
rect 18874 17524 18880 17536
rect 18831 17496 18880 17524
rect 18831 17493 18843 17496
rect 18785 17487 18843 17493
rect 18874 17484 18880 17496
rect 18932 17484 18938 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 2038 17280 2044 17332
rect 2096 17320 2102 17332
rect 2774 17320 2780 17332
rect 2096 17292 2780 17320
rect 2096 17280 2102 17292
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 3513 17323 3571 17329
rect 3513 17320 3525 17323
rect 3108 17292 3525 17320
rect 3108 17280 3114 17292
rect 3513 17289 3525 17292
rect 3559 17289 3571 17323
rect 3513 17283 3571 17289
rect 4249 17323 4307 17329
rect 4249 17289 4261 17323
rect 4295 17320 4307 17323
rect 5534 17320 5540 17332
rect 4295 17292 5540 17320
rect 4295 17289 4307 17292
rect 4249 17283 4307 17289
rect 3528 17184 3556 17283
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 5629 17323 5687 17329
rect 5629 17289 5641 17323
rect 5675 17320 5687 17323
rect 7834 17320 7840 17332
rect 5675 17292 7840 17320
rect 5675 17289 5687 17292
rect 5629 17283 5687 17289
rect 7834 17280 7840 17292
rect 7892 17280 7898 17332
rect 8294 17320 8300 17332
rect 8255 17292 8300 17320
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 9398 17320 9404 17332
rect 9359 17292 9404 17320
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 10413 17323 10471 17329
rect 10413 17320 10425 17323
rect 9824 17292 10425 17320
rect 9824 17280 9830 17292
rect 10413 17289 10425 17292
rect 10459 17289 10471 17323
rect 10413 17283 10471 17289
rect 11609 17323 11667 17329
rect 11609 17289 11621 17323
rect 11655 17320 11667 17323
rect 12342 17320 12348 17332
rect 11655 17292 12348 17320
rect 11655 17289 11667 17292
rect 11609 17283 11667 17289
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12492 17292 12537 17320
rect 12492 17280 12498 17292
rect 13722 17280 13728 17332
rect 13780 17320 13786 17332
rect 13780 17292 16427 17320
rect 13780 17280 13786 17292
rect 9033 17255 9091 17261
rect 9033 17221 9045 17255
rect 9079 17252 9091 17255
rect 10778 17252 10784 17264
rect 9079 17224 10784 17252
rect 9079 17221 9091 17224
rect 9033 17215 9091 17221
rect 10778 17212 10784 17224
rect 10836 17212 10842 17264
rect 12250 17252 12256 17264
rect 11072 17224 12256 17252
rect 4246 17184 4252 17196
rect 1412 17156 2268 17184
rect 3528 17156 4252 17184
rect 1412 17125 1440 17156
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17085 1455 17119
rect 1397 17079 1455 17085
rect 2133 17119 2191 17125
rect 2133 17085 2145 17119
rect 2179 17085 2191 17119
rect 2240 17116 2268 17156
rect 4246 17144 4252 17156
rect 4304 17184 4310 17196
rect 4706 17184 4712 17196
rect 4304 17156 4712 17184
rect 4304 17144 4310 17156
rect 4706 17144 4712 17156
rect 4764 17184 4770 17196
rect 4801 17187 4859 17193
rect 4801 17184 4813 17187
rect 4764 17156 4813 17184
rect 4764 17144 4770 17156
rect 4801 17153 4813 17156
rect 4847 17153 4859 17187
rect 4801 17147 4859 17153
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 6181 17187 6239 17193
rect 6181 17184 6193 17187
rect 5316 17156 6193 17184
rect 5316 17144 5322 17156
rect 6181 17153 6193 17156
rect 6227 17153 6239 17187
rect 6181 17147 6239 17153
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17184 6423 17187
rect 6454 17184 6460 17196
rect 6411 17156 6460 17184
rect 6411 17153 6423 17156
rect 6365 17147 6423 17153
rect 6454 17144 6460 17156
rect 6512 17144 6518 17196
rect 6638 17144 6644 17196
rect 6696 17184 6702 17196
rect 6917 17187 6975 17193
rect 6917 17184 6929 17187
rect 6696 17156 6929 17184
rect 6696 17144 6702 17156
rect 6917 17153 6929 17156
rect 6963 17153 6975 17187
rect 6917 17147 6975 17153
rect 2866 17116 2872 17128
rect 2240 17088 2872 17116
rect 2133 17079 2191 17085
rect 1670 17048 1676 17060
rect 1631 17020 1676 17048
rect 1670 17008 1676 17020
rect 1728 17008 1734 17060
rect 2148 17048 2176 17079
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 3878 17076 3884 17128
rect 3936 17116 3942 17128
rect 3936 17088 4752 17116
rect 3936 17076 3942 17088
rect 2222 17048 2228 17060
rect 2148 17020 2228 17048
rect 2222 17008 2228 17020
rect 2280 17008 2286 17060
rect 2406 17057 2412 17060
rect 2400 17048 2412 17057
rect 2367 17020 2412 17048
rect 2400 17011 2412 17020
rect 2406 17008 2412 17011
rect 2464 17008 2470 17060
rect 4617 17051 4675 17057
rect 4617 17048 4629 17051
rect 2516 17020 4629 17048
rect 1762 16940 1768 16992
rect 1820 16980 1826 16992
rect 2516 16980 2544 17020
rect 4617 17017 4629 17020
rect 4663 17017 4675 17051
rect 4724 17048 4752 17088
rect 4890 17076 4896 17128
rect 4948 17116 4954 17128
rect 6089 17119 6147 17125
rect 6089 17116 6101 17119
rect 4948 17088 6101 17116
rect 4948 17076 4954 17088
rect 6089 17085 6101 17088
rect 6135 17085 6147 17119
rect 6932 17116 6960 17147
rect 8018 17144 8024 17196
rect 8076 17184 8082 17196
rect 8076 17156 8984 17184
rect 8076 17144 8082 17156
rect 7650 17116 7656 17128
rect 6932 17088 7656 17116
rect 6089 17079 6147 17085
rect 7650 17076 7656 17088
rect 7708 17076 7714 17128
rect 8846 17116 8852 17128
rect 8807 17088 8852 17116
rect 8846 17076 8852 17088
rect 8904 17076 8910 17128
rect 8956 17116 8984 17156
rect 9582 17144 9588 17196
rect 9640 17184 9646 17196
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 9640 17156 9965 17184
rect 9640 17144 9646 17156
rect 9953 17153 9965 17156
rect 9999 17153 10011 17187
rect 10962 17184 10968 17196
rect 10923 17156 10968 17184
rect 9953 17147 10011 17153
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 11072 17116 11100 17224
rect 12250 17212 12256 17224
rect 12308 17252 12314 17264
rect 13446 17252 13452 17264
rect 12308 17224 13452 17252
rect 12308 17212 12314 17224
rect 13446 17212 13452 17224
rect 13504 17212 13510 17264
rect 15197 17255 15255 17261
rect 15197 17221 15209 17255
rect 15243 17221 15255 17255
rect 16399 17252 16427 17292
rect 16574 17280 16580 17332
rect 16632 17320 16638 17332
rect 16853 17323 16911 17329
rect 16853 17320 16865 17323
rect 16632 17292 16865 17320
rect 16632 17280 16638 17292
rect 16853 17289 16865 17292
rect 16899 17289 16911 17323
rect 19058 17320 19064 17332
rect 19019 17292 19064 17320
rect 16853 17283 16911 17289
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 19150 17280 19156 17332
rect 19208 17320 19214 17332
rect 20257 17323 20315 17329
rect 20257 17320 20269 17323
rect 19208 17292 20269 17320
rect 19208 17280 19214 17292
rect 20257 17289 20269 17292
rect 20303 17289 20315 17323
rect 20257 17283 20315 17289
rect 16666 17252 16672 17264
rect 16399 17224 16672 17252
rect 15197 17215 15255 17221
rect 11606 17144 11612 17196
rect 11664 17184 11670 17196
rect 12897 17187 12955 17193
rect 12897 17184 12909 17187
rect 11664 17156 12909 17184
rect 11664 17144 11670 17156
rect 12897 17153 12909 17156
rect 12943 17153 12955 17187
rect 12897 17147 12955 17153
rect 12986 17144 12992 17196
rect 13044 17184 13050 17196
rect 13081 17187 13139 17193
rect 13081 17184 13093 17187
rect 13044 17156 13093 17184
rect 13044 17144 13050 17156
rect 13081 17153 13093 17156
rect 13127 17184 13139 17187
rect 13630 17184 13636 17196
rect 13127 17156 13636 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 15212 17184 15240 17215
rect 16666 17212 16672 17224
rect 16724 17212 16730 17264
rect 18049 17255 18107 17261
rect 18049 17221 18061 17255
rect 18095 17252 18107 17255
rect 19334 17252 19340 17264
rect 18095 17224 19340 17252
rect 18095 17221 18107 17224
rect 18049 17215 18107 17221
rect 19334 17212 19340 17224
rect 19392 17212 19398 17264
rect 19518 17212 19524 17264
rect 19576 17252 19582 17264
rect 19702 17252 19708 17264
rect 19576 17224 19708 17252
rect 19576 17212 19582 17224
rect 19702 17212 19708 17224
rect 19760 17212 19766 17264
rect 18693 17187 18751 17193
rect 15212 17156 15424 17184
rect 8956 17088 11100 17116
rect 11146 17076 11152 17128
rect 11204 17116 11210 17128
rect 11425 17119 11483 17125
rect 11425 17116 11437 17119
rect 11204 17088 11437 17116
rect 11204 17076 11210 17088
rect 11425 17085 11437 17088
rect 11471 17085 11483 17119
rect 11425 17079 11483 17085
rect 11790 17076 11796 17128
rect 11848 17116 11854 17128
rect 12526 17116 12532 17128
rect 11848 17088 12532 17116
rect 11848 17076 11854 17088
rect 12526 17076 12532 17088
rect 12584 17076 12590 17128
rect 14090 17125 14096 17128
rect 13817 17119 13875 17125
rect 13817 17116 13829 17119
rect 12912 17088 13829 17116
rect 12912 17060 12940 17088
rect 13817 17085 13829 17088
rect 13863 17085 13875 17119
rect 14084 17116 14096 17125
rect 14003 17088 14096 17116
rect 13817 17079 13875 17085
rect 14084 17079 14096 17088
rect 14148 17116 14154 17128
rect 15286 17116 15292 17128
rect 14148 17088 15292 17116
rect 14090 17076 14096 17079
rect 14148 17076 14154 17088
rect 15286 17076 15292 17088
rect 15344 17076 15350 17128
rect 5537 17051 5595 17057
rect 5537 17048 5549 17051
rect 4724 17020 5549 17048
rect 4617 17011 4675 17017
rect 5537 17017 5549 17020
rect 5583 17017 5595 17051
rect 7184 17051 7242 17057
rect 5537 17011 5595 17017
rect 5736 17020 7144 17048
rect 1820 16952 2544 16980
rect 3789 16983 3847 16989
rect 1820 16940 1826 16952
rect 3789 16949 3801 16983
rect 3835 16980 3847 16983
rect 4430 16980 4436 16992
rect 3835 16952 4436 16980
rect 3835 16949 3847 16952
rect 3789 16943 3847 16949
rect 4430 16940 4436 16952
rect 4488 16940 4494 16992
rect 4706 16980 4712 16992
rect 4667 16952 4712 16980
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 5261 16983 5319 16989
rect 5261 16949 5273 16983
rect 5307 16980 5319 16983
rect 5626 16980 5632 16992
rect 5307 16952 5632 16980
rect 5307 16949 5319 16952
rect 5261 16943 5319 16949
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 5736 16989 5764 17020
rect 5721 16983 5779 16989
rect 5721 16949 5733 16983
rect 5767 16949 5779 16983
rect 7116 16980 7144 17020
rect 7184 17017 7196 17051
rect 7230 17048 7242 17051
rect 7466 17048 7472 17060
rect 7230 17020 7472 17048
rect 7230 17017 7242 17020
rect 7184 17011 7242 17017
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 8570 17008 8576 17060
rect 8628 17048 8634 17060
rect 9861 17051 9919 17057
rect 9861 17048 9873 17051
rect 8628 17020 9873 17048
rect 8628 17008 8634 17020
rect 9861 17017 9873 17020
rect 9907 17017 9919 17051
rect 9861 17011 9919 17017
rect 10781 17051 10839 17057
rect 10781 17017 10793 17051
rect 10827 17048 10839 17051
rect 12710 17048 12716 17060
rect 10827 17020 12716 17048
rect 10827 17017 10839 17020
rect 10781 17011 10839 17017
rect 12710 17008 12716 17020
rect 12768 17008 12774 17060
rect 12894 17008 12900 17060
rect 12952 17008 12958 17060
rect 13722 17008 13728 17060
rect 13780 17048 13786 17060
rect 14182 17048 14188 17060
rect 13780 17020 14188 17048
rect 13780 17008 13786 17020
rect 14182 17008 14188 17020
rect 14240 17008 14246 17060
rect 15396 17048 15424 17156
rect 18693 17153 18705 17187
rect 18739 17184 18751 17187
rect 18874 17184 18880 17196
rect 18739 17156 18880 17184
rect 18739 17153 18751 17156
rect 18693 17147 18751 17153
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 19613 17187 19671 17193
rect 19613 17153 19625 17187
rect 19659 17184 19671 17187
rect 20438 17184 20444 17196
rect 19659 17156 20444 17184
rect 19659 17153 19671 17156
rect 19613 17147 19671 17153
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 20898 17184 20904 17196
rect 20811 17156 20904 17184
rect 20898 17144 20904 17156
rect 20956 17184 20962 17196
rect 21821 17187 21879 17193
rect 21821 17184 21833 17187
rect 20956 17156 21833 17184
rect 20956 17144 20962 17156
rect 21821 17153 21833 17156
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 15473 17119 15531 17125
rect 15473 17085 15485 17119
rect 15519 17116 15531 17119
rect 15519 17088 16160 17116
rect 15519 17085 15531 17088
rect 15473 17079 15531 17085
rect 15718 17051 15776 17057
rect 15718 17048 15730 17051
rect 15396 17020 15730 17048
rect 15718 17017 15730 17020
rect 15764 17048 15776 17051
rect 16022 17048 16028 17060
rect 15764 17020 16028 17048
rect 15764 17017 15776 17020
rect 15718 17011 15776 17017
rect 16022 17008 16028 17020
rect 16080 17008 16086 17060
rect 9674 16980 9680 16992
rect 7116 16952 9680 16980
rect 5721 16943 5779 16949
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 9769 16983 9827 16989
rect 9769 16949 9781 16983
rect 9815 16980 9827 16983
rect 10042 16980 10048 16992
rect 9815 16952 10048 16980
rect 9815 16949 9827 16952
rect 9769 16943 9827 16949
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10502 16940 10508 16992
rect 10560 16980 10566 16992
rect 10873 16983 10931 16989
rect 10873 16980 10885 16983
rect 10560 16952 10885 16980
rect 10560 16940 10566 16952
rect 10873 16949 10885 16952
rect 10919 16949 10931 16983
rect 12802 16980 12808 16992
rect 12763 16952 12808 16980
rect 10873 16943 10931 16949
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 15930 16940 15936 16992
rect 15988 16980 15994 16992
rect 16132 16980 16160 17088
rect 16574 17076 16580 17128
rect 16632 17116 16638 17128
rect 17405 17119 17463 17125
rect 17405 17116 17417 17119
rect 16632 17088 17417 17116
rect 16632 17076 16638 17088
rect 17405 17085 17417 17088
rect 17451 17085 17463 17119
rect 17405 17079 17463 17085
rect 18509 17119 18567 17125
rect 18509 17085 18521 17119
rect 18555 17116 18567 17119
rect 19058 17116 19064 17128
rect 18555 17088 19064 17116
rect 18555 17085 18567 17088
rect 18509 17079 18567 17085
rect 19058 17076 19064 17088
rect 19116 17076 19122 17128
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 19521 17119 19579 17125
rect 19521 17116 19533 17119
rect 19392 17088 19533 17116
rect 19392 17076 19398 17088
rect 19521 17085 19533 17088
rect 19567 17085 19579 17119
rect 19521 17079 19579 17085
rect 20530 17076 20536 17128
rect 20588 17116 20594 17128
rect 20625 17119 20683 17125
rect 20625 17116 20637 17119
rect 20588 17088 20637 17116
rect 20588 17076 20594 17088
rect 20625 17085 20637 17088
rect 20671 17085 20683 17119
rect 20625 17079 20683 17085
rect 19150 17008 19156 17060
rect 19208 17048 19214 17060
rect 21634 17048 21640 17060
rect 19208 17020 21640 17048
rect 19208 17008 19214 17020
rect 21634 17008 21640 17020
rect 21692 17008 21698 17060
rect 15988 16952 16160 16980
rect 17589 16983 17647 16989
rect 15988 16940 15994 16952
rect 17589 16949 17601 16983
rect 17635 16980 17647 16983
rect 17954 16980 17960 16992
rect 17635 16952 17960 16980
rect 17635 16949 17647 16952
rect 17589 16943 17647 16949
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 18414 16980 18420 16992
rect 18375 16952 18420 16980
rect 18414 16940 18420 16952
rect 18472 16940 18478 16992
rect 19426 16980 19432 16992
rect 19387 16952 19432 16980
rect 19426 16940 19432 16952
rect 19484 16940 19490 16992
rect 20622 16940 20628 16992
rect 20680 16980 20686 16992
rect 20717 16983 20775 16989
rect 20717 16980 20729 16983
rect 20680 16952 20729 16980
rect 20680 16940 20686 16952
rect 20717 16949 20729 16952
rect 20763 16949 20775 16983
rect 20717 16943 20775 16949
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1581 16779 1639 16785
rect 1581 16745 1593 16779
rect 1627 16776 1639 16779
rect 1762 16776 1768 16788
rect 1627 16748 1768 16776
rect 1627 16745 1639 16748
rect 1581 16739 1639 16745
rect 1762 16736 1768 16748
rect 1820 16736 1826 16788
rect 2038 16776 2044 16788
rect 1999 16748 2044 16776
rect 2038 16736 2044 16748
rect 2096 16736 2102 16788
rect 2590 16776 2596 16788
rect 2551 16748 2596 16776
rect 2590 16736 2596 16748
rect 2648 16736 2654 16788
rect 4065 16779 4123 16785
rect 4065 16745 4077 16779
rect 4111 16745 4123 16779
rect 4430 16776 4436 16788
rect 4391 16748 4436 16776
rect 4065 16739 4123 16745
rect 1949 16711 2007 16717
rect 1949 16677 1961 16711
rect 1995 16708 2007 16711
rect 2774 16708 2780 16720
rect 1995 16680 2780 16708
rect 1995 16677 2007 16680
rect 1949 16671 2007 16677
rect 2774 16668 2780 16680
rect 2832 16668 2838 16720
rect 3234 16668 3240 16720
rect 3292 16668 3298 16720
rect 3970 16668 3976 16720
rect 4028 16708 4034 16720
rect 4080 16708 4108 16739
rect 4430 16736 4436 16748
rect 4488 16736 4494 16788
rect 4522 16736 4528 16788
rect 4580 16776 4586 16788
rect 4580 16748 6132 16776
rect 4580 16736 4586 16748
rect 4028 16680 4108 16708
rect 4028 16668 4034 16680
rect 4338 16668 4344 16720
rect 4396 16708 4402 16720
rect 5994 16708 6000 16720
rect 4396 16680 6000 16708
rect 4396 16668 4402 16680
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 6104 16708 6132 16748
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 6917 16779 6975 16785
rect 6917 16776 6929 16779
rect 6880 16748 6929 16776
rect 6880 16736 6886 16748
rect 6917 16745 6929 16748
rect 6963 16745 6975 16779
rect 6917 16739 6975 16745
rect 7098 16736 7104 16788
rect 7156 16776 7162 16788
rect 7377 16779 7435 16785
rect 7377 16776 7389 16779
rect 7156 16748 7389 16776
rect 7156 16736 7162 16748
rect 7377 16745 7389 16748
rect 7423 16745 7435 16779
rect 7377 16739 7435 16745
rect 9309 16779 9367 16785
rect 9309 16745 9321 16779
rect 9355 16776 9367 16779
rect 9582 16776 9588 16788
rect 9355 16748 9588 16776
rect 9355 16745 9367 16748
rect 9309 16739 9367 16745
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 10137 16779 10195 16785
rect 10137 16745 10149 16779
rect 10183 16776 10195 16779
rect 11054 16776 11060 16788
rect 10183 16748 11060 16776
rect 10183 16745 10195 16748
rect 10137 16739 10195 16745
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 11974 16736 11980 16788
rect 12032 16776 12038 16788
rect 12345 16779 12403 16785
rect 12345 16776 12357 16779
rect 12032 16748 12357 16776
rect 12032 16736 12038 16748
rect 12345 16745 12357 16748
rect 12391 16745 12403 16779
rect 12345 16739 12403 16745
rect 15289 16779 15347 16785
rect 15289 16745 15301 16779
rect 15335 16776 15347 16779
rect 15562 16776 15568 16788
rect 15335 16748 15568 16776
rect 15335 16745 15347 16748
rect 15289 16739 15347 16745
rect 15562 16736 15568 16748
rect 15620 16736 15626 16788
rect 15654 16736 15660 16788
rect 15712 16776 15718 16788
rect 15749 16779 15807 16785
rect 15749 16776 15761 16779
rect 15712 16748 15761 16776
rect 15712 16736 15718 16748
rect 15749 16745 15761 16748
rect 15795 16745 15807 16779
rect 16298 16776 16304 16788
rect 16259 16748 16304 16776
rect 15749 16739 15807 16745
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 16390 16736 16396 16788
rect 16448 16776 16454 16788
rect 17313 16779 17371 16785
rect 17313 16776 17325 16779
rect 16448 16748 17325 16776
rect 16448 16736 16454 16748
rect 17313 16745 17325 16748
rect 17359 16745 17371 16779
rect 18322 16776 18328 16788
rect 18283 16748 18328 16776
rect 17313 16739 17371 16745
rect 18322 16736 18328 16748
rect 18380 16736 18386 16788
rect 19429 16779 19487 16785
rect 19429 16745 19441 16779
rect 19475 16776 19487 16779
rect 19610 16776 19616 16788
rect 19475 16748 19616 16776
rect 19475 16745 19487 16748
rect 19429 16739 19487 16745
rect 19610 16736 19616 16748
rect 19668 16736 19674 16788
rect 19797 16779 19855 16785
rect 19797 16745 19809 16779
rect 19843 16776 19855 16779
rect 20070 16776 20076 16788
rect 19843 16748 20076 16776
rect 19843 16745 19855 16748
rect 19797 16739 19855 16745
rect 20070 16736 20076 16748
rect 20128 16736 20134 16788
rect 8196 16711 8254 16717
rect 6104 16680 7420 16708
rect 1854 16600 1860 16652
rect 1912 16640 1918 16652
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 1912 16612 2973 16640
rect 1912 16600 1918 16612
rect 2961 16609 2973 16612
rect 3007 16609 3019 16643
rect 3252 16640 3280 16668
rect 2961 16603 3019 16609
rect 3068 16612 3280 16640
rect 3068 16581 3096 16612
rect 3418 16600 3424 16652
rect 3476 16640 3482 16652
rect 4525 16643 4583 16649
rect 4525 16640 4537 16643
rect 3476 16612 4537 16640
rect 3476 16600 3482 16612
rect 4525 16609 4537 16612
rect 4571 16609 4583 16643
rect 5350 16640 5356 16652
rect 4525 16603 4583 16609
rect 5276 16612 5356 16640
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16541 2283 16575
rect 2225 16535 2283 16541
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16541 3111 16575
rect 3053 16535 3111 16541
rect 3237 16575 3295 16581
rect 3237 16541 3249 16575
rect 3283 16572 3295 16575
rect 3326 16572 3332 16584
rect 3283 16544 3332 16572
rect 3283 16541 3295 16544
rect 3237 16535 3295 16541
rect 2240 16504 2268 16535
rect 2406 16504 2412 16516
rect 2240 16476 2412 16504
rect 2406 16464 2412 16476
rect 2464 16504 2470 16516
rect 3252 16504 3280 16535
rect 3326 16532 3332 16544
rect 3384 16572 3390 16584
rect 4709 16575 4767 16581
rect 4709 16572 4721 16575
rect 3384 16544 4721 16572
rect 3384 16532 3390 16544
rect 4709 16541 4721 16544
rect 4755 16572 4767 16575
rect 5166 16572 5172 16584
rect 4755 16544 5172 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 5166 16532 5172 16544
rect 5224 16532 5230 16584
rect 5276 16581 5304 16612
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 5534 16649 5540 16652
rect 5528 16640 5540 16649
rect 5495 16612 5540 16640
rect 5528 16603 5540 16612
rect 5534 16600 5540 16603
rect 5592 16600 5598 16652
rect 7282 16640 7288 16652
rect 7243 16612 7288 16640
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 7392 16640 7420 16680
rect 8196 16677 8208 16711
rect 8242 16708 8254 16711
rect 8294 16708 8300 16720
rect 8242 16680 8300 16708
rect 8242 16677 8254 16680
rect 8196 16671 8254 16677
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 10962 16708 10968 16720
rect 8404 16680 10968 16708
rect 8404 16640 8432 16680
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 12066 16668 12072 16720
rect 12124 16708 12130 16720
rect 13256 16711 13314 16717
rect 12124 16680 12296 16708
rect 12124 16668 12130 16680
rect 9950 16640 9956 16652
rect 7392 16612 8432 16640
rect 9911 16612 9956 16640
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16640 10563 16643
rect 10594 16640 10600 16652
rect 10551 16612 10600 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 10772 16643 10830 16649
rect 10772 16609 10784 16643
rect 10818 16640 10830 16643
rect 11882 16640 11888 16652
rect 10818 16612 11888 16640
rect 10818 16609 10830 16612
rect 10772 16603 10830 16609
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 11974 16600 11980 16652
rect 12032 16640 12038 16652
rect 12161 16643 12219 16649
rect 12161 16640 12173 16643
rect 12032 16612 12173 16640
rect 12032 16600 12038 16612
rect 12161 16609 12173 16612
rect 12207 16609 12219 16643
rect 12268 16640 12296 16680
rect 13256 16677 13268 16711
rect 13302 16708 13314 16711
rect 13302 16680 15424 16708
rect 13302 16677 13314 16680
rect 13256 16671 13314 16677
rect 14366 16640 14372 16652
rect 12268 16612 14372 16640
rect 12161 16603 12219 16609
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 14550 16600 14556 16652
rect 14608 16640 14614 16652
rect 14645 16643 14703 16649
rect 14645 16640 14657 16643
rect 14608 16612 14657 16640
rect 14608 16600 14614 16612
rect 14645 16609 14657 16612
rect 14691 16609 14703 16643
rect 15396 16640 15424 16680
rect 15470 16668 15476 16720
rect 15528 16708 15534 16720
rect 17681 16711 17739 16717
rect 17681 16708 17693 16711
rect 15528 16680 17693 16708
rect 15528 16668 15534 16680
rect 17681 16677 17693 16680
rect 17727 16677 17739 16711
rect 17681 16671 17739 16677
rect 18046 16668 18052 16720
rect 18104 16708 18110 16720
rect 18693 16711 18751 16717
rect 18693 16708 18705 16711
rect 18104 16680 18705 16708
rect 18104 16668 18110 16680
rect 18693 16677 18705 16680
rect 18739 16677 18751 16711
rect 18693 16671 18751 16677
rect 18966 16668 18972 16720
rect 19024 16668 19030 16720
rect 19150 16668 19156 16720
rect 19208 16708 19214 16720
rect 19208 16680 20116 16708
rect 19208 16668 19214 16680
rect 15654 16640 15660 16652
rect 15396 16612 15516 16640
rect 15615 16612 15660 16640
rect 14645 16603 14703 16609
rect 5261 16575 5319 16581
rect 5261 16541 5273 16575
rect 5307 16541 5319 16575
rect 7466 16572 7472 16584
rect 7427 16544 7472 16572
rect 5261 16535 5319 16541
rect 2464 16476 3280 16504
rect 2464 16464 2470 16476
rect 3878 16464 3884 16516
rect 3936 16504 3942 16516
rect 5276 16504 5304 16535
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 7650 16532 7656 16584
rect 7708 16572 7714 16584
rect 7929 16575 7987 16581
rect 7929 16572 7941 16575
rect 7708 16544 7941 16572
rect 7708 16532 7714 16544
rect 7929 16541 7941 16544
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 12894 16532 12900 16584
rect 12952 16572 12958 16584
rect 12989 16575 13047 16581
rect 12989 16572 13001 16575
rect 12952 16544 13001 16572
rect 12952 16532 12958 16544
rect 12989 16541 13001 16544
rect 13035 16541 13047 16575
rect 15488 16572 15516 16612
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 16482 16640 16488 16652
rect 15764 16612 16488 16640
rect 15764 16572 15792 16612
rect 16482 16600 16488 16612
rect 16540 16600 16546 16652
rect 16574 16600 16580 16652
rect 16632 16640 16638 16652
rect 16669 16643 16727 16649
rect 16669 16640 16681 16643
rect 16632 16612 16681 16640
rect 16632 16600 16638 16612
rect 16669 16609 16681 16612
rect 16715 16609 16727 16643
rect 17770 16640 17776 16652
rect 17731 16612 17776 16640
rect 16669 16603 16727 16609
rect 17770 16600 17776 16612
rect 17828 16600 17834 16652
rect 18785 16643 18843 16649
rect 18785 16640 18797 16643
rect 18708 16612 18797 16640
rect 15488 16544 15792 16572
rect 15933 16575 15991 16581
rect 12989 16535 13047 16541
rect 15933 16541 15945 16575
rect 15979 16572 15991 16575
rect 16022 16572 16028 16584
rect 15979 16544 16028 16572
rect 15979 16541 15991 16544
rect 15933 16535 15991 16541
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 16758 16572 16764 16584
rect 16719 16544 16764 16572
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16572 16911 16575
rect 17865 16575 17923 16581
rect 17865 16572 17877 16575
rect 16899 16544 17877 16572
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 17865 16541 17877 16544
rect 17911 16541 17923 16575
rect 17865 16535 17923 16541
rect 3936 16476 5304 16504
rect 3936 16464 3942 16476
rect 6270 16464 6276 16516
rect 6328 16504 6334 16516
rect 16040 16504 16068 16532
rect 16868 16504 16896 16535
rect 6328 16476 7052 16504
rect 16040 16476 16896 16504
rect 6328 16464 6334 16476
rect 6641 16439 6699 16445
rect 6641 16405 6653 16439
rect 6687 16436 6699 16439
rect 6914 16436 6920 16448
rect 6687 16408 6920 16436
rect 6687 16405 6699 16408
rect 6641 16399 6699 16405
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 7024 16436 7052 16476
rect 8570 16436 8576 16448
rect 7024 16408 8576 16436
rect 8570 16396 8576 16408
rect 8628 16396 8634 16448
rect 8846 16396 8852 16448
rect 8904 16436 8910 16448
rect 11790 16436 11796 16448
rect 8904 16408 11796 16436
rect 8904 16396 8910 16408
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 11885 16439 11943 16445
rect 11885 16405 11897 16439
rect 11931 16436 11943 16439
rect 12986 16436 12992 16448
rect 11931 16408 12992 16436
rect 11931 16405 11943 16408
rect 11885 16399 11943 16405
rect 12986 16396 12992 16408
rect 13044 16396 13050 16448
rect 14090 16396 14096 16448
rect 14148 16436 14154 16448
rect 14369 16439 14427 16445
rect 14369 16436 14381 16439
rect 14148 16408 14381 16436
rect 14148 16396 14154 16408
rect 14369 16405 14381 16408
rect 14415 16405 14427 16439
rect 14369 16399 14427 16405
rect 14829 16439 14887 16445
rect 14829 16405 14841 16439
rect 14875 16436 14887 16439
rect 18598 16436 18604 16448
rect 14875 16408 18604 16436
rect 14875 16405 14887 16408
rect 14829 16399 14887 16405
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 18708 16436 18736 16612
rect 18785 16609 18797 16612
rect 18831 16609 18843 16643
rect 18984 16640 19012 16668
rect 20088 16652 20116 16680
rect 19889 16643 19947 16649
rect 19889 16640 19901 16643
rect 18984 16612 19901 16640
rect 18785 16603 18843 16609
rect 19889 16609 19901 16612
rect 19935 16609 19947 16643
rect 19889 16603 19947 16609
rect 20070 16600 20076 16652
rect 20128 16600 20134 16652
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16541 18935 16575
rect 18877 16535 18935 16541
rect 18782 16464 18788 16516
rect 18840 16504 18846 16516
rect 18892 16504 18920 16535
rect 19242 16532 19248 16584
rect 19300 16572 19306 16584
rect 19981 16575 20039 16581
rect 19981 16572 19993 16575
rect 19300 16544 19993 16572
rect 19300 16532 19306 16544
rect 19981 16541 19993 16544
rect 20027 16541 20039 16575
rect 19981 16535 20039 16541
rect 18840 16476 18920 16504
rect 18840 16464 18846 16476
rect 18966 16436 18972 16448
rect 18708 16408 18972 16436
rect 18966 16396 18972 16408
rect 19024 16436 19030 16448
rect 20622 16436 20628 16448
rect 19024 16408 20628 16436
rect 19024 16396 19030 16408
rect 20622 16396 20628 16408
rect 20680 16396 20686 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1486 16192 1492 16244
rect 1544 16232 1550 16244
rect 1673 16235 1731 16241
rect 1673 16232 1685 16235
rect 1544 16204 1685 16232
rect 1544 16192 1550 16204
rect 1673 16201 1685 16204
rect 1719 16201 1731 16235
rect 1673 16195 1731 16201
rect 2777 16235 2835 16241
rect 2777 16201 2789 16235
rect 2823 16232 2835 16235
rect 4706 16232 4712 16244
rect 2823 16204 4712 16232
rect 2823 16201 2835 16204
rect 2777 16195 2835 16201
rect 4706 16192 4712 16204
rect 4764 16192 4770 16244
rect 5350 16192 5356 16244
rect 5408 16232 5414 16244
rect 5994 16232 6000 16244
rect 5408 16204 5856 16232
rect 5955 16204 6000 16232
rect 5408 16192 5414 16204
rect 3789 16167 3847 16173
rect 3789 16133 3801 16167
rect 3835 16164 3847 16167
rect 5442 16164 5448 16176
rect 3835 16136 5448 16164
rect 3835 16133 3847 16136
rect 3789 16127 3847 16133
rect 5442 16124 5448 16136
rect 5500 16124 5506 16176
rect 5828 16164 5856 16204
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 7466 16192 7472 16244
rect 7524 16232 7530 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 7524 16204 8217 16232
rect 7524 16192 7530 16204
rect 8205 16201 8217 16204
rect 8251 16201 8263 16235
rect 8205 16195 8263 16201
rect 9493 16235 9551 16241
rect 9493 16201 9505 16235
rect 9539 16232 9551 16235
rect 10134 16232 10140 16244
rect 9539 16204 10140 16232
rect 9539 16201 9551 16204
rect 9493 16195 9551 16201
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 10376 16204 11744 16232
rect 10376 16192 10382 16204
rect 6365 16167 6423 16173
rect 6365 16164 6377 16167
rect 5828 16136 6377 16164
rect 6365 16133 6377 16136
rect 6411 16133 6423 16167
rect 6365 16127 6423 16133
rect 8481 16167 8539 16173
rect 8481 16133 8493 16167
rect 8527 16164 8539 16167
rect 10502 16164 10508 16176
rect 8527 16136 10508 16164
rect 8527 16133 8539 16136
rect 8481 16127 8539 16133
rect 10502 16124 10508 16136
rect 10560 16124 10566 16176
rect 3326 16096 3332 16108
rect 3287 16068 3332 16096
rect 3326 16056 3332 16068
rect 3384 16056 3390 16108
rect 4246 16056 4252 16108
rect 4304 16096 4310 16108
rect 4341 16099 4399 16105
rect 4341 16096 4353 16099
rect 4304 16068 4353 16096
rect 4304 16056 4310 16068
rect 4341 16065 4353 16068
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 5166 16056 5172 16108
rect 5224 16096 5230 16108
rect 5353 16099 5411 16105
rect 5353 16096 5365 16099
rect 5224 16068 5365 16096
rect 5224 16056 5230 16068
rect 5353 16065 5365 16068
rect 5399 16065 5411 16099
rect 5353 16059 5411 16065
rect 5626 16056 5632 16108
rect 5684 16096 5690 16108
rect 9125 16099 9183 16105
rect 5684 16068 6960 16096
rect 5684 16056 5690 16068
rect 1486 16028 1492 16040
rect 1447 16000 1492 16028
rect 1486 15988 1492 16000
rect 1544 15988 1550 16040
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 16028 2099 16031
rect 2130 16028 2136 16040
rect 2087 16000 2136 16028
rect 2087 15997 2099 16000
rect 2041 15991 2099 15997
rect 2130 15988 2136 16000
rect 2188 15988 2194 16040
rect 2314 16028 2320 16040
rect 2275 16000 2320 16028
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 4154 16028 4160 16040
rect 4115 16000 4160 16028
rect 4154 15988 4160 16000
rect 4212 15988 4218 16040
rect 5813 16031 5871 16037
rect 5813 15997 5825 16031
rect 5859 16028 5871 16031
rect 6270 16028 6276 16040
rect 5859 16000 6276 16028
rect 5859 15997 5871 16000
rect 5813 15991 5871 15997
rect 6270 15988 6276 16000
rect 6328 15988 6334 16040
rect 6454 15988 6460 16040
rect 6512 16028 6518 16040
rect 6549 16031 6607 16037
rect 6549 16028 6561 16031
rect 6512 16000 6561 16028
rect 6512 15988 6518 16000
rect 6549 15997 6561 16000
rect 6595 15997 6607 16031
rect 6549 15991 6607 15997
rect 6638 15988 6644 16040
rect 6696 16028 6702 16040
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6696 16000 6837 16028
rect 6696 15988 6702 16000
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 6932 16028 6960 16068
rect 9125 16065 9137 16099
rect 9171 16096 9183 16099
rect 9582 16096 9588 16108
rect 9171 16068 9588 16096
rect 9171 16065 9183 16068
rect 9125 16059 9183 16065
rect 9582 16056 9588 16068
rect 9640 16096 9646 16108
rect 10045 16099 10103 16105
rect 10045 16096 10057 16099
rect 9640 16068 10057 16096
rect 9640 16056 9646 16068
rect 10045 16065 10057 16068
rect 10091 16065 10103 16099
rect 11716 16096 11744 16204
rect 12158 16192 12164 16244
rect 12216 16232 12222 16244
rect 12437 16235 12495 16241
rect 12437 16232 12449 16235
rect 12216 16204 12449 16232
rect 12216 16192 12222 16204
rect 12437 16201 12449 16204
rect 12483 16201 12495 16235
rect 13814 16232 13820 16244
rect 12437 16195 12495 16201
rect 12544 16204 13820 16232
rect 11790 16124 11796 16176
rect 11848 16164 11854 16176
rect 12544 16164 12572 16204
rect 13814 16192 13820 16204
rect 13872 16232 13878 16244
rect 14366 16232 14372 16244
rect 13872 16204 14372 16232
rect 13872 16192 13878 16204
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 14553 16235 14611 16241
rect 14553 16201 14565 16235
rect 14599 16232 14611 16235
rect 15010 16232 15016 16244
rect 14599 16204 15016 16232
rect 14599 16201 14611 16204
rect 14553 16195 14611 16201
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 15565 16235 15623 16241
rect 15565 16201 15577 16235
rect 15611 16232 15623 16235
rect 15654 16232 15660 16244
rect 15611 16204 15660 16232
rect 15611 16201 15623 16204
rect 15565 16195 15623 16201
rect 15654 16192 15660 16204
rect 15712 16192 15718 16244
rect 16577 16235 16635 16241
rect 16577 16201 16589 16235
rect 16623 16232 16635 16235
rect 16758 16232 16764 16244
rect 16623 16204 16764 16232
rect 16623 16201 16635 16204
rect 16577 16195 16635 16201
rect 16758 16192 16764 16204
rect 16816 16192 16822 16244
rect 17586 16192 17592 16244
rect 17644 16232 17650 16244
rect 20073 16235 20131 16241
rect 20073 16232 20085 16235
rect 17644 16204 20085 16232
rect 17644 16192 17650 16204
rect 20073 16201 20085 16204
rect 20119 16201 20131 16235
rect 20073 16195 20131 16201
rect 11848 16136 12572 16164
rect 11848 16124 11854 16136
rect 13538 16124 13544 16176
rect 13596 16164 13602 16176
rect 19061 16167 19119 16173
rect 13596 16136 18552 16164
rect 13596 16124 13602 16136
rect 12986 16096 12992 16108
rect 11716 16068 12020 16096
rect 12947 16068 12992 16096
rect 10045 16059 10103 16065
rect 8754 16028 8760 16040
rect 6932 16000 8760 16028
rect 6825 15991 6883 15997
rect 8754 15988 8760 16000
rect 8812 15988 8818 16040
rect 10505 16031 10563 16037
rect 10505 15997 10517 16031
rect 10551 16028 10563 16031
rect 10594 16028 10600 16040
rect 10551 16000 10600 16028
rect 10551 15997 10563 16000
rect 10505 15991 10563 15997
rect 10594 15988 10600 16000
rect 10652 16028 10658 16040
rect 11238 16028 11244 16040
rect 10652 16000 11244 16028
rect 10652 15988 10658 16000
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 11330 15988 11336 16040
rect 11388 16028 11394 16040
rect 11992 16028 12020 16068
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 13262 16056 13268 16108
rect 13320 16096 13326 16108
rect 13909 16099 13967 16105
rect 13909 16096 13921 16099
rect 13320 16068 13921 16096
rect 13320 16056 13326 16068
rect 13909 16065 13921 16068
rect 13955 16065 13967 16099
rect 14090 16096 14096 16108
rect 14051 16068 14096 16096
rect 13909 16059 13967 16065
rect 14090 16056 14096 16068
rect 14148 16056 14154 16108
rect 15194 16096 15200 16108
rect 15155 16068 15200 16096
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 15286 16056 15292 16108
rect 15344 16096 15350 16108
rect 18524 16105 18552 16136
rect 19061 16133 19073 16167
rect 19107 16133 19119 16167
rect 19061 16127 19119 16133
rect 16209 16099 16267 16105
rect 16209 16096 16221 16099
rect 15344 16068 16221 16096
rect 15344 16056 15350 16068
rect 16209 16065 16221 16068
rect 16255 16096 16267 16099
rect 17129 16099 17187 16105
rect 17129 16096 17141 16099
rect 16255 16068 17141 16096
rect 16255 16065 16267 16068
rect 16209 16059 16267 16065
rect 17129 16065 17141 16068
rect 17175 16065 17187 16099
rect 17129 16059 17187 16065
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16065 18567 16099
rect 18509 16059 18567 16065
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16096 18751 16099
rect 18782 16096 18788 16108
rect 18739 16068 18788 16096
rect 18739 16065 18751 16068
rect 18693 16059 18751 16065
rect 18782 16056 18788 16068
rect 18840 16056 18846 16108
rect 18969 16099 19027 16105
rect 18969 16065 18981 16099
rect 19015 16096 19027 16099
rect 19076 16096 19104 16127
rect 19242 16124 19248 16176
rect 19300 16164 19306 16176
rect 19300 16136 20668 16164
rect 19300 16124 19306 16136
rect 19015 16068 19104 16096
rect 19015 16065 19027 16068
rect 18969 16059 19027 16065
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 19613 16099 19671 16105
rect 19613 16096 19625 16099
rect 19392 16068 19625 16096
rect 19392 16056 19398 16068
rect 19613 16065 19625 16068
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 20346 16056 20352 16108
rect 20404 16096 20410 16108
rect 20640 16105 20668 16136
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 20404 16068 20545 16096
rect 20404 16056 20410 16068
rect 20533 16065 20545 16068
rect 20579 16065 20591 16099
rect 20533 16059 20591 16065
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16065 20683 16099
rect 20625 16059 20683 16065
rect 13817 16031 13875 16037
rect 13817 16028 13829 16031
rect 11388 16000 11928 16028
rect 11992 16000 13829 16028
rect 11388 15988 11394 16000
rect 1394 15920 1400 15972
rect 1452 15960 1458 15972
rect 3145 15963 3203 15969
rect 3145 15960 3157 15963
rect 1452 15932 3157 15960
rect 1452 15920 1458 15932
rect 3145 15929 3157 15932
rect 3191 15960 3203 15963
rect 4706 15960 4712 15972
rect 3191 15932 4712 15960
rect 3191 15929 3203 15932
rect 3145 15923 3203 15929
rect 4706 15920 4712 15932
rect 4764 15920 4770 15972
rect 6914 15920 6920 15972
rect 6972 15960 6978 15972
rect 7092 15963 7150 15969
rect 7092 15960 7104 15963
rect 6972 15932 7104 15960
rect 6972 15920 6978 15932
rect 7092 15929 7104 15932
rect 7138 15960 7150 15963
rect 8202 15960 8208 15972
rect 7138 15932 8208 15960
rect 7138 15929 7150 15932
rect 7092 15923 7150 15929
rect 8202 15920 8208 15932
rect 8260 15920 8266 15972
rect 8386 15920 8392 15972
rect 8444 15960 8450 15972
rect 8941 15963 8999 15969
rect 8941 15960 8953 15963
rect 8444 15932 8953 15960
rect 8444 15920 8450 15932
rect 8941 15929 8953 15932
rect 8987 15929 8999 15963
rect 8941 15923 8999 15929
rect 10772 15963 10830 15969
rect 10772 15929 10784 15963
rect 10818 15960 10830 15963
rect 11790 15960 11796 15972
rect 10818 15932 11796 15960
rect 10818 15929 10830 15932
rect 10772 15923 10830 15929
rect 11790 15920 11796 15932
rect 11848 15920 11854 15972
rect 11900 15960 11928 16000
rect 13817 15997 13829 16000
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 14921 16031 14979 16037
rect 14921 15997 14933 16031
rect 14967 16028 14979 16031
rect 16390 16028 16396 16040
rect 14967 16000 16396 16028
rect 14967 15997 14979 16000
rect 14921 15991 14979 15997
rect 16390 15988 16396 16000
rect 16448 15988 16454 16040
rect 16666 15988 16672 16040
rect 16724 16028 16730 16040
rect 19242 16028 19248 16040
rect 16724 16000 19248 16028
rect 16724 15988 16730 16000
rect 19242 15988 19248 16000
rect 19300 15988 19306 16040
rect 19978 15988 19984 16040
rect 20036 16028 20042 16040
rect 20441 16031 20499 16037
rect 20441 16028 20453 16031
rect 20036 16000 20453 16028
rect 20036 15988 20042 16000
rect 20441 15997 20453 16000
rect 20487 15997 20499 16031
rect 20441 15991 20499 15997
rect 12897 15963 12955 15969
rect 12897 15960 12909 15963
rect 11900 15932 12909 15960
rect 12897 15929 12909 15932
rect 12943 15929 12955 15963
rect 17954 15960 17960 15972
rect 12897 15923 12955 15929
rect 13464 15932 17960 15960
rect 3234 15852 3240 15904
rect 3292 15892 3298 15904
rect 4249 15895 4307 15901
rect 3292 15864 3337 15892
rect 3292 15852 3298 15864
rect 4249 15861 4261 15895
rect 4295 15892 4307 15895
rect 4801 15895 4859 15901
rect 4801 15892 4813 15895
rect 4295 15864 4813 15892
rect 4295 15861 4307 15864
rect 4249 15855 4307 15861
rect 4801 15861 4813 15864
rect 4847 15861 4859 15895
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 4801 15855 4859 15861
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5261 15895 5319 15901
rect 5261 15861 5273 15895
rect 5307 15892 5319 15895
rect 6730 15892 6736 15904
rect 5307 15864 6736 15892
rect 5307 15861 5319 15864
rect 5261 15855 5319 15861
rect 6730 15852 6736 15864
rect 6788 15852 6794 15904
rect 6822 15852 6828 15904
rect 6880 15892 6886 15904
rect 7650 15892 7656 15904
rect 6880 15864 7656 15892
rect 6880 15852 6886 15864
rect 7650 15852 7656 15864
rect 7708 15852 7714 15904
rect 8846 15892 8852 15904
rect 8807 15864 8852 15892
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 9861 15895 9919 15901
rect 9861 15892 9873 15895
rect 9732 15864 9873 15892
rect 9732 15852 9738 15864
rect 9861 15861 9873 15864
rect 9907 15861 9919 15895
rect 9861 15855 9919 15861
rect 9953 15895 10011 15901
rect 9953 15861 9965 15895
rect 9999 15892 10011 15895
rect 10870 15892 10876 15904
rect 9999 15864 10876 15892
rect 9999 15861 10011 15864
rect 9953 15855 10011 15861
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 11882 15892 11888 15904
rect 11843 15864 11888 15892
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 12710 15852 12716 15904
rect 12768 15892 12774 15904
rect 13464 15901 13492 15932
rect 17954 15920 17960 15932
rect 18012 15920 18018 15972
rect 19521 15963 19579 15969
rect 19521 15960 19533 15963
rect 18064 15932 19104 15960
rect 12805 15895 12863 15901
rect 12805 15892 12817 15895
rect 12768 15864 12817 15892
rect 12768 15852 12774 15864
rect 12805 15861 12817 15864
rect 12851 15861 12863 15895
rect 12805 15855 12863 15861
rect 13449 15895 13507 15901
rect 13449 15861 13461 15895
rect 13495 15861 13507 15895
rect 13449 15855 13507 15861
rect 15013 15895 15071 15901
rect 15013 15861 15025 15895
rect 15059 15892 15071 15895
rect 15286 15892 15292 15904
rect 15059 15864 15292 15892
rect 15059 15861 15071 15864
rect 15013 15855 15071 15861
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 15746 15852 15752 15904
rect 15804 15892 15810 15904
rect 15933 15895 15991 15901
rect 15933 15892 15945 15895
rect 15804 15864 15945 15892
rect 15804 15852 15810 15864
rect 15933 15861 15945 15864
rect 15979 15861 15991 15895
rect 15933 15855 15991 15861
rect 16025 15895 16083 15901
rect 16025 15861 16037 15895
rect 16071 15892 16083 15895
rect 16206 15892 16212 15904
rect 16071 15864 16212 15892
rect 16071 15861 16083 15864
rect 16025 15855 16083 15861
rect 16206 15852 16212 15864
rect 16264 15852 16270 15904
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 16945 15895 17003 15901
rect 16945 15892 16957 15895
rect 16908 15864 16957 15892
rect 16908 15852 16914 15864
rect 16945 15861 16957 15864
rect 16991 15861 17003 15895
rect 16945 15855 17003 15861
rect 17037 15895 17095 15901
rect 17037 15861 17049 15895
rect 17083 15892 17095 15895
rect 17126 15892 17132 15904
rect 17083 15864 17132 15892
rect 17083 15861 17095 15864
rect 17037 15855 17095 15861
rect 17126 15852 17132 15864
rect 17184 15852 17190 15904
rect 18064 15901 18092 15932
rect 18049 15895 18107 15901
rect 18049 15861 18061 15895
rect 18095 15861 18107 15895
rect 18049 15855 18107 15861
rect 18138 15852 18144 15904
rect 18196 15892 18202 15904
rect 18417 15895 18475 15901
rect 18417 15892 18429 15895
rect 18196 15864 18429 15892
rect 18196 15852 18202 15864
rect 18417 15861 18429 15864
rect 18463 15861 18475 15895
rect 18417 15855 18475 15861
rect 18506 15852 18512 15904
rect 18564 15892 18570 15904
rect 18969 15895 19027 15901
rect 18969 15892 18981 15895
rect 18564 15864 18981 15892
rect 18564 15852 18570 15864
rect 18969 15861 18981 15864
rect 19015 15861 19027 15895
rect 19076 15892 19104 15932
rect 19260 15932 19533 15960
rect 19260 15892 19288 15932
rect 19521 15929 19533 15932
rect 19567 15929 19579 15963
rect 19521 15923 19579 15929
rect 19076 15864 19288 15892
rect 18969 15855 19027 15861
rect 19334 15852 19340 15904
rect 19392 15892 19398 15904
rect 19429 15895 19487 15901
rect 19429 15892 19441 15895
rect 19392 15864 19441 15892
rect 19392 15852 19398 15864
rect 19429 15861 19441 15864
rect 19475 15861 19487 15895
rect 19429 15855 19487 15861
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1578 15688 1584 15700
rect 1539 15660 1584 15688
rect 1578 15648 1584 15660
rect 1636 15648 1642 15700
rect 1949 15691 2007 15697
rect 1949 15657 1961 15691
rect 1995 15657 2007 15691
rect 1949 15651 2007 15657
rect 2317 15691 2375 15697
rect 2317 15657 2329 15691
rect 2363 15688 2375 15691
rect 2406 15688 2412 15700
rect 2363 15660 2412 15688
rect 2363 15657 2375 15660
rect 2317 15651 2375 15657
rect 1964 15620 1992 15651
rect 2406 15648 2412 15660
rect 2464 15648 2470 15700
rect 3421 15691 3479 15697
rect 3421 15657 3433 15691
rect 3467 15688 3479 15691
rect 3510 15688 3516 15700
rect 3467 15660 3516 15688
rect 3467 15657 3479 15660
rect 3421 15651 3479 15657
rect 3510 15648 3516 15660
rect 3568 15648 3574 15700
rect 4062 15648 4068 15700
rect 4120 15688 4126 15700
rect 4709 15691 4767 15697
rect 4120 15660 4384 15688
rect 4120 15648 4126 15660
rect 4356 15620 4384 15660
rect 4709 15657 4721 15691
rect 4755 15688 4767 15691
rect 5353 15691 5411 15697
rect 5353 15688 5365 15691
rect 4755 15660 5365 15688
rect 4755 15657 4767 15660
rect 4709 15651 4767 15657
rect 5353 15657 5365 15660
rect 5399 15657 5411 15691
rect 5353 15651 5411 15657
rect 5718 15648 5724 15700
rect 5776 15688 5782 15700
rect 6178 15688 6184 15700
rect 5776 15660 6184 15688
rect 5776 15648 5782 15660
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 6549 15691 6607 15697
rect 6549 15657 6561 15691
rect 6595 15688 6607 15691
rect 7190 15688 7196 15700
rect 6595 15660 7196 15688
rect 6595 15657 6607 15660
rect 6549 15651 6607 15657
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 7282 15648 7288 15700
rect 7340 15688 7346 15700
rect 7561 15691 7619 15697
rect 7561 15688 7573 15691
rect 7340 15660 7573 15688
rect 7340 15648 7346 15660
rect 7561 15657 7573 15660
rect 7607 15657 7619 15691
rect 7561 15651 7619 15657
rect 7650 15648 7656 15700
rect 7708 15688 7714 15700
rect 8021 15691 8079 15697
rect 8021 15688 8033 15691
rect 7708 15660 8033 15688
rect 7708 15648 7714 15660
rect 8021 15657 8033 15660
rect 8067 15657 8079 15691
rect 8021 15651 8079 15657
rect 8573 15691 8631 15697
rect 8573 15657 8585 15691
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 6086 15620 6092 15632
rect 1964 15592 4292 15620
rect 4356 15592 6092 15620
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 3234 15512 3240 15564
rect 3292 15552 3298 15564
rect 3329 15555 3387 15561
rect 3329 15552 3341 15555
rect 3292 15524 3341 15552
rect 3292 15512 3298 15524
rect 3329 15521 3341 15524
rect 3375 15521 3387 15555
rect 4264 15552 4292 15592
rect 6086 15580 6092 15592
rect 6144 15580 6150 15632
rect 6917 15623 6975 15629
rect 6917 15589 6929 15623
rect 6963 15620 6975 15623
rect 8588 15620 8616 15651
rect 8846 15648 8852 15700
rect 8904 15688 8910 15700
rect 12986 15688 12992 15700
rect 8904 15660 12992 15688
rect 8904 15648 8910 15660
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 14829 15691 14887 15697
rect 14829 15657 14841 15691
rect 14875 15657 14887 15691
rect 15286 15688 15292 15700
rect 15247 15660 15292 15688
rect 14829 15651 14887 15657
rect 6963 15592 8616 15620
rect 6963 15589 6975 15592
rect 6917 15583 6975 15589
rect 8754 15580 8760 15632
rect 8812 15620 8818 15632
rect 8941 15623 8999 15629
rect 8941 15620 8953 15623
rect 8812 15592 8953 15620
rect 8812 15580 8818 15592
rect 8941 15589 8953 15592
rect 8987 15589 8999 15623
rect 8941 15583 8999 15589
rect 9033 15623 9091 15629
rect 9033 15589 9045 15623
rect 9079 15620 9091 15623
rect 9214 15620 9220 15632
rect 9079 15592 9220 15620
rect 9079 15589 9091 15592
rect 9033 15583 9091 15589
rect 9214 15580 9220 15592
rect 9272 15580 9278 15632
rect 11330 15620 11336 15632
rect 9600 15592 11336 15620
rect 4617 15555 4675 15561
rect 4264 15524 4568 15552
rect 3329 15515 3387 15521
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2409 15487 2467 15493
rect 2409 15484 2421 15487
rect 1820 15456 2421 15484
rect 1820 15444 1826 15456
rect 2409 15453 2421 15456
rect 2455 15453 2467 15487
rect 2590 15484 2596 15496
rect 2551 15456 2596 15484
rect 2409 15447 2467 15453
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 3602 15484 3608 15496
rect 3563 15456 3608 15484
rect 3602 15444 3608 15456
rect 3660 15444 3666 15496
rect 4540 15484 4568 15524
rect 4617 15521 4629 15555
rect 4663 15552 4675 15555
rect 5534 15552 5540 15564
rect 4663 15524 5540 15552
rect 4663 15521 4675 15524
rect 4617 15515 4675 15521
rect 5534 15512 5540 15524
rect 5592 15512 5598 15564
rect 5718 15552 5724 15564
rect 5679 15524 5724 15552
rect 5718 15512 5724 15524
rect 5776 15512 5782 15564
rect 5813 15555 5871 15561
rect 5813 15521 5825 15555
rect 5859 15552 5871 15555
rect 7558 15552 7564 15564
rect 5859 15524 7564 15552
rect 5859 15521 5871 15524
rect 5813 15515 5871 15521
rect 7558 15512 7564 15524
rect 7616 15512 7622 15564
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15521 7987 15555
rect 7929 15515 7987 15521
rect 4798 15484 4804 15496
rect 4540 15456 4660 15484
rect 4759 15456 4804 15484
rect 2961 15419 3019 15425
rect 2961 15385 2973 15419
rect 3007 15416 3019 15419
rect 4154 15416 4160 15428
rect 3007 15388 4160 15416
rect 3007 15385 3019 15388
rect 2961 15379 3019 15385
rect 4154 15376 4160 15388
rect 4212 15376 4218 15428
rect 4632 15416 4660 15456
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 5902 15484 5908 15496
rect 5863 15456 5908 15484
rect 5902 15444 5908 15456
rect 5960 15444 5966 15496
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15484 7067 15487
rect 7098 15484 7104 15496
rect 7055 15456 7104 15484
rect 7055 15453 7067 15456
rect 7009 15447 7067 15453
rect 7098 15444 7104 15456
rect 7156 15444 7162 15496
rect 7193 15487 7251 15493
rect 7193 15453 7205 15487
rect 7239 15484 7251 15487
rect 7466 15484 7472 15496
rect 7239 15456 7472 15484
rect 7239 15453 7251 15456
rect 7193 15447 7251 15453
rect 7466 15444 7472 15456
rect 7524 15444 7530 15496
rect 7944 15416 7972 15515
rect 8570 15512 8576 15564
rect 8628 15552 8634 15564
rect 8846 15552 8852 15564
rect 8628 15524 8852 15552
rect 8628 15512 8634 15524
rect 8846 15512 8852 15524
rect 8904 15512 8910 15564
rect 8202 15484 8208 15496
rect 8115 15456 8208 15484
rect 8202 15444 8208 15456
rect 8260 15484 8266 15496
rect 9217 15487 9275 15493
rect 9217 15484 9229 15487
rect 8260 15456 9229 15484
rect 8260 15444 8266 15456
rect 9217 15453 9229 15456
rect 9263 15484 9275 15487
rect 9306 15484 9312 15496
rect 9263 15456 9312 15484
rect 9263 15453 9275 15456
rect 9217 15447 9275 15453
rect 9306 15444 9312 15456
rect 9364 15444 9370 15496
rect 4632 15388 7972 15416
rect 8478 15376 8484 15428
rect 8536 15416 8542 15428
rect 9600 15416 9628 15592
rect 11330 15580 11336 15592
rect 11388 15580 11394 15632
rect 11508 15623 11566 15629
rect 11508 15589 11520 15623
rect 11554 15620 11566 15623
rect 14090 15620 14096 15632
rect 11554 15592 14096 15620
rect 11554 15589 11566 15592
rect 11508 15583 11566 15589
rect 14090 15580 14096 15592
rect 14148 15580 14154 15632
rect 14844 15620 14872 15651
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 16301 15691 16359 15697
rect 16301 15657 16313 15691
rect 16347 15688 16359 15691
rect 18230 15688 18236 15700
rect 16347 15660 18236 15688
rect 16347 15657 16359 15660
rect 16301 15651 16359 15657
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 18322 15648 18328 15700
rect 18380 15688 18386 15700
rect 18380 15660 18425 15688
rect 18380 15648 18386 15660
rect 18782 15648 18788 15700
rect 18840 15688 18846 15700
rect 19334 15688 19340 15700
rect 18840 15660 18920 15688
rect 19295 15660 19340 15688
rect 18840 15648 18846 15660
rect 17954 15620 17960 15632
rect 14844 15592 17960 15620
rect 17954 15580 17960 15592
rect 18012 15580 18018 15632
rect 18046 15580 18052 15632
rect 18104 15620 18110 15632
rect 18104 15592 18451 15620
rect 18104 15580 18110 15592
rect 10410 15552 10416 15564
rect 10371 15524 10416 15552
rect 10410 15512 10416 15524
rect 10468 15512 10474 15564
rect 11238 15552 11244 15564
rect 11151 15524 11244 15552
rect 11238 15512 11244 15524
rect 11296 15552 11302 15564
rect 11974 15552 11980 15564
rect 11296 15524 11980 15552
rect 11296 15512 11302 15524
rect 11974 15512 11980 15524
rect 12032 15552 12038 15564
rect 12713 15555 12771 15561
rect 12032 15524 12296 15552
rect 12032 15512 12038 15524
rect 10502 15484 10508 15496
rect 10463 15456 10508 15484
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 10686 15484 10692 15496
rect 10647 15456 10692 15484
rect 10686 15444 10692 15456
rect 10744 15444 10750 15496
rect 12268 15484 12296 15524
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 13164 15555 13222 15561
rect 13164 15552 13176 15555
rect 12759 15524 13176 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 13164 15521 13176 15524
rect 13210 15552 13222 15555
rect 13538 15552 13544 15564
rect 13210 15524 13544 15552
rect 13210 15521 13222 15524
rect 13164 15515 13222 15521
rect 13538 15512 13544 15524
rect 13596 15552 13602 15564
rect 14550 15552 14556 15564
rect 13596 15524 14556 15552
rect 13596 15512 13602 15524
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 14645 15555 14703 15561
rect 14645 15521 14657 15555
rect 14691 15552 14703 15555
rect 15010 15552 15016 15564
rect 14691 15524 15016 15552
rect 14691 15521 14703 15524
rect 14645 15515 14703 15521
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 15654 15552 15660 15564
rect 15396 15524 15660 15552
rect 12894 15484 12900 15496
rect 12268 15456 12900 15484
rect 12894 15444 12900 15456
rect 12952 15444 12958 15496
rect 13906 15444 13912 15496
rect 13964 15484 13970 15496
rect 15396 15484 15424 15524
rect 15654 15512 15660 15524
rect 15712 15512 15718 15564
rect 16666 15552 16672 15564
rect 16627 15524 16672 15552
rect 16666 15512 16672 15524
rect 16724 15512 16730 15564
rect 17678 15552 17684 15564
rect 17639 15524 17684 15552
rect 17678 15512 17684 15524
rect 17736 15512 17742 15564
rect 17773 15555 17831 15561
rect 17773 15521 17785 15555
rect 17819 15552 17831 15555
rect 18322 15552 18328 15564
rect 17819 15524 18328 15552
rect 17819 15521 17831 15524
rect 17773 15515 17831 15521
rect 18322 15512 18328 15524
rect 18380 15512 18386 15564
rect 18423 15552 18451 15592
rect 18690 15580 18696 15632
rect 18748 15620 18754 15632
rect 18748 15592 18793 15620
rect 18748 15580 18754 15592
rect 18785 15555 18843 15561
rect 18785 15552 18797 15555
rect 18423 15524 18797 15552
rect 18785 15521 18797 15524
rect 18831 15521 18843 15555
rect 18892 15552 18920 15660
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 19705 15623 19763 15629
rect 19705 15589 19717 15623
rect 19751 15620 19763 15623
rect 19794 15620 19800 15632
rect 19751 15592 19800 15620
rect 19751 15589 19763 15592
rect 19705 15583 19763 15589
rect 19794 15580 19800 15592
rect 19852 15580 19858 15632
rect 18892 15524 20024 15552
rect 18785 15515 18843 15521
rect 13964 15456 15424 15484
rect 13964 15444 13970 15456
rect 15470 15444 15476 15496
rect 15528 15484 15534 15496
rect 15749 15487 15807 15493
rect 15749 15484 15761 15487
rect 15528 15456 15761 15484
rect 15528 15444 15534 15456
rect 15749 15453 15761 15456
rect 15795 15453 15807 15487
rect 15749 15447 15807 15453
rect 15933 15487 15991 15493
rect 15933 15453 15945 15487
rect 15979 15484 15991 15487
rect 16022 15484 16028 15496
rect 15979 15456 16028 15484
rect 15979 15453 15991 15456
rect 15933 15447 15991 15453
rect 8536 15388 9628 15416
rect 12621 15419 12679 15425
rect 8536 15376 8542 15388
rect 12621 15385 12633 15419
rect 12667 15416 12679 15419
rect 12713 15419 12771 15425
rect 12713 15416 12725 15419
rect 12667 15388 12725 15416
rect 12667 15385 12679 15388
rect 12621 15379 12679 15385
rect 12713 15385 12725 15388
rect 12759 15385 12771 15419
rect 15764 15416 15792 15447
rect 16022 15444 16028 15456
rect 16080 15444 16086 15496
rect 16758 15484 16764 15496
rect 16719 15456 16764 15484
rect 16758 15444 16764 15456
rect 16816 15444 16822 15496
rect 16945 15487 17003 15493
rect 16945 15453 16957 15487
rect 16991 15484 17003 15487
rect 17862 15484 17868 15496
rect 16991 15456 17868 15484
rect 16991 15453 17003 15456
rect 16945 15447 17003 15453
rect 17862 15444 17868 15456
rect 17920 15444 17926 15496
rect 18969 15487 19027 15493
rect 18969 15484 18981 15487
rect 18423 15456 18981 15484
rect 16117 15419 16175 15425
rect 16117 15416 16129 15419
rect 15764 15388 16129 15416
rect 12713 15379 12771 15385
rect 16117 15385 16129 15388
rect 16163 15385 16175 15419
rect 18423 15416 18451 15456
rect 18969 15453 18981 15456
rect 19015 15453 19027 15487
rect 19242 15484 19248 15496
rect 18969 15447 19027 15453
rect 19168 15456 19248 15484
rect 16117 15379 16175 15385
rect 16224 15388 18451 15416
rect 4246 15348 4252 15360
rect 4207 15320 4252 15348
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 5166 15308 5172 15360
rect 5224 15348 5230 15360
rect 6914 15348 6920 15360
rect 5224 15320 6920 15348
rect 5224 15308 5230 15320
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 10045 15351 10103 15357
rect 10045 15317 10057 15351
rect 10091 15348 10103 15351
rect 12158 15348 12164 15360
rect 10091 15320 12164 15348
rect 10091 15317 10103 15320
rect 10045 15311 10103 15317
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 14277 15351 14335 15357
rect 14277 15317 14289 15351
rect 14323 15348 14335 15351
rect 14550 15348 14556 15360
rect 14323 15320 14556 15348
rect 14323 15317 14335 15320
rect 14277 15311 14335 15317
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 14642 15308 14648 15360
rect 14700 15348 14706 15360
rect 16224 15348 16252 15388
rect 14700 15320 16252 15348
rect 17313 15351 17371 15357
rect 14700 15308 14706 15320
rect 17313 15317 17325 15351
rect 17359 15348 17371 15351
rect 17954 15348 17960 15360
rect 17359 15320 17960 15348
rect 17359 15317 17371 15320
rect 17313 15311 17371 15317
rect 17954 15308 17960 15320
rect 18012 15308 18018 15360
rect 19168 15348 19196 15456
rect 19242 15444 19248 15456
rect 19300 15444 19306 15496
rect 19996 15493 20024 15524
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15453 19855 15487
rect 19797 15447 19855 15453
rect 19981 15487 20039 15493
rect 19981 15453 19993 15487
rect 20027 15484 20039 15487
rect 20622 15484 20628 15496
rect 20027 15456 20628 15484
rect 20027 15453 20039 15456
rect 19981 15447 20039 15453
rect 19812 15348 19840 15447
rect 20622 15444 20628 15456
rect 20680 15444 20686 15496
rect 19168 15320 19840 15348
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 3786 15144 3792 15156
rect 3436 15116 3792 15144
rect 3436 15017 3464 15116
rect 3786 15104 3792 15116
rect 3844 15104 3850 15156
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 6825 15147 6883 15153
rect 6825 15144 6837 15147
rect 5776 15116 6837 15144
rect 5776 15104 5782 15116
rect 6825 15113 6837 15116
rect 6871 15113 6883 15147
rect 6825 15107 6883 15113
rect 6914 15104 6920 15156
rect 6972 15144 6978 15156
rect 11790 15144 11796 15156
rect 6972 15116 11652 15144
rect 11751 15116 11796 15144
rect 6972 15104 6978 15116
rect 6086 15036 6092 15088
rect 6144 15076 6150 15088
rect 8021 15079 8079 15085
rect 8021 15076 8033 15079
rect 6144 15048 8033 15076
rect 6144 15036 6150 15048
rect 8021 15045 8033 15048
rect 8067 15045 8079 15079
rect 8021 15039 8079 15045
rect 8297 15079 8355 15085
rect 8297 15045 8309 15079
rect 8343 15076 8355 15079
rect 11624 15076 11652 15116
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 12437 15147 12495 15153
rect 12437 15113 12449 15147
rect 12483 15144 12495 15147
rect 12802 15144 12808 15156
rect 12483 15116 12808 15144
rect 12483 15113 12495 15116
rect 12437 15107 12495 15113
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 13817 15147 13875 15153
rect 13817 15113 13829 15147
rect 13863 15144 13875 15147
rect 17494 15144 17500 15156
rect 13863 15116 17500 15144
rect 13863 15113 13875 15116
rect 13817 15107 13875 15113
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 17589 15147 17647 15153
rect 17589 15113 17601 15147
rect 17635 15144 17647 15147
rect 17862 15144 17868 15156
rect 17635 15116 17868 15144
rect 17635 15113 17647 15116
rect 17589 15107 17647 15113
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 13170 15076 13176 15088
rect 8343 15048 8800 15076
rect 11624 15048 13176 15076
rect 8343 15045 8355 15048
rect 8297 15039 8355 15045
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 1765 14943 1823 14949
rect 1765 14909 1777 14943
rect 1811 14940 1823 14943
rect 3436 14940 3464 14971
rect 7190 14968 7196 15020
rect 7248 15008 7254 15020
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 7248 14980 7389 15008
rect 7248 14968 7254 14980
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 8110 14968 8116 15020
rect 8168 15008 8174 15020
rect 8772 15017 8800 15048
rect 13170 15036 13176 15048
rect 13228 15036 13234 15088
rect 18322 15076 18328 15088
rect 17880 15048 18328 15076
rect 8757 15011 8815 15017
rect 8168 14980 8616 15008
rect 8168 14968 8174 14980
rect 3688 14943 3746 14949
rect 3688 14940 3700 14943
rect 1811 14912 3464 14940
rect 3620 14912 3700 14940
rect 1811 14909 1823 14912
rect 1765 14903 1823 14909
rect 2240 14884 2268 14912
rect 2038 14881 2044 14884
rect 2032 14835 2044 14881
rect 2096 14872 2102 14884
rect 2096 14844 2132 14872
rect 2038 14832 2044 14835
rect 2096 14832 2102 14844
rect 2222 14832 2228 14884
rect 2280 14832 2286 14884
rect 3620 14872 3648 14912
rect 3688 14909 3700 14912
rect 3734 14940 3746 14943
rect 4798 14940 4804 14952
rect 3734 14912 4804 14940
rect 3734 14909 3746 14912
rect 3688 14903 3746 14909
rect 4798 14900 4804 14912
rect 4856 14900 4862 14952
rect 5074 14940 5080 14952
rect 5035 14912 5080 14940
rect 5074 14900 5080 14912
rect 5132 14900 5138 14952
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 8588 14949 8616 14980
rect 8757 14977 8769 15011
rect 8803 14977 8815 15011
rect 10413 15011 10471 15017
rect 10413 15008 10425 15011
rect 8757 14971 8815 14977
rect 9784 14980 10425 15008
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 5684 14912 7849 14940
rect 5684 14900 5690 14912
rect 7837 14909 7849 14912
rect 7883 14909 7895 14943
rect 7837 14903 7895 14909
rect 8573 14943 8631 14949
rect 8573 14909 8585 14943
rect 8619 14909 8631 14943
rect 8772 14940 8800 14971
rect 9784 14940 9812 14980
rect 10413 14977 10425 14980
rect 10459 14977 10471 15011
rect 10413 14971 10471 14977
rect 11882 14968 11888 15020
rect 11940 15008 11946 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 11940 14980 13001 15008
rect 11940 14968 11946 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 12253 14943 12311 14949
rect 8772 14912 9812 14940
rect 10522 14912 10815 14940
rect 8573 14903 8631 14909
rect 5350 14881 5356 14884
rect 5344 14872 5356 14881
rect 3160 14844 3648 14872
rect 5311 14844 5356 14872
rect 3160 14813 3188 14844
rect 5344 14835 5356 14844
rect 5350 14832 5356 14835
rect 5408 14832 5414 14884
rect 9024 14875 9082 14881
rect 9024 14841 9036 14875
rect 9070 14872 9082 14875
rect 9122 14872 9128 14884
rect 9070 14844 9128 14872
rect 9070 14841 9082 14844
rect 9024 14835 9082 14841
rect 9122 14832 9128 14844
rect 9180 14832 9186 14884
rect 9582 14832 9588 14884
rect 9640 14872 9646 14884
rect 10522 14872 10550 14912
rect 10686 14881 10692 14884
rect 10680 14872 10692 14881
rect 9640 14844 10550 14872
rect 10599 14844 10692 14872
rect 9640 14832 9646 14844
rect 10680 14835 10692 14844
rect 10686 14832 10692 14835
rect 10744 14832 10750 14884
rect 10787 14872 10815 14912
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 13262 14940 13268 14952
rect 12299 14912 13268 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13906 14940 13912 14952
rect 13679 14912 13912 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 13906 14900 13912 14912
rect 13964 14900 13970 14952
rect 14185 14943 14243 14949
rect 14185 14909 14197 14943
rect 14231 14909 14243 14943
rect 14185 14903 14243 14909
rect 12434 14872 12440 14884
rect 10787 14844 12440 14872
rect 12434 14832 12440 14844
rect 12492 14832 12498 14884
rect 14200 14872 14228 14903
rect 16022 14900 16028 14952
rect 16080 14940 16086 14952
rect 16209 14943 16267 14949
rect 16209 14940 16221 14943
rect 16080 14912 16221 14940
rect 16080 14900 16086 14912
rect 16209 14909 16221 14912
rect 16255 14909 16267 14943
rect 17880 14940 17908 15048
rect 18322 15036 18328 15048
rect 18380 15036 18386 15088
rect 18414 14968 18420 15020
rect 18472 15008 18478 15020
rect 18601 15011 18659 15017
rect 18601 15008 18613 15011
rect 18472 14980 18613 15008
rect 18472 14968 18478 14980
rect 18601 14977 18613 14980
rect 18647 14977 18659 15011
rect 19702 15008 19708 15020
rect 18601 14971 18659 14977
rect 18984 14980 19564 15008
rect 19663 14980 19708 15008
rect 16209 14903 16267 14909
rect 16408 14912 17908 14940
rect 13648 14844 14228 14872
rect 14452 14875 14510 14881
rect 3145 14807 3203 14813
rect 3145 14773 3157 14807
rect 3191 14773 3203 14807
rect 3145 14767 3203 14773
rect 3510 14764 3516 14816
rect 3568 14804 3574 14816
rect 4801 14807 4859 14813
rect 4801 14804 4813 14807
rect 3568 14776 4813 14804
rect 3568 14764 3574 14776
rect 4801 14773 4813 14776
rect 4847 14804 4859 14807
rect 5442 14804 5448 14816
rect 4847 14776 5448 14804
rect 4847 14773 4859 14776
rect 4801 14767 4859 14773
rect 5442 14764 5448 14776
rect 5500 14764 5506 14816
rect 5902 14764 5908 14816
rect 5960 14804 5966 14816
rect 6457 14807 6515 14813
rect 6457 14804 6469 14807
rect 5960 14776 6469 14804
rect 5960 14764 5966 14776
rect 6457 14773 6469 14776
rect 6503 14773 6515 14807
rect 6457 14767 6515 14773
rect 6914 14764 6920 14816
rect 6972 14804 6978 14816
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 6972 14776 7205 14804
rect 6972 14764 6978 14776
rect 7193 14773 7205 14776
rect 7239 14773 7251 14807
rect 7193 14767 7251 14773
rect 7285 14807 7343 14813
rect 7285 14773 7297 14807
rect 7331 14804 7343 14807
rect 7466 14804 7472 14816
rect 7331 14776 7472 14804
rect 7331 14773 7343 14776
rect 7285 14767 7343 14773
rect 7466 14764 7472 14776
rect 7524 14764 7530 14816
rect 7650 14764 7656 14816
rect 7708 14804 7714 14816
rect 8297 14807 8355 14813
rect 8297 14804 8309 14807
rect 7708 14776 8309 14804
rect 7708 14764 7714 14776
rect 8297 14773 8309 14776
rect 8343 14804 8355 14807
rect 8389 14807 8447 14813
rect 8389 14804 8401 14807
rect 8343 14776 8401 14804
rect 8343 14773 8355 14776
rect 8297 14767 8355 14773
rect 8389 14773 8401 14776
rect 8435 14773 8447 14807
rect 8389 14767 8447 14773
rect 10137 14807 10195 14813
rect 10137 14773 10149 14807
rect 10183 14804 10195 14807
rect 10695 14804 10723 14832
rect 13648 14816 13676 14844
rect 14452 14841 14464 14875
rect 14498 14872 14510 14875
rect 14550 14872 14556 14884
rect 14498 14844 14556 14872
rect 14498 14841 14510 14844
rect 14452 14835 14510 14841
rect 14550 14832 14556 14844
rect 14608 14832 14614 14884
rect 15286 14832 15292 14884
rect 15344 14872 15350 14884
rect 16408 14872 16436 14912
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 18012 14912 18460 14940
rect 18012 14900 18018 14912
rect 15344 14844 16436 14872
rect 16476 14875 16534 14881
rect 15344 14832 15350 14844
rect 16476 14841 16488 14875
rect 16522 14872 16534 14875
rect 17218 14872 17224 14884
rect 16522 14844 17224 14872
rect 16522 14841 16534 14844
rect 16476 14835 16534 14841
rect 17218 14832 17224 14844
rect 17276 14832 17282 14884
rect 18432 14881 18460 14912
rect 18506 14900 18512 14952
rect 18564 14940 18570 14952
rect 18564 14912 18609 14940
rect 18564 14900 18570 14912
rect 18417 14875 18475 14881
rect 17880 14844 18368 14872
rect 11882 14804 11888 14816
rect 10183 14776 11888 14804
rect 10183 14773 10195 14776
rect 10137 14767 10195 14773
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 11974 14764 11980 14816
rect 12032 14804 12038 14816
rect 12069 14807 12127 14813
rect 12069 14804 12081 14807
rect 12032 14776 12081 14804
rect 12032 14764 12038 14776
rect 12069 14773 12081 14776
rect 12115 14804 12127 14807
rect 12526 14804 12532 14816
rect 12115 14776 12532 14804
rect 12115 14773 12127 14776
rect 12069 14767 12127 14773
rect 12526 14764 12532 14776
rect 12584 14764 12590 14816
rect 12802 14804 12808 14816
rect 12763 14776 12808 14804
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 12897 14807 12955 14813
rect 12897 14773 12909 14807
rect 12943 14804 12955 14807
rect 13078 14804 13084 14816
rect 12943 14776 13084 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 13630 14764 13636 14816
rect 13688 14764 13694 14816
rect 15562 14804 15568 14816
rect 15523 14776 15568 14804
rect 15562 14764 15568 14776
rect 15620 14764 15626 14816
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 17880 14804 17908 14844
rect 16264 14776 17908 14804
rect 16264 14764 16270 14776
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18049 14807 18107 14813
rect 18049 14804 18061 14807
rect 18012 14776 18061 14804
rect 18012 14764 18018 14776
rect 18049 14773 18061 14776
rect 18095 14773 18107 14807
rect 18340 14804 18368 14844
rect 18417 14841 18429 14875
rect 18463 14841 18475 14875
rect 18417 14835 18475 14841
rect 18984 14804 19012 14980
rect 19426 14940 19432 14952
rect 19387 14912 19432 14940
rect 19426 14900 19432 14912
rect 19484 14900 19490 14952
rect 19536 14940 19564 14980
rect 19702 14968 19708 14980
rect 19760 14968 19766 15020
rect 20346 14968 20352 15020
rect 20404 15008 20410 15020
rect 20625 15011 20683 15017
rect 20625 15008 20637 15011
rect 20404 14980 20637 15008
rect 20404 14968 20410 14980
rect 20625 14977 20637 14980
rect 20671 14977 20683 15011
rect 20625 14971 20683 14977
rect 20806 14940 20812 14952
rect 19536 14912 20812 14940
rect 20806 14900 20812 14912
rect 20864 14900 20870 14952
rect 20441 14875 20499 14881
rect 20441 14872 20453 14875
rect 19076 14844 20453 14872
rect 19076 14813 19104 14844
rect 20441 14841 20453 14844
rect 20487 14841 20499 14875
rect 20441 14835 20499 14841
rect 18340 14776 19012 14804
rect 19061 14807 19119 14813
rect 18049 14767 18107 14773
rect 19061 14773 19073 14807
rect 19107 14773 19119 14807
rect 19518 14804 19524 14816
rect 19479 14776 19524 14804
rect 19061 14767 19119 14773
rect 19518 14764 19524 14776
rect 19576 14764 19582 14816
rect 19978 14764 19984 14816
rect 20036 14804 20042 14816
rect 20073 14807 20131 14813
rect 20073 14804 20085 14807
rect 20036 14776 20085 14804
rect 20036 14764 20042 14776
rect 20073 14773 20085 14776
rect 20119 14773 20131 14807
rect 20530 14804 20536 14816
rect 20491 14776 20536 14804
rect 20073 14767 20131 14773
rect 20530 14764 20536 14776
rect 20588 14764 20594 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 2866 14600 2872 14612
rect 2827 14572 2872 14600
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 3237 14603 3295 14609
rect 3237 14569 3249 14603
rect 3283 14600 3295 14603
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 3283 14572 4077 14600
rect 3283 14569 3295 14572
rect 3237 14563 3295 14569
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 4065 14563 4123 14569
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 4525 14603 4583 14609
rect 4525 14600 4537 14603
rect 4212 14572 4537 14600
rect 4212 14560 4218 14572
rect 4525 14569 4537 14572
rect 4571 14569 4583 14603
rect 5902 14600 5908 14612
rect 4525 14563 4583 14569
rect 4908 14572 5908 14600
rect 2317 14535 2375 14541
rect 2317 14501 2329 14535
rect 2363 14532 2375 14535
rect 2685 14535 2743 14541
rect 2685 14532 2697 14535
rect 2363 14504 2697 14532
rect 2363 14501 2375 14504
rect 2317 14495 2375 14501
rect 2685 14501 2697 14504
rect 2731 14501 2743 14535
rect 2685 14495 2743 14501
rect 3329 14535 3387 14541
rect 3329 14501 3341 14535
rect 3375 14532 3387 14535
rect 4246 14532 4252 14544
rect 3375 14504 4252 14532
rect 3375 14501 3387 14504
rect 3329 14495 3387 14501
rect 4246 14492 4252 14504
rect 4304 14492 4310 14544
rect 4908 14532 4936 14572
rect 5902 14560 5908 14572
rect 5960 14560 5966 14612
rect 6362 14560 6368 14612
rect 6420 14600 6426 14612
rect 7929 14603 7987 14609
rect 7929 14600 7941 14603
rect 6420 14572 7941 14600
rect 6420 14560 6426 14572
rect 7929 14569 7941 14572
rect 7975 14600 7987 14603
rect 8754 14600 8760 14612
rect 7975 14572 8760 14600
rect 7975 14569 7987 14572
rect 7929 14563 7987 14569
rect 8754 14560 8760 14572
rect 8812 14560 8818 14612
rect 9582 14600 9588 14612
rect 8864 14572 9588 14600
rect 4356 14504 4936 14532
rect 5353 14535 5411 14541
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 2225 14467 2283 14473
rect 2225 14464 2237 14467
rect 1443 14436 2237 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2225 14433 2237 14436
rect 2271 14433 2283 14467
rect 3602 14464 3608 14476
rect 2225 14427 2283 14433
rect 2424 14436 3608 14464
rect 2038 14356 2044 14408
rect 2096 14396 2102 14408
rect 2424 14405 2452 14436
rect 3602 14424 3608 14436
rect 3660 14464 3666 14476
rect 4356 14464 4384 14504
rect 5353 14501 5365 14535
rect 5399 14532 5411 14535
rect 5626 14532 5632 14544
rect 5399 14504 5632 14532
rect 5399 14501 5411 14504
rect 5353 14495 5411 14501
rect 5626 14492 5632 14504
rect 5684 14492 5690 14544
rect 6086 14492 6092 14544
rect 6144 14541 6150 14544
rect 6144 14535 6208 14541
rect 6144 14501 6162 14535
rect 6196 14501 6208 14535
rect 6144 14495 6208 14501
rect 6144 14492 6150 14495
rect 6546 14492 6552 14544
rect 6604 14532 6610 14544
rect 8018 14532 8024 14544
rect 6604 14504 8024 14532
rect 6604 14492 6610 14504
rect 8018 14492 8024 14504
rect 8076 14492 8082 14544
rect 3660 14436 4384 14464
rect 4433 14467 4491 14473
rect 3660 14424 3666 14436
rect 4433 14433 4445 14467
rect 4479 14433 4491 14467
rect 4433 14427 4491 14433
rect 5077 14467 5135 14473
rect 5077 14433 5089 14467
rect 5123 14464 5135 14467
rect 7558 14464 7564 14476
rect 5123 14436 7564 14464
rect 5123 14433 5135 14436
rect 5077 14427 5135 14433
rect 2409 14399 2467 14405
rect 2409 14396 2421 14399
rect 2096 14368 2421 14396
rect 2096 14356 2102 14368
rect 2409 14365 2421 14368
rect 2455 14365 2467 14399
rect 3510 14396 3516 14408
rect 3471 14368 3516 14396
rect 2409 14359 2467 14365
rect 3510 14356 3516 14368
rect 3568 14356 3574 14408
rect 1857 14331 1915 14337
rect 1857 14297 1869 14331
rect 1903 14328 1915 14331
rect 4448 14328 4476 14427
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 8864 14464 8892 14572
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 9953 14603 10011 14609
rect 9953 14569 9965 14603
rect 9999 14600 10011 14603
rect 10502 14600 10508 14612
rect 9999 14572 10508 14600
rect 9999 14569 10011 14572
rect 9953 14563 10011 14569
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 10962 14560 10968 14612
rect 11020 14600 11026 14612
rect 12345 14603 12403 14609
rect 12345 14600 12357 14603
rect 11020 14572 12357 14600
rect 11020 14560 11026 14572
rect 12345 14569 12357 14572
rect 12391 14569 12403 14603
rect 12345 14563 12403 14569
rect 13354 14560 13360 14612
rect 13412 14600 13418 14612
rect 16393 14603 16451 14609
rect 16393 14600 16405 14603
rect 13412 14572 16405 14600
rect 13412 14560 13418 14572
rect 16393 14569 16405 14572
rect 16439 14569 16451 14603
rect 16393 14563 16451 14569
rect 16853 14603 16911 14609
rect 16853 14569 16865 14603
rect 16899 14600 16911 14603
rect 18414 14600 18420 14612
rect 16899 14572 18000 14600
rect 18375 14572 18420 14600
rect 16899 14569 16911 14572
rect 16853 14563 16911 14569
rect 9766 14492 9772 14544
rect 9824 14532 9830 14544
rect 10413 14535 10471 14541
rect 10413 14532 10425 14535
rect 9824 14504 10425 14532
rect 9824 14492 9830 14504
rect 10413 14501 10425 14504
rect 10459 14501 10471 14535
rect 10413 14495 10471 14501
rect 10686 14492 10692 14544
rect 10744 14532 10750 14544
rect 12437 14535 12495 14541
rect 12437 14532 12449 14535
rect 10744 14504 12449 14532
rect 10744 14492 10750 14504
rect 12437 14501 12449 14504
rect 12483 14501 12495 14535
rect 12437 14495 12495 14501
rect 14642 14492 14648 14544
rect 14700 14532 14706 14544
rect 15102 14532 15108 14544
rect 14700 14504 15108 14532
rect 14700 14492 14706 14504
rect 15102 14492 15108 14504
rect 15160 14492 15166 14544
rect 15565 14535 15623 14541
rect 15565 14501 15577 14535
rect 15611 14532 15623 14535
rect 16206 14532 16212 14544
rect 15611 14504 16212 14532
rect 15611 14501 15623 14504
rect 15565 14495 15623 14501
rect 16206 14492 16212 14504
rect 16264 14492 16270 14544
rect 17304 14535 17362 14541
rect 17304 14501 17316 14535
rect 17350 14532 17362 14535
rect 17862 14532 17868 14544
rect 17350 14504 17868 14532
rect 17350 14501 17362 14504
rect 17304 14495 17362 14501
rect 17862 14492 17868 14504
rect 17920 14492 17926 14544
rect 17972 14532 18000 14572
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 18598 14560 18604 14612
rect 18656 14600 18662 14612
rect 18693 14603 18751 14609
rect 18693 14600 18705 14603
rect 18656 14572 18705 14600
rect 18656 14560 18662 14572
rect 18693 14569 18705 14572
rect 18739 14569 18751 14603
rect 18693 14563 18751 14569
rect 19705 14603 19763 14609
rect 19705 14569 19717 14603
rect 19751 14600 19763 14603
rect 20530 14600 20536 14612
rect 19751 14572 20536 14600
rect 19751 14569 19763 14572
rect 19705 14563 19763 14569
rect 20530 14560 20536 14572
rect 20588 14560 20594 14612
rect 18782 14532 18788 14544
rect 17972 14504 18788 14532
rect 18782 14492 18788 14504
rect 18840 14492 18846 14544
rect 19242 14492 19248 14544
rect 19300 14492 19306 14544
rect 19610 14492 19616 14544
rect 19668 14532 19674 14544
rect 20165 14535 20223 14541
rect 20165 14532 20177 14535
rect 19668 14504 20177 14532
rect 19668 14492 19674 14504
rect 20165 14501 20177 14504
rect 20211 14501 20223 14535
rect 20165 14495 20223 14501
rect 8036 14436 8892 14464
rect 8941 14467 8999 14473
rect 4709 14399 4767 14405
rect 4709 14365 4721 14399
rect 4755 14396 4767 14399
rect 4798 14396 4804 14408
rect 4755 14368 4804 14396
rect 4755 14365 4767 14368
rect 4709 14359 4767 14365
rect 4798 14356 4804 14368
rect 4856 14356 4862 14408
rect 5905 14399 5963 14405
rect 5905 14365 5917 14399
rect 5951 14365 5963 14399
rect 5905 14359 5963 14365
rect 1903 14300 4476 14328
rect 1903 14297 1915 14300
rect 1857 14291 1915 14297
rect 5074 14288 5080 14340
rect 5132 14328 5138 14340
rect 5920 14328 5948 14359
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 8036 14405 8064 14436
rect 8941 14433 8953 14467
rect 8987 14464 8999 14467
rect 9582 14464 9588 14476
rect 8987 14436 9588 14464
rect 8987 14433 8999 14436
rect 8941 14427 8999 14433
rect 9582 14424 9588 14436
rect 9640 14424 9646 14476
rect 10042 14464 10048 14476
rect 9784 14436 10048 14464
rect 9784 14408 9812 14436
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 10321 14467 10379 14473
rect 10321 14433 10333 14467
rect 10367 14464 10379 14467
rect 11146 14464 11152 14476
rect 10367 14436 11152 14464
rect 10367 14433 10379 14436
rect 10321 14427 10379 14433
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 11330 14464 11336 14476
rect 11256 14436 11336 14464
rect 8021 14399 8079 14405
rect 8021 14396 8033 14399
rect 7432 14368 8033 14396
rect 7432 14356 7438 14368
rect 8021 14365 8033 14368
rect 8067 14365 8079 14399
rect 8021 14359 8079 14365
rect 8110 14356 8116 14408
rect 8168 14396 8174 14408
rect 9033 14399 9091 14405
rect 8168 14368 8213 14396
rect 8168 14356 8174 14368
rect 9033 14365 9045 14399
rect 9079 14365 9091 14399
rect 9033 14359 9091 14365
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14396 9183 14399
rect 9306 14396 9312 14408
rect 9171 14368 9312 14396
rect 9171 14365 9183 14368
rect 9125 14359 9183 14365
rect 5132 14300 5948 14328
rect 5132 14288 5138 14300
rect 2685 14263 2743 14269
rect 2685 14229 2697 14263
rect 2731 14260 2743 14263
rect 3602 14260 3608 14272
rect 2731 14232 3608 14260
rect 2731 14229 2743 14232
rect 2685 14223 2743 14229
rect 3602 14220 3608 14232
rect 3660 14220 3666 14272
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 5442 14260 5448 14272
rect 4120 14232 5448 14260
rect 4120 14220 4126 14232
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 5920 14260 5948 14300
rect 7098 14288 7104 14340
rect 7156 14328 7162 14340
rect 8573 14331 8631 14337
rect 8573 14328 8585 14331
rect 7156 14300 8585 14328
rect 7156 14288 7162 14300
rect 8573 14297 8585 14300
rect 8619 14297 8631 14331
rect 9048 14328 9076 14359
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 9766 14356 9772 14408
rect 9824 14356 9830 14408
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14396 10563 14399
rect 10778 14396 10784 14408
rect 10551 14368 10784 14396
rect 10551 14365 10563 14368
rect 10505 14359 10563 14365
rect 10042 14328 10048 14340
rect 9048 14300 10048 14328
rect 8573 14291 8631 14297
rect 10042 14288 10048 14300
rect 10100 14288 10106 14340
rect 10520 14328 10548 14359
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 11256 14396 11284 14436
rect 11330 14424 11336 14436
rect 11388 14424 11394 14476
rect 13354 14464 13360 14476
rect 13315 14436 13360 14464
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 14366 14464 14372 14476
rect 14327 14436 14372 14464
rect 14366 14424 14372 14436
rect 14424 14424 14430 14476
rect 14461 14467 14519 14473
rect 14461 14433 14473 14467
rect 14507 14464 14519 14467
rect 15286 14464 15292 14476
rect 14507 14436 14679 14464
rect 15247 14436 15292 14464
rect 14507 14433 14519 14436
rect 14461 14427 14519 14433
rect 11422 14396 11428 14408
rect 11112 14368 11284 14396
rect 11383 14368 11428 14396
rect 11112 14356 11118 14368
rect 11422 14356 11428 14368
rect 11480 14356 11486 14408
rect 11514 14356 11520 14408
rect 11572 14396 11578 14408
rect 11572 14368 11617 14396
rect 11572 14356 11578 14368
rect 11882 14356 11888 14408
rect 11940 14396 11946 14408
rect 12529 14399 12587 14405
rect 12529 14396 12541 14399
rect 11940 14368 12541 14396
rect 11940 14356 11946 14368
rect 12529 14365 12541 14368
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 12710 14356 12716 14408
rect 12768 14396 12774 14408
rect 13449 14399 13507 14405
rect 13449 14396 13461 14399
rect 12768 14368 13461 14396
rect 12768 14356 12774 14368
rect 13449 14365 13461 14368
rect 13495 14365 13507 14399
rect 13449 14359 13507 14365
rect 13538 14356 13544 14408
rect 13596 14396 13602 14408
rect 13596 14368 13641 14396
rect 13596 14356 13602 14368
rect 14090 14356 14096 14408
rect 14148 14396 14154 14408
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 14148 14368 14565 14396
rect 14148 14356 14154 14368
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 14651 14396 14679 14436
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 16022 14424 16028 14476
rect 16080 14464 16086 14476
rect 17037 14467 17095 14473
rect 17037 14464 17049 14467
rect 16080 14436 17049 14464
rect 16080 14424 16086 14436
rect 17037 14433 17049 14436
rect 17083 14464 17095 14467
rect 17586 14464 17592 14476
rect 17083 14436 17592 14464
rect 17083 14433 17095 14436
rect 17037 14427 17095 14433
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 18690 14424 18696 14476
rect 18748 14464 18754 14476
rect 19061 14467 19119 14473
rect 19061 14464 19073 14467
rect 18748 14436 19073 14464
rect 18748 14424 18754 14436
rect 19061 14433 19073 14436
rect 19107 14433 19119 14467
rect 19260 14464 19288 14492
rect 20073 14467 20131 14473
rect 20073 14464 20085 14467
rect 19260 14436 20085 14464
rect 19061 14427 19119 14433
rect 20073 14433 20085 14436
rect 20119 14433 20131 14467
rect 20073 14427 20131 14433
rect 16206 14396 16212 14408
rect 14651 14368 16212 14396
rect 14553 14359 14611 14365
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 16482 14396 16488 14408
rect 16443 14368 16488 14396
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14396 16635 14399
rect 16623 14368 16988 14396
rect 16623 14365 16635 14368
rect 16577 14359 16635 14365
rect 10428 14300 10548 14328
rect 6638 14260 6644 14272
rect 5920 14232 6644 14260
rect 6638 14220 6644 14232
rect 6696 14220 6702 14272
rect 7285 14263 7343 14269
rect 7285 14229 7297 14263
rect 7331 14260 7343 14263
rect 7374 14260 7380 14272
rect 7331 14232 7380 14260
rect 7331 14229 7343 14232
rect 7285 14223 7343 14229
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 7466 14220 7472 14272
rect 7524 14260 7530 14272
rect 7561 14263 7619 14269
rect 7561 14260 7573 14263
rect 7524 14232 7573 14260
rect 7524 14220 7530 14232
rect 7561 14229 7573 14232
rect 7607 14229 7619 14263
rect 7561 14223 7619 14229
rect 9122 14220 9128 14272
rect 9180 14260 9186 14272
rect 10428 14260 10456 14300
rect 13170 14288 13176 14340
rect 13228 14328 13234 14340
rect 15930 14328 15936 14340
rect 13228 14300 15936 14328
rect 13228 14288 13234 14300
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 16025 14331 16083 14337
rect 16025 14297 16037 14331
rect 16071 14328 16083 14331
rect 16666 14328 16672 14340
rect 16071 14300 16672 14328
rect 16071 14297 16083 14300
rect 16025 14291 16083 14297
rect 16666 14288 16672 14300
rect 16724 14288 16730 14340
rect 9180 14232 10456 14260
rect 9180 14220 9186 14232
rect 10594 14220 10600 14272
rect 10652 14260 10658 14272
rect 10965 14263 11023 14269
rect 10965 14260 10977 14263
rect 10652 14232 10977 14260
rect 10652 14220 10658 14232
rect 10965 14229 10977 14232
rect 11011 14229 11023 14263
rect 11974 14260 11980 14272
rect 11935 14232 11980 14260
rect 10965 14223 11023 14229
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 12989 14263 13047 14269
rect 12989 14229 13001 14263
rect 13035 14260 13047 14263
rect 13906 14260 13912 14272
rect 13035 14232 13912 14260
rect 13035 14229 13047 14232
rect 12989 14223 13047 14229
rect 13906 14220 13912 14232
rect 13964 14220 13970 14272
rect 14001 14263 14059 14269
rect 14001 14229 14013 14263
rect 14047 14260 14059 14263
rect 16853 14263 16911 14269
rect 16853 14260 16865 14263
rect 14047 14232 16865 14260
rect 14047 14229 14059 14232
rect 14001 14223 14059 14229
rect 16853 14229 16865 14232
rect 16899 14229 16911 14263
rect 16960 14260 16988 14368
rect 18046 14356 18052 14408
rect 18104 14396 18110 14408
rect 19153 14399 19211 14405
rect 19153 14396 19165 14399
rect 18104 14368 19165 14396
rect 18104 14356 18110 14368
rect 19153 14365 19165 14368
rect 19199 14365 19211 14399
rect 19153 14359 19211 14365
rect 19245 14399 19303 14405
rect 19245 14365 19257 14399
rect 19291 14365 19303 14399
rect 19245 14359 19303 14365
rect 18138 14288 18144 14340
rect 18196 14328 18202 14340
rect 18782 14328 18788 14340
rect 18196 14300 18788 14328
rect 18196 14288 18202 14300
rect 18782 14288 18788 14300
rect 18840 14288 18846 14340
rect 17218 14260 17224 14272
rect 16960 14232 17224 14260
rect 16853 14223 16911 14229
rect 17218 14220 17224 14232
rect 17276 14260 17282 14272
rect 17402 14260 17408 14272
rect 17276 14232 17408 14260
rect 17276 14220 17282 14232
rect 17402 14220 17408 14232
rect 17460 14260 17466 14272
rect 19260 14260 19288 14359
rect 19702 14356 19708 14408
rect 19760 14396 19766 14408
rect 20257 14399 20315 14405
rect 20257 14396 20269 14399
rect 19760 14368 20269 14396
rect 19760 14356 19766 14368
rect 20257 14365 20269 14368
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20772 14368 20913 14396
rect 20772 14356 20778 14368
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 17460 14232 19288 14260
rect 17460 14220 17466 14232
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 4154 14056 4160 14068
rect 3436 14028 4160 14056
rect 2866 13988 2872 14000
rect 2424 13960 2872 13988
rect 2424 13929 2452 13960
rect 2866 13948 2872 13960
rect 2924 13988 2930 14000
rect 3326 13988 3332 14000
rect 2924 13960 3332 13988
rect 2924 13948 2930 13960
rect 3326 13948 3332 13960
rect 3384 13948 3390 14000
rect 3436 13929 3464 14028
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 5350 14056 5356 14068
rect 5311 14028 5356 14056
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 5592 14028 5641 14056
rect 5592 14016 5598 14028
rect 5629 14025 5641 14028
rect 5675 14025 5687 14059
rect 5629 14019 5687 14025
rect 6270 14016 6276 14068
rect 6328 14056 6334 14068
rect 6638 14056 6644 14068
rect 6328 14028 6644 14056
rect 6328 14016 6334 14028
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 7190 14016 7196 14068
rect 7248 14056 7254 14068
rect 8110 14056 8116 14068
rect 7248 14028 8116 14056
rect 7248 14016 7254 14028
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 9122 14016 9128 14068
rect 9180 14056 9186 14068
rect 9217 14059 9275 14065
rect 9217 14056 9229 14059
rect 9180 14028 9229 14056
rect 9180 14016 9186 14028
rect 9217 14025 9229 14028
rect 9263 14025 9275 14059
rect 9217 14019 9275 14025
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 9858 14056 9864 14068
rect 9815 14028 9864 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 10137 14059 10195 14065
rect 10137 14025 10149 14059
rect 10183 14056 10195 14059
rect 10410 14056 10416 14068
rect 10183 14028 10416 14056
rect 10183 14025 10195 14028
rect 10137 14019 10195 14025
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 11146 14056 11152 14068
rect 11107 14028 11152 14056
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 14093 14059 14151 14065
rect 14093 14025 14105 14059
rect 14139 14056 14151 14059
rect 14182 14056 14188 14068
rect 14139 14028 14188 14056
rect 14139 14025 14151 14028
rect 14093 14019 14151 14025
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 14737 14059 14795 14065
rect 14737 14025 14749 14059
rect 14783 14056 14795 14059
rect 16758 14056 16764 14068
rect 14783 14028 16620 14056
rect 16719 14028 16764 14056
rect 14783 14025 14795 14028
rect 14737 14019 14795 14025
rect 5368 13988 5396 14016
rect 7208 13988 7236 14016
rect 5368 13960 7420 13988
rect 2409 13923 2467 13929
rect 2409 13889 2421 13923
rect 2455 13889 2467 13923
rect 2409 13883 2467 13889
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13889 2651 13923
rect 2593 13883 2651 13889
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13889 3479 13923
rect 3421 13883 3479 13889
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 3694 13920 3700 13932
rect 3651 13892 3700 13920
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 1670 13852 1676 13864
rect 1443 13824 1676 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 2608 13852 2636 13883
rect 3694 13880 3700 13892
rect 3752 13920 3758 13932
rect 3752 13892 4108 13920
rect 3752 13880 3758 13892
rect 2608 13824 3832 13852
rect 1578 13744 1584 13796
rect 1636 13784 1642 13796
rect 3329 13787 3387 13793
rect 3329 13784 3341 13787
rect 1636 13756 3341 13784
rect 1636 13744 1642 13756
rect 3329 13753 3341 13756
rect 3375 13753 3387 13787
rect 3804 13784 3832 13824
rect 3878 13812 3884 13864
rect 3936 13852 3942 13864
rect 3973 13855 4031 13861
rect 3973 13852 3985 13855
rect 3936 13824 3985 13852
rect 3936 13812 3942 13824
rect 3973 13821 3985 13824
rect 4019 13821 4031 13855
rect 4080 13852 4108 13892
rect 5902 13880 5908 13932
rect 5960 13920 5966 13932
rect 6181 13923 6239 13929
rect 6181 13920 6193 13923
rect 5960 13892 6193 13920
rect 5960 13880 5966 13892
rect 6181 13889 6193 13892
rect 6227 13889 6239 13923
rect 6730 13920 6736 13932
rect 6181 13883 6239 13889
rect 6472 13892 6736 13920
rect 4229 13855 4287 13861
rect 4229 13852 4241 13855
rect 4080 13824 4241 13852
rect 3973 13815 4031 13821
rect 4229 13821 4241 13824
rect 4275 13821 4287 13855
rect 6472 13852 6500 13892
rect 6730 13880 6736 13892
rect 6788 13880 6794 13932
rect 7392 13929 7420 13960
rect 8938 13948 8944 14000
rect 8996 13988 9002 14000
rect 11882 13988 11888 14000
rect 8996 13960 11888 13988
rect 8996 13948 9002 13960
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 16485 13991 16543 13997
rect 16485 13957 16497 13991
rect 16531 13957 16543 13991
rect 16592 13988 16620 14028
rect 16758 14016 16764 14028
rect 16816 14016 16822 14068
rect 18690 14056 18696 14068
rect 18064 14028 18696 14056
rect 18064 13988 18092 14028
rect 18690 14016 18696 14028
rect 18748 14016 18754 14068
rect 19610 14016 19616 14068
rect 19668 14016 19674 14068
rect 19705 14059 19763 14065
rect 19705 14025 19717 14059
rect 19751 14056 19763 14059
rect 20162 14056 20168 14068
rect 19751 14028 20168 14056
rect 19751 14025 19763 14028
rect 19705 14019 19763 14025
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 20898 14056 20904 14068
rect 20859 14028 20904 14056
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 16592 13960 18092 13988
rect 19628 13988 19656 14016
rect 19628 13960 20300 13988
rect 16485 13951 16543 13957
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13889 7435 13923
rect 7377 13883 7435 13889
rect 7466 13880 7472 13932
rect 7524 13880 7530 13932
rect 7650 13880 7656 13932
rect 7708 13920 7714 13932
rect 7837 13923 7895 13929
rect 7837 13920 7849 13923
rect 7708 13892 7849 13920
rect 7708 13880 7714 13892
rect 7837 13889 7849 13892
rect 7883 13889 7895 13923
rect 10594 13920 10600 13932
rect 7837 13883 7895 13889
rect 9508 13892 10456 13920
rect 10555 13892 10600 13920
rect 4229 13815 4287 13821
rect 4356 13824 6500 13852
rect 7285 13855 7343 13861
rect 4356 13784 4384 13824
rect 7285 13821 7297 13855
rect 7331 13852 7343 13855
rect 7484 13852 7512 13880
rect 8110 13861 8116 13864
rect 8104 13852 8116 13861
rect 7331 13824 7512 13852
rect 8071 13824 8116 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 8104 13815 8116 13824
rect 8168 13852 8174 13864
rect 9508 13852 9536 13892
rect 8168 13824 9536 13852
rect 9585 13855 9643 13861
rect 8110 13812 8116 13815
rect 8168 13812 8174 13824
rect 9585 13821 9597 13855
rect 9631 13821 9643 13855
rect 10428 13852 10456 13892
rect 10594 13880 10600 13892
rect 10652 13880 10658 13932
rect 10778 13920 10784 13932
rect 10739 13892 10784 13920
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 11514 13920 11520 13932
rect 10971 13892 11520 13920
rect 10971 13852 10999 13892
rect 11514 13880 11520 13892
rect 11572 13920 11578 13932
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 11572 13892 11713 13920
rect 11572 13880 11578 13892
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 16500 13920 16528 13951
rect 17402 13920 17408 13932
rect 11701 13883 11759 13889
rect 13740 13892 15148 13920
rect 16500 13892 17408 13920
rect 11606 13852 11612 13864
rect 10428 13824 10999 13852
rect 11567 13824 11612 13852
rect 9585 13815 9643 13821
rect 3804 13756 4384 13784
rect 3329 13747 3387 13753
rect 5442 13744 5448 13796
rect 5500 13784 5506 13796
rect 5902 13784 5908 13796
rect 5500 13756 5908 13784
rect 5500 13744 5506 13756
rect 5902 13744 5908 13756
rect 5960 13744 5966 13796
rect 5997 13787 6055 13793
rect 5997 13753 6009 13787
rect 6043 13784 6055 13787
rect 6362 13784 6368 13796
rect 6043 13756 6368 13784
rect 6043 13753 6055 13756
rect 5997 13747 6055 13753
rect 6362 13744 6368 13756
rect 6420 13744 6426 13796
rect 7193 13787 7251 13793
rect 7193 13753 7205 13787
rect 7239 13784 7251 13787
rect 7466 13784 7472 13796
rect 7239 13756 7472 13784
rect 7239 13753 7251 13756
rect 7193 13747 7251 13753
rect 7466 13744 7472 13756
rect 7524 13744 7530 13796
rect 8294 13744 8300 13796
rect 8352 13784 8358 13796
rect 9122 13784 9128 13796
rect 8352 13756 9128 13784
rect 8352 13744 8358 13756
rect 9122 13744 9128 13756
rect 9180 13784 9186 13796
rect 9600 13784 9628 13815
rect 11606 13812 11612 13824
rect 11664 13812 11670 13864
rect 12713 13855 12771 13861
rect 12713 13821 12725 13855
rect 12759 13852 12771 13855
rect 13538 13852 13544 13864
rect 12759 13824 13544 13852
rect 12759 13821 12771 13824
rect 12713 13815 12771 13821
rect 13538 13812 13544 13824
rect 13596 13852 13602 13864
rect 13740 13852 13768 13892
rect 15120 13861 15148 13892
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 20070 13880 20076 13932
rect 20128 13920 20134 13932
rect 20272 13929 20300 13960
rect 20165 13923 20223 13929
rect 20165 13920 20177 13923
rect 20128 13892 20177 13920
rect 20128 13880 20134 13892
rect 20165 13889 20177 13892
rect 20211 13889 20223 13923
rect 20165 13883 20223 13889
rect 20257 13923 20315 13929
rect 20257 13889 20269 13923
rect 20303 13889 20315 13923
rect 20257 13883 20315 13889
rect 15378 13861 15384 13864
rect 13596 13824 13768 13852
rect 14553 13855 14611 13861
rect 13596 13812 13602 13824
rect 14553 13821 14565 13855
rect 14599 13852 14611 13855
rect 15105 13855 15163 13861
rect 14599 13824 15056 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 9180 13756 9628 13784
rect 9180 13744 9186 13756
rect 10134 13744 10140 13796
rect 10192 13784 10198 13796
rect 10505 13787 10563 13793
rect 10505 13784 10517 13787
rect 10192 13756 10517 13784
rect 10192 13744 10198 13756
rect 10505 13753 10517 13756
rect 10551 13784 10563 13787
rect 12980 13787 13038 13793
rect 10551 13756 11652 13784
rect 10551 13753 10563 13756
rect 10505 13747 10563 13753
rect 1946 13716 1952 13728
rect 1907 13688 1952 13716
rect 1946 13676 1952 13688
rect 2004 13676 2010 13728
rect 2038 13676 2044 13728
rect 2096 13716 2102 13728
rect 2317 13719 2375 13725
rect 2317 13716 2329 13719
rect 2096 13688 2329 13716
rect 2096 13676 2102 13688
rect 2317 13685 2329 13688
rect 2363 13685 2375 13719
rect 2958 13716 2964 13728
rect 2919 13688 2964 13716
rect 2317 13679 2375 13685
rect 2958 13676 2964 13688
rect 3016 13676 3022 13728
rect 6089 13719 6147 13725
rect 6089 13685 6101 13719
rect 6135 13716 6147 13719
rect 6825 13719 6883 13725
rect 6825 13716 6837 13719
rect 6135 13688 6837 13716
rect 6135 13685 6147 13688
rect 6089 13679 6147 13685
rect 6825 13685 6837 13688
rect 6871 13685 6883 13719
rect 6825 13679 6883 13685
rect 7098 13676 7104 13728
rect 7156 13716 7162 13728
rect 11054 13716 11060 13728
rect 7156 13688 11060 13716
rect 7156 13676 7162 13688
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 11514 13716 11520 13728
rect 11475 13688 11520 13716
rect 11514 13676 11520 13688
rect 11572 13676 11578 13728
rect 11624 13716 11652 13756
rect 12980 13753 12992 13787
rect 13026 13784 13038 13787
rect 14090 13784 14096 13796
rect 13026 13756 14096 13784
rect 13026 13753 13038 13756
rect 12980 13747 13038 13753
rect 14090 13744 14096 13756
rect 14148 13784 14154 13796
rect 14642 13784 14648 13796
rect 14148 13756 14648 13784
rect 14148 13744 14154 13756
rect 14642 13744 14648 13756
rect 14700 13744 14706 13796
rect 13814 13716 13820 13728
rect 11624 13688 13820 13716
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 15028 13716 15056 13824
rect 15105 13821 15117 13855
rect 15151 13821 15163 13855
rect 15372 13852 15384 13861
rect 15339 13824 15384 13852
rect 15105 13815 15163 13821
rect 15372 13815 15384 13824
rect 15120 13784 15148 13815
rect 15378 13812 15384 13815
rect 15436 13812 15442 13864
rect 17586 13812 17592 13864
rect 17644 13852 17650 13864
rect 17954 13852 17960 13864
rect 17644 13824 17960 13852
rect 17644 13812 17650 13824
rect 17954 13812 17960 13824
rect 18012 13852 18018 13864
rect 18322 13861 18328 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 18012 13824 18061 13852
rect 18012 13812 18018 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18316 13852 18328 13861
rect 18283 13824 18328 13852
rect 18049 13815 18107 13821
rect 18316 13815 18328 13824
rect 18322 13812 18328 13815
rect 18380 13812 18386 13864
rect 20717 13855 20775 13861
rect 20717 13852 20729 13855
rect 18423 13824 20729 13852
rect 15286 13784 15292 13796
rect 15120 13756 15292 13784
rect 15286 13744 15292 13756
rect 15344 13744 15350 13796
rect 15930 13744 15936 13796
rect 15988 13784 15994 13796
rect 18423 13784 18451 13824
rect 20717 13821 20729 13824
rect 20763 13821 20775 13855
rect 20717 13815 20775 13821
rect 15988 13756 18451 13784
rect 15988 13744 15994 13756
rect 18782 13744 18788 13796
rect 18840 13784 18846 13796
rect 20073 13787 20131 13793
rect 20073 13784 20085 13787
rect 18840 13756 20085 13784
rect 18840 13744 18846 13756
rect 20073 13753 20085 13756
rect 20119 13753 20131 13787
rect 20073 13747 20131 13753
rect 16206 13716 16212 13728
rect 15028 13688 16212 13716
rect 16206 13676 16212 13688
rect 16264 13676 16270 13728
rect 16574 13676 16580 13728
rect 16632 13716 16638 13728
rect 17129 13719 17187 13725
rect 17129 13716 17141 13719
rect 16632 13688 17141 13716
rect 16632 13676 16638 13688
rect 17129 13685 17141 13688
rect 17175 13685 17187 13719
rect 17129 13679 17187 13685
rect 17218 13676 17224 13728
rect 17276 13716 17282 13728
rect 17276 13688 17321 13716
rect 17276 13676 17282 13688
rect 17586 13676 17592 13728
rect 17644 13716 17650 13728
rect 19429 13719 19487 13725
rect 19429 13716 19441 13719
rect 17644 13688 19441 13716
rect 17644 13676 17650 13688
rect 19429 13685 19441 13688
rect 19475 13685 19487 13719
rect 19429 13679 19487 13685
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 2038 13472 2044 13524
rect 2096 13512 2102 13524
rect 3418 13512 3424 13524
rect 2096 13484 3424 13512
rect 2096 13472 2102 13484
rect 3418 13472 3424 13484
rect 3476 13472 3482 13524
rect 3694 13512 3700 13524
rect 3655 13484 3700 13512
rect 3694 13472 3700 13484
rect 3752 13472 3758 13524
rect 4154 13512 4160 13524
rect 4115 13484 4160 13512
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 4525 13515 4583 13521
rect 4525 13481 4537 13515
rect 4571 13512 4583 13515
rect 5169 13515 5227 13521
rect 5169 13512 5181 13515
rect 4571 13484 5181 13512
rect 4571 13481 4583 13484
rect 4525 13475 4583 13481
rect 5169 13481 5181 13484
rect 5215 13481 5227 13515
rect 5169 13475 5227 13481
rect 5537 13515 5595 13521
rect 5537 13481 5549 13515
rect 5583 13512 5595 13515
rect 5626 13512 5632 13524
rect 5583 13484 5632 13512
rect 5583 13481 5595 13484
rect 5537 13475 5595 13481
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 6822 13512 6828 13524
rect 6783 13484 6828 13512
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 8202 13512 8208 13524
rect 8163 13484 8208 13512
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10045 13515 10103 13521
rect 10045 13512 10057 13515
rect 10008 13484 10057 13512
rect 10008 13472 10014 13484
rect 10045 13481 10057 13484
rect 10091 13512 10103 13515
rect 10502 13512 10508 13524
rect 10091 13484 10508 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 10686 13512 10692 13524
rect 10647 13484 10692 13512
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 11146 13512 11152 13524
rect 11107 13484 11152 13512
rect 11146 13472 11152 13484
rect 11204 13472 11210 13524
rect 11698 13512 11704 13524
rect 11659 13484 11704 13512
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 11974 13472 11980 13524
rect 12032 13512 12038 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 12032 13484 12081 13512
rect 12032 13472 12038 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 12158 13472 12164 13524
rect 12216 13512 12222 13524
rect 12216 13484 12261 13512
rect 12216 13472 12222 13484
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 15010 13512 15016 13524
rect 13504 13484 15016 13512
rect 13504 13472 13510 13484
rect 15010 13472 15016 13484
rect 15068 13472 15074 13524
rect 15289 13515 15347 13521
rect 15289 13481 15301 13515
rect 15335 13512 15347 13515
rect 15746 13512 15752 13524
rect 15335 13484 15516 13512
rect 15707 13484 15752 13512
rect 15335 13481 15347 13484
rect 15289 13475 15347 13481
rect 2958 13444 2964 13456
rect 1596 13416 2964 13444
rect 1596 13385 1624 13416
rect 2958 13404 2964 13416
rect 3016 13404 3022 13456
rect 6730 13404 6736 13456
rect 6788 13444 6794 13456
rect 7285 13447 7343 13453
rect 7285 13444 7297 13447
rect 6788 13416 7297 13444
rect 6788 13404 6794 13416
rect 7285 13413 7297 13416
rect 7331 13413 7343 13447
rect 7285 13407 7343 13413
rect 7374 13404 7380 13456
rect 7432 13444 7438 13456
rect 7834 13444 7840 13456
rect 7432 13416 7840 13444
rect 7432 13404 7438 13416
rect 7834 13404 7840 13416
rect 7892 13444 7898 13456
rect 7892 13416 8248 13444
rect 7892 13404 7898 13416
rect 1581 13379 1639 13385
rect 1581 13345 1593 13379
rect 1627 13345 1639 13379
rect 1581 13339 1639 13345
rect 2406 13336 2412 13388
rect 2464 13376 2470 13388
rect 2584 13379 2642 13385
rect 2584 13376 2596 13379
rect 2464 13348 2596 13376
rect 2464 13336 2470 13348
rect 2584 13345 2596 13348
rect 2630 13376 2642 13379
rect 4617 13379 4675 13385
rect 2630 13348 4108 13376
rect 2630 13345 2642 13348
rect 2584 13339 2642 13345
rect 4080 13320 4108 13348
rect 4617 13345 4629 13379
rect 4663 13376 4675 13379
rect 5442 13376 5448 13388
rect 4663 13348 5448 13376
rect 4663 13345 4675 13348
rect 4617 13339 4675 13345
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 6089 13379 6147 13385
rect 6089 13345 6101 13379
rect 6135 13345 6147 13379
rect 6089 13339 6147 13345
rect 1857 13311 1915 13317
rect 1857 13277 1869 13311
rect 1903 13277 1915 13311
rect 2314 13308 2320 13320
rect 2275 13280 2320 13308
rect 1857 13271 1915 13277
rect 1872 13172 1900 13271
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4709 13311 4767 13317
rect 4709 13308 4721 13311
rect 4120 13280 4721 13308
rect 4120 13268 4126 13280
rect 4709 13277 4721 13280
rect 4755 13277 4767 13311
rect 5626 13308 5632 13320
rect 5587 13280 5632 13308
rect 4709 13271 4767 13277
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 5776 13280 5821 13308
rect 5776 13268 5782 13280
rect 6104 13240 6132 13339
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 7193 13379 7251 13385
rect 7193 13376 7205 13379
rect 7156 13348 7205 13376
rect 7156 13336 7162 13348
rect 7193 13345 7205 13348
rect 7239 13345 7251 13379
rect 8220 13376 8248 13416
rect 9582 13404 9588 13456
rect 9640 13444 9646 13456
rect 10597 13447 10655 13453
rect 10597 13444 10609 13447
rect 9640 13416 10609 13444
rect 9640 13404 9646 13416
rect 10597 13413 10609 13416
rect 10643 13413 10655 13447
rect 10597 13407 10655 13413
rect 10778 13404 10784 13456
rect 10836 13444 10842 13456
rect 10836 13416 11284 13444
rect 10836 13404 10842 13416
rect 8849 13379 8907 13385
rect 8220 13348 8800 13376
rect 7193 13339 7251 13345
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 6822 13308 6828 13320
rect 6604 13280 6828 13308
rect 6604 13268 6610 13280
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 7374 13308 7380 13320
rect 7335 13280 7380 13308
rect 7374 13268 7380 13280
rect 7432 13268 7438 13320
rect 8294 13308 8300 13320
rect 8255 13280 8300 13308
rect 8294 13268 8300 13280
rect 8352 13268 8358 13320
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13308 8539 13311
rect 8662 13308 8668 13320
rect 8527 13280 8668 13308
rect 8527 13277 8539 13280
rect 8481 13271 8539 13277
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 8772 13308 8800 13348
rect 8849 13345 8861 13379
rect 8895 13376 8907 13379
rect 9122 13376 9128 13388
rect 8895 13348 9128 13376
rect 8895 13345 8907 13348
rect 8849 13339 8907 13345
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 10226 13376 10232 13388
rect 10183 13348 10232 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 10226 13336 10232 13348
rect 10284 13376 10290 13388
rect 10284 13348 10640 13376
rect 10284 13336 10290 13348
rect 10321 13311 10379 13317
rect 10321 13308 10333 13311
rect 8772 13280 10333 13308
rect 10321 13277 10333 13280
rect 10367 13308 10379 13311
rect 10502 13308 10508 13320
rect 10367 13280 10508 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10502 13268 10508 13280
rect 10560 13268 10566 13320
rect 10612 13308 10640 13348
rect 10686 13336 10692 13388
rect 10744 13376 10750 13388
rect 11057 13379 11115 13385
rect 11057 13376 11069 13379
rect 10744 13348 11069 13376
rect 10744 13336 10750 13348
rect 11057 13345 11069 13348
rect 11103 13345 11115 13379
rect 11057 13339 11115 13345
rect 11256 13317 11284 13416
rect 12618 13404 12624 13456
rect 12676 13444 12682 13456
rect 13722 13444 13728 13456
rect 12676 13416 13728 13444
rect 12676 13404 12682 13416
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 15488 13444 15516 13484
rect 15746 13472 15752 13484
rect 15804 13472 15810 13524
rect 16393 13515 16451 13521
rect 16393 13481 16405 13515
rect 16439 13512 16451 13515
rect 16574 13512 16580 13524
rect 16439 13484 16580 13512
rect 16439 13481 16451 13484
rect 16393 13475 16451 13481
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 16761 13515 16819 13521
rect 16761 13481 16773 13515
rect 16807 13512 16819 13515
rect 17405 13515 17463 13521
rect 16807 13484 17356 13512
rect 16807 13481 16819 13484
rect 16761 13475 16819 13481
rect 17218 13444 17224 13456
rect 15488 13416 17224 13444
rect 17218 13404 17224 13416
rect 17276 13404 17282 13456
rect 17328 13444 17356 13484
rect 17405 13481 17417 13515
rect 17451 13512 17463 13515
rect 17678 13512 17684 13524
rect 17451 13484 17684 13512
rect 17451 13481 17463 13484
rect 17405 13475 17463 13481
rect 17678 13472 17684 13484
rect 17736 13472 17742 13524
rect 17773 13515 17831 13521
rect 17773 13481 17785 13515
rect 17819 13512 17831 13515
rect 20714 13512 20720 13524
rect 17819 13484 20720 13512
rect 17819 13481 17831 13484
rect 17773 13475 17831 13481
rect 20714 13472 20720 13484
rect 20772 13472 20778 13524
rect 18046 13444 18052 13456
rect 17328 13416 18052 13444
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 18138 13404 18144 13456
rect 18196 13444 18202 13456
rect 18196 13416 18451 13444
rect 18196 13404 18202 13416
rect 11790 13336 11796 13388
rect 11848 13376 11854 13388
rect 12897 13379 12955 13385
rect 11848 13348 12296 13376
rect 11848 13336 11854 13348
rect 12268 13317 12296 13348
rect 12897 13345 12909 13379
rect 12943 13345 12955 13379
rect 12897 13339 12955 13345
rect 11241 13311 11299 13317
rect 10612 13280 11192 13308
rect 9950 13240 9956 13252
rect 6104 13212 9956 13240
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 11164 13240 11192 13280
rect 11241 13277 11253 13311
rect 11287 13277 11299 13311
rect 11241 13271 11299 13277
rect 12253 13311 12311 13317
rect 12253 13277 12265 13311
rect 12299 13277 12311 13311
rect 12912 13308 12940 13339
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 13538 13376 13544 13388
rect 13044 13348 13089 13376
rect 13499 13348 13544 13376
rect 13044 13336 13050 13348
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 13808 13379 13866 13385
rect 13808 13345 13820 13379
rect 13854 13376 13866 13379
rect 14182 13376 14188 13388
rect 13854 13348 14188 13376
rect 13854 13345 13866 13348
rect 13808 13339 13866 13345
rect 14182 13336 14188 13348
rect 14240 13336 14246 13388
rect 14918 13336 14924 13388
rect 14976 13376 14982 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 14976 13348 15669 13376
rect 14976 13336 14982 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 16574 13376 16580 13388
rect 15657 13339 15715 13345
rect 15764 13348 16580 13376
rect 12912 13280 13584 13308
rect 12253 13271 12311 13277
rect 13556 13252 13584 13280
rect 15194 13268 15200 13320
rect 15252 13308 15258 13320
rect 15764 13308 15792 13348
rect 16574 13336 16580 13348
rect 16632 13376 16638 13388
rect 16853 13379 16911 13385
rect 16853 13376 16865 13379
rect 16632 13348 16865 13376
rect 16632 13336 16638 13348
rect 16853 13345 16865 13348
rect 16899 13345 16911 13379
rect 16853 13339 16911 13345
rect 17034 13336 17040 13388
rect 17092 13376 17098 13388
rect 17865 13379 17923 13385
rect 17865 13376 17877 13379
rect 17092 13348 17877 13376
rect 17092 13336 17098 13348
rect 17865 13345 17877 13348
rect 17911 13376 17923 13379
rect 18423 13376 18451 13416
rect 18598 13404 18604 13456
rect 18656 13444 18662 13456
rect 18656 13416 18701 13444
rect 18656 13404 18662 13416
rect 18782 13404 18788 13456
rect 18840 13444 18846 13456
rect 19337 13447 19395 13453
rect 19337 13444 19349 13447
rect 18840 13416 19349 13444
rect 18840 13404 18846 13416
rect 19337 13413 19349 13416
rect 19383 13444 19395 13447
rect 19797 13447 19855 13453
rect 19797 13444 19809 13447
rect 19383 13416 19809 13444
rect 19383 13413 19395 13416
rect 19337 13407 19395 13413
rect 19797 13413 19809 13416
rect 19843 13413 19855 13447
rect 19797 13407 19855 13413
rect 18693 13379 18751 13385
rect 18693 13376 18705 13379
rect 17911 13348 18081 13376
rect 18423 13348 18705 13376
rect 17911 13345 17923 13348
rect 17865 13339 17923 13345
rect 15930 13308 15936 13320
rect 15252 13280 15792 13308
rect 15843 13280 15936 13308
rect 15252 13268 15258 13280
rect 15930 13268 15936 13280
rect 15988 13308 15994 13320
rect 16758 13308 16764 13320
rect 15988 13280 16764 13308
rect 15988 13268 15994 13280
rect 16758 13268 16764 13280
rect 16816 13308 16822 13320
rect 16945 13311 17003 13317
rect 16945 13308 16957 13311
rect 16816 13280 16957 13308
rect 16816 13268 16822 13280
rect 16945 13277 16957 13280
rect 16991 13277 17003 13311
rect 16945 13271 17003 13277
rect 17402 13268 17408 13320
rect 17460 13308 17466 13320
rect 17957 13311 18015 13317
rect 17957 13308 17969 13311
rect 17460 13280 17969 13308
rect 17460 13268 17466 13280
rect 17957 13277 17969 13280
rect 18003 13277 18015 13311
rect 18053 13308 18081 13348
rect 18693 13345 18705 13348
rect 18739 13345 18751 13379
rect 18693 13339 18751 13345
rect 18877 13311 18935 13317
rect 18053 13280 18552 13308
rect 17957 13271 18015 13277
rect 11790 13240 11796 13252
rect 11164 13212 11796 13240
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 12713 13243 12771 13249
rect 12713 13209 12725 13243
rect 12759 13240 12771 13243
rect 13262 13240 13268 13252
rect 12759 13212 13268 13240
rect 12759 13209 12771 13212
rect 12713 13203 12771 13209
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 13538 13200 13544 13252
rect 13596 13200 13602 13252
rect 18414 13240 18420 13252
rect 14844 13212 18420 13240
rect 5074 13172 5080 13184
rect 1872 13144 5080 13172
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 5902 13132 5908 13184
rect 5960 13172 5966 13184
rect 6273 13175 6331 13181
rect 6273 13172 6285 13175
rect 5960 13144 6285 13172
rect 5960 13132 5966 13144
rect 6273 13141 6285 13144
rect 6319 13141 6331 13175
rect 6730 13172 6736 13184
rect 6691 13144 6736 13172
rect 6273 13135 6331 13141
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 7006 13132 7012 13184
rect 7064 13172 7070 13184
rect 7742 13172 7748 13184
rect 7064 13144 7748 13172
rect 7064 13132 7070 13144
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 7837 13175 7895 13181
rect 7837 13141 7849 13175
rect 7883 13172 7895 13175
rect 8202 13172 8208 13184
rect 7883 13144 8208 13172
rect 7883 13141 7895 13144
rect 7837 13135 7895 13141
rect 8202 13132 8208 13144
rect 8260 13132 8266 13184
rect 8570 13132 8576 13184
rect 8628 13172 8634 13184
rect 9033 13175 9091 13181
rect 9033 13172 9045 13175
rect 8628 13144 9045 13172
rect 8628 13132 8634 13144
rect 9033 13141 9045 13144
rect 9079 13141 9091 13175
rect 9033 13135 9091 13141
rect 9306 13132 9312 13184
rect 9364 13172 9370 13184
rect 9677 13175 9735 13181
rect 9677 13172 9689 13175
rect 9364 13144 9689 13172
rect 9364 13132 9370 13144
rect 9677 13141 9689 13144
rect 9723 13141 9735 13175
rect 9677 13135 9735 13141
rect 10597 13175 10655 13181
rect 10597 13141 10609 13175
rect 10643 13172 10655 13175
rect 12342 13172 12348 13184
rect 10643 13144 12348 13172
rect 10643 13141 10655 13144
rect 10597 13135 10655 13141
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 13173 13175 13231 13181
rect 13173 13141 13185 13175
rect 13219 13172 13231 13175
rect 14844 13172 14872 13212
rect 18414 13200 18420 13212
rect 18472 13200 18478 13252
rect 18524 13240 18552 13280
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 18966 13308 18972 13320
rect 18923 13280 18972 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 18966 13268 18972 13280
rect 19024 13268 19030 13320
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13277 19947 13311
rect 19889 13271 19947 13277
rect 19981 13311 20039 13317
rect 19981 13277 19993 13311
rect 20027 13308 20039 13311
rect 20162 13308 20168 13320
rect 20027 13280 20168 13308
rect 20027 13277 20039 13280
rect 19981 13271 20039 13277
rect 19904 13240 19932 13271
rect 20162 13268 20168 13280
rect 20220 13268 20226 13320
rect 18524 13212 19932 13240
rect 13219 13144 14872 13172
rect 14921 13175 14979 13181
rect 13219 13141 13231 13144
rect 13173 13135 13231 13141
rect 14921 13141 14933 13175
rect 14967 13172 14979 13175
rect 15378 13172 15384 13184
rect 14967 13144 15384 13172
rect 14967 13141 14979 13144
rect 14921 13135 14979 13141
rect 15378 13132 15384 13144
rect 15436 13172 15442 13184
rect 15930 13172 15936 13184
rect 15436 13144 15936 13172
rect 15436 13132 15442 13144
rect 15930 13132 15936 13144
rect 15988 13132 15994 13184
rect 17218 13132 17224 13184
rect 17276 13172 17282 13184
rect 17494 13172 17500 13184
rect 17276 13144 17500 13172
rect 17276 13132 17282 13144
rect 17494 13132 17500 13144
rect 17552 13132 17558 13184
rect 18233 13175 18291 13181
rect 18233 13141 18245 13175
rect 18279 13172 18291 13175
rect 18690 13172 18696 13184
rect 18279 13144 18696 13172
rect 18279 13141 18291 13144
rect 18233 13135 18291 13141
rect 18690 13132 18696 13144
rect 18748 13132 18754 13184
rect 19429 13175 19487 13181
rect 19429 13141 19441 13175
rect 19475 13172 19487 13175
rect 19702 13172 19708 13184
rect 19475 13144 19708 13172
rect 19475 13141 19487 13144
rect 19429 13135 19487 13141
rect 19702 13132 19708 13144
rect 19760 13132 19766 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 4249 12971 4307 12977
rect 4249 12968 4261 12971
rect 2148 12940 4261 12968
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12832 2099 12835
rect 2148 12832 2176 12940
rect 4249 12937 4261 12940
rect 4295 12937 4307 12971
rect 5442 12968 5448 12980
rect 5403 12940 5448 12968
rect 4249 12931 4307 12937
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 6454 12968 6460 12980
rect 6415 12940 6460 12968
rect 6454 12928 6460 12940
rect 6512 12928 6518 12980
rect 7193 12971 7251 12977
rect 7193 12937 7205 12971
rect 7239 12968 7251 12971
rect 7239 12940 8239 12968
rect 7239 12937 7251 12940
rect 7193 12931 7251 12937
rect 3973 12903 4031 12909
rect 3973 12869 3985 12903
rect 4019 12900 4031 12903
rect 4062 12900 4068 12912
rect 4019 12872 4068 12900
rect 4019 12869 4031 12872
rect 3973 12863 4031 12869
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 6638 12900 6644 12912
rect 6380 12872 6644 12900
rect 2087 12804 2176 12832
rect 2225 12835 2283 12841
rect 2087 12801 2099 12804
rect 2041 12795 2099 12801
rect 2225 12801 2237 12835
rect 2271 12832 2283 12835
rect 2406 12832 2412 12844
rect 2271 12804 2412 12832
rect 2271 12801 2283 12804
rect 2225 12795 2283 12801
rect 2406 12792 2412 12804
rect 2464 12792 2470 12844
rect 4801 12835 4859 12841
rect 4801 12832 4813 12835
rect 4540 12804 4813 12832
rect 2314 12724 2320 12776
rect 2372 12764 2378 12776
rect 2590 12764 2596 12776
rect 2372 12736 2596 12764
rect 2372 12724 2378 12736
rect 2590 12724 2596 12736
rect 2648 12764 2654 12776
rect 3878 12764 3884 12776
rect 2648 12736 3884 12764
rect 2648 12724 2654 12736
rect 3878 12724 3884 12736
rect 3936 12764 3942 12776
rect 4430 12764 4436 12776
rect 3936 12736 4436 12764
rect 3936 12724 3942 12736
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 2860 12699 2918 12705
rect 2860 12665 2872 12699
rect 2906 12696 2918 12699
rect 3510 12696 3516 12708
rect 2906 12668 3516 12696
rect 2906 12665 2918 12668
rect 2860 12659 2918 12665
rect 3510 12656 3516 12668
rect 3568 12696 3574 12708
rect 4540 12696 4568 12804
rect 4801 12801 4813 12804
rect 4847 12832 4859 12835
rect 5718 12832 5724 12844
rect 4847 12804 5724 12832
rect 4847 12801 4859 12804
rect 4801 12795 4859 12801
rect 5718 12792 5724 12804
rect 5776 12832 5782 12844
rect 5997 12835 6055 12841
rect 5997 12832 6009 12835
rect 5776 12804 6009 12832
rect 5776 12792 5782 12804
rect 5997 12801 6009 12804
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6380 12776 6408 12872
rect 6638 12860 6644 12872
rect 6696 12860 6702 12912
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 7208 12832 7236 12931
rect 8211 12900 8239 12940
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 9953 12971 10011 12977
rect 9953 12968 9965 12971
rect 8352 12940 9965 12968
rect 8352 12928 8358 12940
rect 9953 12937 9965 12940
rect 9999 12937 10011 12971
rect 14369 12971 14427 12977
rect 9953 12931 10011 12937
rect 10152 12940 14320 12968
rect 8662 12900 8668 12912
rect 8211 12872 8340 12900
rect 8623 12872 8668 12900
rect 6871 12804 7236 12832
rect 8312 12832 8340 12872
rect 8662 12860 8668 12872
rect 8720 12900 8726 12912
rect 8720 12872 9536 12900
rect 8720 12860 8726 12872
rect 9508 12841 9536 12872
rect 9493 12835 9551 12841
rect 8312 12804 9444 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 4709 12767 4767 12773
rect 4709 12733 4721 12767
rect 4755 12764 4767 12767
rect 4890 12764 4896 12776
rect 4755 12736 4896 12764
rect 4755 12733 4767 12736
rect 4709 12727 4767 12733
rect 4890 12724 4896 12736
rect 4948 12724 4954 12776
rect 6362 12724 6368 12776
rect 6420 12724 6426 12776
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 7552 12767 7610 12773
rect 7552 12733 7564 12767
rect 7598 12764 7610 12767
rect 7834 12764 7840 12776
rect 7598 12736 7840 12764
rect 7598 12733 7610 12736
rect 7552 12727 7610 12733
rect 3568 12668 4568 12696
rect 4617 12699 4675 12705
rect 3568 12656 3574 12668
rect 4617 12665 4629 12699
rect 4663 12696 4675 12699
rect 5442 12696 5448 12708
rect 4663 12668 5448 12696
rect 4663 12665 4675 12668
rect 4617 12659 4675 12665
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 5813 12699 5871 12705
rect 5813 12665 5825 12699
rect 5859 12696 5871 12699
rect 6270 12696 6276 12708
rect 5859 12668 6276 12696
rect 5859 12665 5871 12668
rect 5813 12659 5871 12665
rect 6270 12656 6276 12668
rect 6328 12656 6334 12708
rect 1949 12631 2007 12637
rect 1949 12597 1961 12631
rect 1995 12628 2007 12631
rect 2958 12628 2964 12640
rect 1995 12600 2964 12628
rect 1995 12597 2007 12600
rect 1949 12591 2007 12597
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 5902 12588 5908 12640
rect 5960 12628 5966 12640
rect 6656 12628 6684 12727
rect 6822 12656 6828 12708
rect 6880 12696 6886 12708
rect 7300 12696 7328 12727
rect 7834 12724 7840 12736
rect 7892 12724 7898 12776
rect 9306 12764 9312 12776
rect 9267 12736 9312 12764
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 9416 12764 9444 12804
rect 9493 12801 9505 12835
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 10152 12764 10180 12940
rect 11422 12900 11428 12912
rect 10520 12872 11428 12900
rect 10520 12844 10548 12872
rect 11422 12860 11428 12872
rect 11480 12860 11486 12912
rect 14090 12900 14096 12912
rect 14051 12872 14096 12900
rect 14090 12860 14096 12872
rect 14148 12860 14154 12912
rect 14292 12900 14320 12940
rect 14369 12937 14381 12971
rect 14415 12968 14427 12971
rect 14458 12968 14464 12980
rect 14415 12940 14464 12968
rect 14415 12937 14427 12940
rect 14369 12931 14427 12937
rect 14458 12928 14464 12940
rect 14516 12928 14522 12980
rect 16209 12971 16267 12977
rect 16209 12937 16221 12971
rect 16255 12968 16267 12971
rect 16482 12968 16488 12980
rect 16255 12940 16488 12968
rect 16255 12937 16267 12940
rect 16209 12931 16267 12937
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 16666 12928 16672 12980
rect 16724 12968 16730 12980
rect 17865 12971 17923 12977
rect 17865 12968 17877 12971
rect 16724 12940 17877 12968
rect 16724 12928 16730 12940
rect 17865 12937 17877 12940
rect 17911 12937 17923 12971
rect 17865 12931 17923 12937
rect 18782 12928 18788 12980
rect 18840 12968 18846 12980
rect 20438 12968 20444 12980
rect 18840 12940 20444 12968
rect 18840 12928 18846 12940
rect 20438 12928 20444 12940
rect 20496 12928 20502 12980
rect 20640 12940 20944 12968
rect 17678 12900 17684 12912
rect 14292 12872 17684 12900
rect 17678 12860 17684 12872
rect 17736 12860 17742 12912
rect 19150 12900 19156 12912
rect 17788 12872 19156 12900
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10284 12804 10456 12832
rect 10284 12792 10290 12804
rect 10428 12773 10456 12804
rect 10502 12792 10508 12844
rect 10560 12832 10566 12844
rect 10560 12804 10605 12832
rect 10560 12792 10566 12804
rect 10778 12792 10784 12844
rect 10836 12832 10842 12844
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 10836 12804 11529 12832
rect 10836 12792 10842 12804
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 14550 12792 14556 12844
rect 14608 12832 14614 12844
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14608 12804 14933 12832
rect 14608 12792 14614 12804
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 16390 12832 16396 12844
rect 14921 12795 14979 12801
rect 15488 12804 16396 12832
rect 9416 12736 10180 12764
rect 10413 12767 10471 12773
rect 10413 12733 10425 12767
rect 10459 12733 10471 12767
rect 10413 12727 10471 12733
rect 10962 12724 10968 12776
rect 11020 12724 11026 12776
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11425 12767 11483 12773
rect 11425 12764 11437 12767
rect 11204 12736 11437 12764
rect 11204 12724 11210 12736
rect 11425 12733 11437 12736
rect 11471 12764 11483 12767
rect 12066 12764 12072 12776
rect 11471 12736 12072 12764
rect 11471 12733 11483 12736
rect 11425 12727 11483 12733
rect 12066 12724 12072 12736
rect 12124 12724 12130 12776
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12713 12767 12771 12773
rect 12713 12764 12725 12767
rect 12492 12736 12725 12764
rect 12492 12724 12498 12736
rect 12713 12733 12725 12736
rect 12759 12733 12771 12767
rect 12713 12727 12771 12733
rect 13906 12724 13912 12776
rect 13964 12764 13970 12776
rect 14737 12767 14795 12773
rect 14737 12764 14749 12767
rect 13964 12736 14749 12764
rect 13964 12724 13970 12736
rect 14737 12733 14749 12736
rect 14783 12733 14795 12767
rect 14737 12727 14795 12733
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 15488 12764 15516 12804
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 16758 12832 16764 12844
rect 16500 12804 16620 12832
rect 16719 12804 16764 12832
rect 14875 12736 15516 12764
rect 15565 12767 15623 12773
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 15565 12733 15577 12767
rect 15611 12733 15623 12767
rect 15565 12727 15623 12733
rect 9401 12699 9459 12705
rect 6880 12668 9067 12696
rect 6880 12656 6886 12668
rect 7374 12628 7380 12640
rect 5960 12600 6005 12628
rect 6656 12600 7380 12628
rect 5960 12588 5966 12600
rect 7374 12588 7380 12600
rect 7432 12588 7438 12640
rect 8938 12628 8944 12640
rect 8899 12600 8944 12628
rect 8938 12588 8944 12600
rect 8996 12588 9002 12640
rect 9039 12628 9067 12668
rect 9401 12665 9413 12699
rect 9447 12696 9459 12699
rect 9447 12668 10272 12696
rect 9447 12665 9459 12668
rect 9401 12659 9459 12665
rect 10244 12640 10272 12668
rect 9858 12628 9864 12640
rect 9039 12600 9864 12628
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 10226 12588 10232 12640
rect 10284 12588 10290 12640
rect 10321 12631 10379 12637
rect 10321 12597 10333 12631
rect 10367 12628 10379 12631
rect 10410 12628 10416 12640
rect 10367 12600 10416 12628
rect 10367 12597 10379 12600
rect 10321 12591 10379 12597
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 10980 12637 11008 12724
rect 12980 12699 13038 12705
rect 12980 12665 12992 12699
rect 13026 12696 13038 12699
rect 13170 12696 13176 12708
rect 13026 12668 13176 12696
rect 13026 12665 13038 12668
rect 12980 12659 13038 12665
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 15580 12696 15608 12727
rect 15654 12724 15660 12776
rect 15712 12764 15718 12776
rect 15712 12736 15757 12764
rect 15712 12724 15718 12736
rect 16500 12696 16528 12804
rect 16592 12764 16620 12804
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 17788 12832 17816 12872
rect 19150 12860 19156 12872
rect 19208 12860 19214 12912
rect 20162 12900 20168 12912
rect 19260 12872 20168 12900
rect 17144 12804 17816 12832
rect 17865 12835 17923 12841
rect 17144 12764 17172 12804
rect 17865 12801 17877 12835
rect 17911 12832 17923 12835
rect 18785 12835 18843 12841
rect 18785 12832 18797 12835
rect 17911 12804 18797 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 18785 12801 18797 12804
rect 18831 12801 18843 12835
rect 18966 12832 18972 12844
rect 18927 12804 18972 12832
rect 18785 12795 18843 12801
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 16592 12736 17172 12764
rect 17218 12724 17224 12776
rect 17276 12764 17282 12776
rect 17276 12736 17321 12764
rect 17276 12724 17282 12736
rect 18506 12724 18512 12776
rect 18564 12764 18570 12776
rect 18874 12764 18880 12776
rect 18564 12736 18880 12764
rect 18564 12724 18570 12736
rect 18874 12724 18880 12736
rect 18932 12724 18938 12776
rect 14200 12668 15608 12696
rect 15856 12668 16528 12696
rect 16669 12699 16727 12705
rect 10965 12631 11023 12637
rect 10965 12597 10977 12631
rect 11011 12597 11023 12631
rect 11330 12628 11336 12640
rect 11291 12600 11336 12628
rect 10965 12591 11023 12597
rect 11330 12588 11336 12600
rect 11388 12588 11394 12640
rect 13262 12588 13268 12640
rect 13320 12628 13326 12640
rect 14200 12628 14228 12668
rect 13320 12600 14228 12628
rect 13320 12588 13326 12600
rect 15194 12588 15200 12640
rect 15252 12628 15258 12640
rect 15856 12637 15884 12668
rect 16669 12665 16681 12699
rect 16715 12696 16727 12699
rect 17034 12696 17040 12708
rect 16715 12668 17040 12696
rect 16715 12665 16727 12668
rect 16669 12659 16727 12665
rect 17034 12656 17040 12668
rect 17092 12656 17098 12708
rect 17494 12696 17500 12708
rect 17455 12668 17500 12696
rect 17494 12656 17500 12668
rect 17552 12656 17558 12708
rect 17678 12656 17684 12708
rect 17736 12696 17742 12708
rect 19260 12696 19288 12872
rect 20162 12860 20168 12872
rect 20220 12900 20226 12912
rect 20640 12900 20668 12940
rect 20220 12872 20668 12900
rect 20220 12860 20226 12872
rect 20714 12860 20720 12912
rect 20772 12860 20778 12912
rect 19426 12792 19432 12844
rect 19484 12832 19490 12844
rect 19889 12835 19947 12841
rect 19889 12832 19901 12835
rect 19484 12804 19901 12832
rect 19484 12792 19490 12804
rect 19889 12801 19901 12804
rect 19935 12801 19947 12835
rect 19889 12795 19947 12801
rect 19702 12764 19708 12776
rect 19663 12736 19708 12764
rect 19702 12724 19708 12736
rect 19760 12724 19766 12776
rect 19794 12724 19800 12776
rect 19852 12764 19858 12776
rect 20732 12773 20760 12860
rect 20916 12841 20944 12940
rect 20901 12835 20959 12841
rect 20901 12801 20913 12835
rect 20947 12801 20959 12835
rect 20901 12795 20959 12801
rect 20717 12767 20775 12773
rect 19852 12736 19897 12764
rect 19852 12724 19858 12736
rect 20717 12733 20729 12767
rect 20763 12733 20775 12767
rect 20717 12727 20775 12733
rect 17736 12668 19288 12696
rect 17736 12656 17742 12668
rect 15381 12631 15439 12637
rect 15381 12628 15393 12631
rect 15252 12600 15393 12628
rect 15252 12588 15258 12600
rect 15381 12597 15393 12600
rect 15427 12597 15439 12631
rect 15381 12591 15439 12597
rect 15841 12631 15899 12637
rect 15841 12597 15853 12631
rect 15887 12597 15899 12631
rect 15841 12591 15899 12597
rect 16298 12588 16304 12640
rect 16356 12628 16362 12640
rect 16577 12631 16635 12637
rect 16577 12628 16589 12631
rect 16356 12600 16589 12628
rect 16356 12588 16362 12600
rect 16577 12597 16589 12600
rect 16623 12597 16635 12631
rect 16577 12591 16635 12597
rect 18138 12588 18144 12640
rect 18196 12628 18202 12640
rect 18325 12631 18383 12637
rect 18325 12628 18337 12631
rect 18196 12600 18337 12628
rect 18196 12588 18202 12600
rect 18325 12597 18337 12600
rect 18371 12597 18383 12631
rect 18325 12591 18383 12597
rect 18414 12588 18420 12640
rect 18472 12628 18478 12640
rect 18693 12631 18751 12637
rect 18693 12628 18705 12631
rect 18472 12600 18705 12628
rect 18472 12588 18478 12600
rect 18693 12597 18705 12600
rect 18739 12597 18751 12631
rect 18693 12591 18751 12597
rect 19150 12588 19156 12640
rect 19208 12628 19214 12640
rect 19337 12631 19395 12637
rect 19337 12628 19349 12631
rect 19208 12600 19349 12628
rect 19208 12588 19214 12600
rect 19337 12597 19349 12600
rect 19383 12597 19395 12631
rect 19337 12591 19395 12597
rect 20162 12588 20168 12640
rect 20220 12628 20226 12640
rect 20349 12631 20407 12637
rect 20349 12628 20361 12631
rect 20220 12600 20361 12628
rect 20220 12588 20226 12600
rect 20349 12597 20361 12600
rect 20395 12597 20407 12631
rect 20349 12591 20407 12597
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 20864 12600 20909 12628
rect 20864 12588 20870 12600
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 2774 12424 2780 12436
rect 1627 12396 2780 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 2774 12384 2780 12396
rect 2832 12384 2838 12436
rect 2958 12424 2964 12436
rect 2919 12396 2964 12424
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 3970 12384 3976 12436
rect 4028 12424 4034 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 4028 12396 4261 12424
rect 4028 12384 4034 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 4249 12387 4307 12393
rect 5718 12384 5724 12436
rect 5776 12424 5782 12436
rect 6089 12427 6147 12433
rect 6089 12424 6101 12427
rect 5776 12396 6101 12424
rect 5776 12384 5782 12396
rect 6089 12393 6101 12396
rect 6135 12393 6147 12427
rect 6089 12387 6147 12393
rect 6362 12384 6368 12436
rect 6420 12424 6426 12436
rect 6638 12424 6644 12436
rect 6420 12396 6644 12424
rect 6420 12384 6426 12396
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 7377 12427 7435 12433
rect 7377 12393 7389 12427
rect 7423 12424 7435 12427
rect 7558 12424 7564 12436
rect 7423 12396 7564 12424
rect 7423 12393 7435 12396
rect 7377 12387 7435 12393
rect 7558 12384 7564 12396
rect 7616 12384 7622 12436
rect 8205 12427 8263 12433
rect 7668 12396 8064 12424
rect 1486 12316 1492 12368
rect 1544 12356 1550 12368
rect 7668 12356 7696 12396
rect 1544 12328 7696 12356
rect 7745 12359 7803 12365
rect 1544 12316 1550 12328
rect 7745 12325 7757 12359
rect 7791 12356 7803 12359
rect 7926 12356 7932 12368
rect 7791 12328 7932 12356
rect 7791 12325 7803 12328
rect 7745 12319 7803 12325
rect 7926 12316 7932 12328
rect 7984 12316 7990 12368
rect 8036 12356 8064 12396
rect 8205 12393 8217 12427
rect 8251 12424 8263 12427
rect 8849 12427 8907 12433
rect 8849 12424 8861 12427
rect 8251 12396 8861 12424
rect 8251 12393 8263 12396
rect 8205 12387 8263 12393
rect 8849 12393 8861 12396
rect 8895 12393 8907 12427
rect 8849 12387 8907 12393
rect 10226 12384 10232 12436
rect 10284 12424 10290 12436
rect 11517 12427 11575 12433
rect 11517 12424 11529 12427
rect 10284 12396 11529 12424
rect 10284 12384 10290 12396
rect 11517 12393 11529 12396
rect 11563 12393 11575 12427
rect 11882 12424 11888 12436
rect 11843 12396 11888 12424
rect 11517 12387 11575 12393
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 11977 12427 12035 12433
rect 11977 12393 11989 12427
rect 12023 12424 12035 12427
rect 12158 12424 12164 12436
rect 12023 12396 12164 12424
rect 12023 12393 12035 12396
rect 11977 12387 12035 12393
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 12710 12424 12716 12436
rect 12671 12396 12716 12424
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 13081 12427 13139 12433
rect 13081 12393 13093 12427
rect 13127 12424 13139 12427
rect 13262 12424 13268 12436
rect 13127 12396 13268 12424
rect 13127 12393 13139 12396
rect 13081 12387 13139 12393
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 13354 12384 13360 12436
rect 13412 12424 13418 12436
rect 13725 12427 13783 12433
rect 13725 12424 13737 12427
rect 13412 12396 13737 12424
rect 13412 12384 13418 12396
rect 13725 12393 13737 12396
rect 13771 12393 13783 12427
rect 13725 12387 13783 12393
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 15654 12424 15660 12436
rect 15528 12396 15660 12424
rect 15528 12384 15534 12396
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 16574 12424 16580 12436
rect 16040 12396 16580 12424
rect 8757 12359 8815 12365
rect 8757 12356 8769 12359
rect 8036 12328 8769 12356
rect 8757 12325 8769 12328
rect 8803 12325 8815 12359
rect 15841 12359 15899 12365
rect 15841 12356 15853 12359
rect 8757 12319 8815 12325
rect 8864 12328 15853 12356
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1762 12288 1768 12300
rect 1443 12260 1768 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1762 12248 1768 12260
rect 1820 12248 1826 12300
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12288 2375 12291
rect 2958 12288 2964 12300
rect 2363 12260 2964 12288
rect 2363 12257 2375 12260
rect 2317 12251 2375 12257
rect 2958 12248 2964 12260
rect 3016 12248 3022 12300
rect 3326 12288 3332 12300
rect 3287 12260 3332 12288
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 3881 12291 3939 12297
rect 3881 12257 3893 12291
rect 3927 12288 3939 12291
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 3927 12260 4077 12288
rect 3927 12257 3939 12260
rect 3881 12251 3939 12257
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 4065 12251 4123 12257
rect 4430 12248 4436 12300
rect 4488 12288 4494 12300
rect 4982 12297 4988 12300
rect 4709 12291 4767 12297
rect 4709 12288 4721 12291
rect 4488 12260 4721 12288
rect 4488 12248 4494 12260
rect 4709 12257 4721 12260
rect 4755 12257 4767 12291
rect 4976 12288 4988 12297
rect 4943 12260 4988 12288
rect 4709 12251 4767 12257
rect 4976 12251 4988 12260
rect 4982 12248 4988 12251
rect 5040 12248 5046 12300
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12288 6791 12291
rect 7650 12288 7656 12300
rect 6779 12260 7656 12288
rect 6779 12257 6791 12260
rect 6733 12251 6791 12257
rect 7650 12248 7656 12260
rect 7708 12248 7714 12300
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 8864 12288 8892 12328
rect 15841 12325 15853 12328
rect 15887 12325 15899 12359
rect 15841 12319 15899 12325
rect 9858 12288 9864 12300
rect 8628 12260 8892 12288
rect 9819 12260 9864 12288
rect 8628 12248 8634 12260
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 9950 12248 9956 12300
rect 10008 12288 10014 12300
rect 10117 12291 10175 12297
rect 10117 12288 10129 12291
rect 10008 12260 10129 12288
rect 10008 12248 10014 12260
rect 10117 12257 10129 12260
rect 10163 12288 10175 12291
rect 10870 12288 10876 12300
rect 10163 12260 10876 12288
rect 10163 12257 10175 12260
rect 10117 12251 10175 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 13998 12288 14004 12300
rect 13280 12260 14004 12288
rect 1946 12180 1952 12232
rect 2004 12220 2010 12232
rect 2130 12220 2136 12232
rect 2004 12192 2136 12220
rect 2004 12180 2010 12192
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12220 2651 12223
rect 2774 12220 2780 12232
rect 2639 12192 2780 12220
rect 2639 12189 2651 12192
rect 2593 12183 2651 12189
rect 2424 12152 2452 12183
rect 2774 12180 2780 12192
rect 2832 12180 2838 12232
rect 3418 12220 3424 12232
rect 3379 12192 3424 12220
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3510 12180 3516 12232
rect 3568 12220 3574 12232
rect 3568 12192 3613 12220
rect 3568 12180 3574 12192
rect 6178 12180 6184 12232
rect 6236 12220 6242 12232
rect 6822 12220 6828 12232
rect 6236 12192 6828 12220
rect 6236 12180 6242 12192
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 3234 12152 3240 12164
rect 2424 12124 3240 12152
rect 3234 12112 3240 12124
rect 3292 12112 3298 12164
rect 5902 12112 5908 12164
rect 5960 12152 5966 12164
rect 6365 12155 6423 12161
rect 6365 12152 6377 12155
rect 5960 12124 6377 12152
rect 5960 12112 5966 12124
rect 6365 12121 6377 12124
rect 6411 12121 6423 12155
rect 6365 12115 6423 12121
rect 6546 12112 6552 12164
rect 6604 12152 6610 12164
rect 6932 12152 6960 12183
rect 7834 12180 7840 12232
rect 7892 12220 7898 12232
rect 8021 12223 8079 12229
rect 7892 12192 7937 12220
rect 7892 12180 7898 12192
rect 8021 12189 8033 12223
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 8941 12223 8999 12229
rect 8941 12189 8953 12223
rect 8987 12189 8999 12223
rect 11330 12220 11336 12232
rect 11291 12192 11336 12220
rect 8941 12183 8999 12189
rect 6604 12124 6960 12152
rect 6604 12112 6610 12124
rect 1949 12087 2007 12093
rect 1949 12053 1961 12087
rect 1995 12084 2007 12087
rect 2130 12084 2136 12096
rect 1995 12056 2136 12084
rect 1995 12053 2007 12056
rect 1949 12047 2007 12053
rect 2130 12044 2136 12056
rect 2188 12044 2194 12096
rect 3881 12087 3939 12093
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 6454 12084 6460 12096
rect 3927 12056 6460 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 8036 12084 8064 12183
rect 8110 12112 8116 12164
rect 8168 12152 8174 12164
rect 8205 12155 8263 12161
rect 8205 12152 8217 12155
rect 8168 12124 8217 12152
rect 8168 12112 8174 12124
rect 8205 12121 8217 12124
rect 8251 12121 8263 12155
rect 8205 12115 8263 12121
rect 8662 12112 8668 12164
rect 8720 12152 8726 12164
rect 8956 12152 8984 12183
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 11422 12180 11428 12232
rect 11480 12220 11486 12232
rect 12069 12223 12127 12229
rect 12069 12220 12081 12223
rect 11480 12192 12081 12220
rect 11480 12180 11486 12192
rect 12069 12189 12081 12192
rect 12115 12189 12127 12223
rect 12069 12183 12127 12189
rect 12526 12180 12532 12232
rect 12584 12220 12590 12232
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 12584 12192 13185 12220
rect 12584 12180 12590 12192
rect 13173 12189 13185 12192
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 8720 12124 9628 12152
rect 8720 12112 8726 12124
rect 9600 12096 9628 12124
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 9858 12152 9864 12164
rect 9732 12124 9864 12152
rect 9732 12112 9738 12124
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 10870 12112 10876 12164
rect 10928 12152 10934 12164
rect 11241 12155 11299 12161
rect 11241 12152 11253 12155
rect 10928 12124 11253 12152
rect 10928 12112 10934 12124
rect 11241 12121 11253 12124
rect 11287 12152 11299 12155
rect 13280 12152 13308 12260
rect 13998 12248 14004 12260
rect 14056 12248 14062 12300
rect 14093 12291 14151 12297
rect 14093 12257 14105 12291
rect 14139 12288 14151 12291
rect 14737 12291 14795 12297
rect 14737 12288 14749 12291
rect 14139 12260 14749 12288
rect 14139 12257 14151 12260
rect 14093 12251 14151 12257
rect 14737 12257 14749 12260
rect 14783 12257 14795 12291
rect 14737 12251 14795 12257
rect 13354 12180 13360 12232
rect 13412 12220 13418 12232
rect 13412 12192 13457 12220
rect 13412 12180 13418 12192
rect 13722 12180 13728 12232
rect 13780 12220 13786 12232
rect 14185 12223 14243 12229
rect 14185 12220 14197 12223
rect 13780 12192 14197 12220
rect 13780 12180 13786 12192
rect 14185 12189 14197 12192
rect 14231 12189 14243 12223
rect 14185 12183 14243 12189
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 11287 12124 13308 12152
rect 13372 12152 13400 12180
rect 14292 12152 14320 12183
rect 14458 12180 14464 12232
rect 14516 12220 14522 12232
rect 16040 12229 16068 12396
rect 16574 12384 16580 12396
rect 16632 12424 16638 12436
rect 17586 12424 17592 12436
rect 16632 12396 17592 12424
rect 16632 12384 16638 12396
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 17865 12427 17923 12433
rect 17865 12393 17877 12427
rect 17911 12393 17923 12427
rect 17865 12387 17923 12393
rect 16752 12359 16810 12365
rect 16752 12325 16764 12359
rect 16798 12356 16810 12359
rect 17218 12356 17224 12368
rect 16798 12328 17224 12356
rect 16798 12325 16810 12328
rect 16752 12319 16810 12325
rect 17218 12316 17224 12328
rect 17276 12316 17282 12368
rect 17880 12356 17908 12387
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19610 12424 19616 12436
rect 19392 12396 19616 12424
rect 19392 12384 19398 12396
rect 19610 12384 19616 12396
rect 19668 12384 19674 12436
rect 19797 12427 19855 12433
rect 19797 12393 19809 12427
rect 19843 12424 19855 12427
rect 19886 12424 19892 12436
rect 19843 12396 19892 12424
rect 19843 12393 19855 12396
rect 19797 12387 19855 12393
rect 19886 12384 19892 12396
rect 19944 12384 19950 12436
rect 20070 12384 20076 12436
rect 20128 12424 20134 12436
rect 20165 12427 20223 12433
rect 20165 12424 20177 12427
rect 20128 12396 20177 12424
rect 20128 12384 20134 12396
rect 20165 12393 20177 12396
rect 20211 12393 20223 12427
rect 20165 12387 20223 12393
rect 20901 12427 20959 12433
rect 20901 12393 20913 12427
rect 20947 12424 20959 12427
rect 21450 12424 21456 12436
rect 20947 12396 21456 12424
rect 20947 12393 20959 12396
rect 20901 12387 20959 12393
rect 21450 12384 21456 12396
rect 21508 12384 21514 12436
rect 18408 12359 18466 12365
rect 18408 12356 18420 12359
rect 17880 12328 18420 12356
rect 18408 12325 18420 12328
rect 18454 12356 18466 12359
rect 18506 12356 18512 12368
rect 18454 12328 18512 12356
rect 18454 12325 18466 12328
rect 18408 12319 18466 12325
rect 18506 12316 18512 12328
rect 18564 12356 18570 12368
rect 18782 12356 18788 12368
rect 18564 12328 18788 12356
rect 18564 12316 18570 12328
rect 18782 12316 18788 12328
rect 18840 12316 18846 12368
rect 19058 12316 19064 12368
rect 19116 12356 19122 12368
rect 19242 12356 19248 12368
rect 19116 12328 19248 12356
rect 19116 12316 19122 12328
rect 19242 12316 19248 12328
rect 19300 12316 19306 12368
rect 17957 12291 18015 12297
rect 16408 12260 17540 12288
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 14516 12192 15945 12220
rect 14516 12180 14522 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 13372 12124 14320 12152
rect 15473 12155 15531 12161
rect 11287 12121 11299 12124
rect 11241 12115 11299 12121
rect 15473 12121 15485 12155
rect 15519 12152 15531 12155
rect 15838 12152 15844 12164
rect 15519 12124 15844 12152
rect 15519 12121 15531 12124
rect 15473 12115 15531 12121
rect 15838 12112 15844 12124
rect 15896 12112 15902 12164
rect 15948 12152 15976 12183
rect 16408 12152 16436 12260
rect 16485 12223 16543 12229
rect 16485 12189 16497 12223
rect 16531 12189 16543 12223
rect 17512 12220 17540 12260
rect 17957 12257 17969 12291
rect 18003 12288 18015 12291
rect 18046 12288 18052 12300
rect 18003 12260 18052 12288
rect 18003 12257 18015 12260
rect 17957 12251 18015 12257
rect 18046 12248 18052 12260
rect 18104 12288 18110 12300
rect 18141 12291 18199 12297
rect 18141 12288 18153 12291
rect 18104 12260 18153 12288
rect 18104 12248 18110 12260
rect 18141 12257 18153 12260
rect 18187 12257 18199 12291
rect 20438 12288 20444 12300
rect 18141 12251 18199 12257
rect 18248 12260 20444 12288
rect 18248 12220 18276 12260
rect 20438 12248 20444 12260
rect 20496 12248 20502 12300
rect 17512 12192 18276 12220
rect 16485 12183 16543 12189
rect 15948 12124 16436 12152
rect 7156 12056 8064 12084
rect 8389 12087 8447 12093
rect 7156 12044 7162 12056
rect 8389 12053 8401 12087
rect 8435 12084 8447 12087
rect 9214 12084 9220 12096
rect 8435 12056 9220 12084
rect 8435 12053 8447 12056
rect 8389 12047 8447 12053
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 9582 12044 9588 12096
rect 9640 12044 9646 12096
rect 10226 12044 10232 12096
rect 10284 12084 10290 12096
rect 11333 12087 11391 12093
rect 11333 12084 11345 12087
rect 10284 12056 11345 12084
rect 10284 12044 10290 12056
rect 11333 12053 11345 12056
rect 11379 12053 11391 12087
rect 11333 12047 11391 12053
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 14734 12084 14740 12096
rect 13228 12056 14740 12084
rect 13228 12044 13234 12056
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 15194 12044 15200 12096
rect 15252 12084 15258 12096
rect 16390 12084 16396 12096
rect 15252 12056 16396 12084
rect 15252 12044 15258 12056
rect 16390 12044 16396 12056
rect 16448 12084 16454 12096
rect 16500 12084 16528 12183
rect 19794 12180 19800 12232
rect 19852 12220 19858 12232
rect 20257 12223 20315 12229
rect 20257 12220 20269 12223
rect 19852 12192 20269 12220
rect 19852 12180 19858 12192
rect 20257 12189 20269 12192
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 20349 12223 20407 12229
rect 20349 12189 20361 12223
rect 20395 12189 20407 12223
rect 20349 12183 20407 12189
rect 20364 12152 20392 12183
rect 19536 12124 20392 12152
rect 17957 12087 18015 12093
rect 17957 12084 17969 12087
rect 16448 12056 17969 12084
rect 16448 12044 16454 12056
rect 17957 12053 17969 12056
rect 18003 12053 18015 12087
rect 17957 12047 18015 12053
rect 18874 12044 18880 12096
rect 18932 12084 18938 12096
rect 19536 12093 19564 12124
rect 19521 12087 19579 12093
rect 19521 12084 19533 12087
rect 18932 12056 19533 12084
rect 18932 12044 18938 12056
rect 19521 12053 19533 12056
rect 19567 12053 19579 12087
rect 19521 12047 19579 12053
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 4985 11883 5043 11889
rect 4985 11880 4997 11883
rect 4632 11852 4997 11880
rect 4632 11824 4660 11852
rect 4985 11849 4997 11852
rect 5031 11849 5043 11883
rect 4985 11843 5043 11849
rect 5537 11883 5595 11889
rect 5537 11849 5549 11883
rect 5583 11880 5595 11883
rect 5626 11880 5632 11892
rect 5583 11852 5632 11880
rect 5583 11849 5595 11852
rect 5537 11843 5595 11849
rect 5626 11840 5632 11852
rect 5684 11840 5690 11892
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 6825 11883 6883 11889
rect 6825 11880 6837 11883
rect 6328 11852 6837 11880
rect 6328 11840 6334 11852
rect 6825 11849 6837 11852
rect 6871 11849 6883 11883
rect 7834 11880 7840 11892
rect 7795 11852 7840 11880
rect 6825 11843 6883 11849
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 7926 11840 7932 11892
rect 7984 11880 7990 11892
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 7984 11852 8861 11880
rect 7984 11840 7990 11852
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 8849 11843 8907 11849
rect 8956 11852 9444 11880
rect 4614 11772 4620 11824
rect 4672 11772 4678 11824
rect 4709 11815 4767 11821
rect 4709 11781 4721 11815
rect 4755 11812 4767 11815
rect 4890 11812 4896 11824
rect 4755 11784 4896 11812
rect 4755 11781 4767 11784
rect 4709 11775 4767 11781
rect 4890 11772 4896 11784
rect 4948 11812 4954 11824
rect 6546 11812 6552 11824
rect 4948 11784 6552 11812
rect 4948 11772 4954 11784
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 3234 11744 3240 11756
rect 2915 11716 3240 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 3234 11704 3240 11716
rect 3292 11744 3298 11756
rect 6104 11753 6132 11784
rect 6546 11772 6552 11784
rect 6604 11772 6610 11824
rect 7742 11772 7748 11824
rect 7800 11812 7806 11824
rect 8662 11812 8668 11824
rect 7800 11784 8668 11812
rect 7800 11772 7806 11784
rect 8662 11772 8668 11784
rect 8720 11772 8726 11824
rect 6089 11747 6147 11753
rect 3292 11716 3464 11744
rect 3292 11704 3298 11716
rect 1489 11679 1547 11685
rect 1489 11645 1501 11679
rect 1535 11676 1547 11679
rect 1535 11648 2268 11676
rect 1535 11645 1547 11648
rect 1489 11639 1547 11645
rect 1394 11568 1400 11620
rect 1452 11608 1458 11620
rect 1765 11611 1823 11617
rect 1765 11608 1777 11611
rect 1452 11580 1777 11608
rect 1452 11568 1458 11580
rect 1765 11577 1777 11580
rect 1811 11577 1823 11611
rect 1765 11571 1823 11577
rect 2240 11549 2268 11648
rect 2590 11636 2596 11688
rect 2648 11676 2654 11688
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 2648 11648 3341 11676
rect 2648 11636 2654 11648
rect 3329 11645 3341 11648
rect 3375 11645 3387 11679
rect 3436 11676 3464 11716
rect 6089 11713 6101 11747
rect 6135 11713 6147 11747
rect 6564 11744 6592 11772
rect 7377 11747 7435 11753
rect 7377 11744 7389 11747
rect 6564 11716 7389 11744
rect 6089 11707 6147 11713
rect 7377 11713 7389 11716
rect 7423 11713 7435 11747
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 7377 11707 7435 11713
rect 8036 11716 8493 11744
rect 3585 11679 3643 11685
rect 3585 11676 3597 11679
rect 3436 11648 3597 11676
rect 3329 11639 3387 11645
rect 3585 11645 3597 11648
rect 3631 11645 3643 11679
rect 3585 11639 3643 11645
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11645 4859 11679
rect 4801 11639 4859 11645
rect 4246 11568 4252 11620
rect 4304 11608 4310 11620
rect 4614 11608 4620 11620
rect 4304 11580 4620 11608
rect 4304 11568 4310 11580
rect 4614 11568 4620 11580
rect 4672 11568 4678 11620
rect 2225 11543 2283 11549
rect 2225 11509 2237 11543
rect 2271 11509 2283 11543
rect 2225 11503 2283 11509
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 2593 11543 2651 11549
rect 2593 11540 2605 11543
rect 2372 11512 2605 11540
rect 2372 11500 2378 11512
rect 2593 11509 2605 11512
rect 2639 11509 2651 11543
rect 2593 11503 2651 11509
rect 2685 11543 2743 11549
rect 2685 11509 2697 11543
rect 2731 11540 2743 11543
rect 4062 11540 4068 11552
rect 2731 11512 4068 11540
rect 2731 11509 2743 11512
rect 2685 11503 2743 11509
rect 4062 11500 4068 11512
rect 4120 11500 4126 11552
rect 4816 11540 4844 11639
rect 4982 11636 4988 11688
rect 5040 11676 5046 11688
rect 5445 11679 5503 11685
rect 5445 11676 5457 11679
rect 5040 11648 5457 11676
rect 5040 11636 5046 11648
rect 5445 11645 5457 11648
rect 5491 11676 5503 11679
rect 5902 11676 5908 11688
rect 5491 11648 5908 11676
rect 5491 11645 5503 11648
rect 5445 11639 5503 11645
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 6730 11636 6736 11688
rect 6788 11676 6794 11688
rect 8036 11676 8064 11716
rect 8481 11713 8493 11716
rect 8527 11744 8539 11747
rect 8754 11744 8760 11756
rect 8527 11716 8760 11744
rect 8527 11713 8539 11716
rect 8481 11707 8539 11713
rect 8754 11704 8760 11716
rect 8812 11744 8818 11756
rect 8956 11744 8984 11852
rect 9214 11772 9220 11824
rect 9272 11772 9278 11824
rect 8812 11716 8984 11744
rect 8812 11704 8818 11716
rect 8202 11676 8208 11688
rect 6788 11648 8064 11676
rect 8163 11648 8208 11676
rect 6788 11636 6794 11648
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11676 8355 11679
rect 8938 11676 8944 11688
rect 8343 11648 8944 11676
rect 8343 11645 8355 11648
rect 8297 11639 8355 11645
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 9232 11685 9260 11772
rect 9416 11753 9444 11852
rect 9582 11840 9588 11892
rect 9640 11840 9646 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 12158 11880 12164 11892
rect 9732 11852 12164 11880
rect 9732 11840 9738 11852
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 14093 11883 14151 11889
rect 14093 11880 14105 11883
rect 13596 11852 14105 11880
rect 13596 11840 13602 11852
rect 14093 11849 14105 11852
rect 14139 11849 14151 11883
rect 14093 11843 14151 11849
rect 14734 11840 14740 11892
rect 14792 11880 14798 11892
rect 15749 11883 15807 11889
rect 15749 11880 15761 11883
rect 14792 11852 15761 11880
rect 14792 11840 14798 11852
rect 15749 11849 15761 11852
rect 15795 11880 15807 11883
rect 16022 11880 16028 11892
rect 15795 11852 16028 11880
rect 15795 11849 15807 11852
rect 15749 11843 15807 11849
rect 16022 11840 16028 11852
rect 16080 11840 16086 11892
rect 16206 11840 16212 11892
rect 16264 11880 16270 11892
rect 16264 11852 18368 11880
rect 16264 11840 16270 11852
rect 9600 11812 9628 11840
rect 9600 11784 10272 11812
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11713 9459 11747
rect 9401 11707 9459 11713
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 9950 11744 9956 11756
rect 9640 11716 9956 11744
rect 9640 11704 9646 11716
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 10244 11753 10272 11784
rect 11882 11772 11888 11824
rect 11940 11812 11946 11824
rect 11977 11815 12035 11821
rect 11977 11812 11989 11815
rect 11940 11784 11989 11812
rect 11940 11772 11946 11784
rect 11977 11781 11989 11784
rect 12023 11781 12035 11815
rect 11977 11775 12035 11781
rect 13817 11815 13875 11821
rect 13817 11781 13829 11815
rect 13863 11812 13875 11815
rect 14366 11812 14372 11824
rect 13863 11784 14372 11812
rect 13863 11781 13875 11784
rect 13817 11775 13875 11781
rect 14366 11772 14372 11784
rect 14424 11772 14430 11824
rect 17770 11772 17776 11824
rect 17828 11772 17834 11824
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 11790 11704 11796 11756
rect 11848 11744 11854 11756
rect 11848 11716 12572 11744
rect 11848 11704 11854 11716
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11645 9275 11679
rect 9217 11639 9275 11645
rect 9490 11636 9496 11688
rect 9548 11676 9554 11688
rect 10045 11679 10103 11685
rect 10045 11676 10057 11679
rect 9548 11648 10057 11676
rect 9548 11636 9554 11648
rect 10045 11645 10057 11648
rect 10091 11645 10103 11679
rect 10045 11639 10103 11645
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11676 10655 11679
rect 12434 11676 12440 11688
rect 10643 11648 12440 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 12434 11636 12440 11648
rect 12492 11636 12498 11688
rect 12544 11676 12572 11716
rect 15562 11704 15568 11756
rect 15620 11744 15626 11756
rect 16206 11744 16212 11756
rect 15620 11716 16212 11744
rect 15620 11704 15626 11716
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 17310 11704 17316 11756
rect 17368 11744 17374 11756
rect 17788 11744 17816 11772
rect 18340 11753 18368 11852
rect 18598 11840 18604 11892
rect 18656 11880 18662 11892
rect 18785 11883 18843 11889
rect 18785 11880 18797 11883
rect 18656 11852 18797 11880
rect 18656 11840 18662 11852
rect 18785 11849 18797 11852
rect 18831 11849 18843 11883
rect 20990 11880 20996 11892
rect 20951 11852 20996 11880
rect 18785 11843 18843 11849
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 19242 11772 19248 11824
rect 19300 11812 19306 11824
rect 21082 11812 21088 11824
rect 19300 11784 21088 11812
rect 19300 11772 19306 11784
rect 21082 11772 21088 11784
rect 21140 11772 21146 11824
rect 18325 11747 18383 11753
rect 17368 11716 18184 11744
rect 17368 11704 17374 11716
rect 14182 11676 14188 11688
rect 12544 11648 14188 11676
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 14277 11679 14335 11685
rect 14277 11645 14289 11679
rect 14323 11645 14335 11679
rect 14277 11639 14335 11645
rect 14369 11679 14427 11685
rect 14369 11645 14381 11679
rect 14415 11676 14427 11679
rect 15194 11676 15200 11688
rect 14415 11648 15200 11676
rect 14415 11645 14427 11648
rect 14369 11639 14427 11645
rect 5997 11611 6055 11617
rect 5997 11577 6009 11611
rect 6043 11608 6055 11611
rect 6086 11608 6092 11620
rect 6043 11580 6092 11608
rect 6043 11577 6055 11580
rect 5997 11571 6055 11577
rect 6086 11568 6092 11580
rect 6144 11568 6150 11620
rect 6362 11568 6368 11620
rect 6420 11608 6426 11620
rect 7006 11608 7012 11620
rect 6420 11580 7012 11608
rect 6420 11568 6426 11580
rect 7006 11568 7012 11580
rect 7064 11568 7070 11620
rect 7285 11611 7343 11617
rect 7285 11577 7297 11611
rect 7331 11608 7343 11611
rect 8662 11608 8668 11620
rect 7331 11580 8668 11608
rect 7331 11577 7343 11580
rect 7285 11571 7343 11577
rect 8662 11568 8668 11580
rect 8720 11568 8726 11620
rect 10686 11608 10692 11620
rect 9232 11580 10692 11608
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 4816 11512 7205 11540
rect 7193 11509 7205 11512
rect 7239 11540 7251 11543
rect 9232 11540 9260 11580
rect 10686 11568 10692 11580
rect 10744 11568 10750 11620
rect 10870 11617 10876 11620
rect 10864 11608 10876 11617
rect 10831 11580 10876 11608
rect 10864 11571 10876 11580
rect 10870 11568 10876 11571
rect 10928 11568 10934 11620
rect 11882 11568 11888 11620
rect 11940 11608 11946 11620
rect 12682 11611 12740 11617
rect 12682 11608 12694 11611
rect 11940 11580 12694 11608
rect 11940 11568 11946 11580
rect 12682 11577 12694 11580
rect 12728 11577 12740 11611
rect 12682 11571 12740 11577
rect 7239 11512 9260 11540
rect 9309 11543 9367 11549
rect 7239 11509 7251 11512
rect 7193 11503 7251 11509
rect 9309 11509 9321 11543
rect 9355 11540 9367 11543
rect 9398 11540 9404 11552
rect 9355 11512 9404 11540
rect 9355 11509 9367 11512
rect 9309 11503 9367 11509
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 9677 11543 9735 11549
rect 9677 11540 9689 11543
rect 9640 11512 9689 11540
rect 9640 11500 9646 11512
rect 9677 11509 9689 11512
rect 9723 11509 9735 11543
rect 9677 11503 9735 11509
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 10137 11543 10195 11549
rect 10137 11540 10149 11543
rect 10008 11512 10149 11540
rect 10008 11500 10014 11512
rect 10137 11509 10149 11512
rect 10183 11540 10195 11543
rect 11974 11540 11980 11552
rect 10183 11512 11980 11540
rect 10183 11509 10195 11512
rect 10137 11503 10195 11509
rect 11974 11500 11980 11512
rect 12032 11500 12038 11552
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 14292 11540 14320 11639
rect 15194 11636 15200 11648
rect 15252 11636 15258 11688
rect 16301 11679 16359 11685
rect 16301 11645 16313 11679
rect 16347 11676 16359 11679
rect 16390 11676 16396 11688
rect 16347 11648 16396 11676
rect 16347 11645 16359 11648
rect 16301 11639 16359 11645
rect 16390 11636 16396 11648
rect 16448 11636 16454 11688
rect 16574 11685 16580 11688
rect 16568 11639 16580 11685
rect 16632 11676 16638 11688
rect 16632 11648 16668 11676
rect 16574 11636 16580 11639
rect 16632 11636 16638 11648
rect 16942 11636 16948 11688
rect 17000 11676 17006 11688
rect 17770 11676 17776 11688
rect 17000 11648 17776 11676
rect 17000 11636 17006 11648
rect 17770 11636 17776 11648
rect 17828 11636 17834 11688
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 18012 11648 18061 11676
rect 18012 11636 18018 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18156 11676 18184 11716
rect 18325 11713 18337 11747
rect 18371 11713 18383 11747
rect 18325 11707 18383 11713
rect 18966 11704 18972 11756
rect 19024 11744 19030 11756
rect 19337 11747 19395 11753
rect 19337 11744 19349 11747
rect 19024 11716 19349 11744
rect 19024 11704 19030 11716
rect 19337 11713 19349 11716
rect 19383 11713 19395 11747
rect 19337 11707 19395 11713
rect 19426 11704 19432 11756
rect 19484 11744 19490 11756
rect 20349 11747 20407 11753
rect 20349 11744 20361 11747
rect 19484 11716 20361 11744
rect 19484 11704 19490 11716
rect 20349 11713 20361 11716
rect 20395 11713 20407 11747
rect 20349 11707 20407 11713
rect 19245 11679 19303 11685
rect 19245 11676 19257 11679
rect 18156 11648 19257 11676
rect 18049 11639 18107 11645
rect 19245 11645 19257 11648
rect 19291 11645 19303 11679
rect 20162 11676 20168 11688
rect 20123 11648 20168 11676
rect 19245 11639 19303 11645
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 20809 11679 20867 11685
rect 20809 11645 20821 11679
rect 20855 11676 20867 11679
rect 20990 11676 20996 11688
rect 20855 11648 20996 11676
rect 20855 11645 20867 11648
rect 20809 11639 20867 11645
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 14636 11611 14694 11617
rect 14636 11577 14648 11611
rect 14682 11608 14694 11611
rect 15562 11608 15568 11620
rect 14682 11580 15568 11608
rect 14682 11577 14694 11580
rect 14636 11571 14694 11577
rect 15562 11568 15568 11580
rect 15620 11568 15626 11620
rect 19610 11608 19616 11620
rect 15678 11580 19616 11608
rect 12124 11512 14320 11540
rect 12124 11500 12130 11512
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15678 11540 15706 11580
rect 19610 11568 19616 11580
rect 19668 11568 19674 11620
rect 15436 11512 15706 11540
rect 15436 11500 15442 11512
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 17681 11543 17739 11549
rect 17681 11540 17693 11543
rect 17184 11512 17693 11540
rect 17184 11500 17190 11512
rect 17681 11509 17693 11512
rect 17727 11540 17739 11543
rect 18966 11540 18972 11552
rect 17727 11512 18972 11540
rect 17727 11509 17739 11512
rect 17681 11503 17739 11509
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 19150 11540 19156 11552
rect 19111 11512 19156 11540
rect 19150 11500 19156 11512
rect 19208 11500 19214 11552
rect 19426 11500 19432 11552
rect 19484 11540 19490 11552
rect 19797 11543 19855 11549
rect 19797 11540 19809 11543
rect 19484 11512 19809 11540
rect 19484 11500 19490 11512
rect 19797 11509 19809 11512
rect 19843 11509 19855 11543
rect 19797 11503 19855 11509
rect 20257 11543 20315 11549
rect 20257 11509 20269 11543
rect 20303 11540 20315 11543
rect 20714 11540 20720 11552
rect 20303 11512 20720 11540
rect 20303 11509 20315 11512
rect 20257 11503 20315 11509
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 1397 11339 1455 11345
rect 1397 11305 1409 11339
rect 1443 11336 1455 11339
rect 1486 11336 1492 11348
rect 1443 11308 1492 11336
rect 1443 11305 1455 11308
rect 1397 11299 1455 11305
rect 1486 11296 1492 11308
rect 1544 11296 1550 11348
rect 3234 11336 3240 11348
rect 3195 11308 3240 11336
rect 3234 11296 3240 11308
rect 3292 11296 3298 11348
rect 3326 11296 3332 11348
rect 3384 11336 3390 11348
rect 3513 11339 3571 11345
rect 3513 11336 3525 11339
rect 3384 11308 3525 11336
rect 3384 11296 3390 11308
rect 3513 11305 3525 11308
rect 3559 11305 3571 11339
rect 4062 11336 4068 11348
rect 4023 11308 4068 11336
rect 3513 11299 3571 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11305 5319 11339
rect 5261 11299 5319 11305
rect 2590 11268 2596 11280
rect 1872 11240 2596 11268
rect 1872 11209 1900 11240
rect 2590 11228 2596 11240
rect 2648 11228 2654 11280
rect 3878 11228 3884 11280
rect 3936 11268 3942 11280
rect 5276 11268 5304 11299
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6270 11336 6276 11348
rect 5868 11308 6276 11336
rect 5868 11296 5874 11308
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 7193 11339 7251 11345
rect 7193 11336 7205 11339
rect 7156 11308 7205 11336
rect 7156 11296 7162 11308
rect 7193 11305 7205 11308
rect 7239 11305 7251 11339
rect 7193 11299 7251 11305
rect 7377 11339 7435 11345
rect 7377 11305 7389 11339
rect 7423 11336 7435 11339
rect 7423 11308 8708 11336
rect 7423 11305 7435 11308
rect 7377 11299 7435 11305
rect 3936 11240 5304 11268
rect 6080 11271 6138 11277
rect 3936 11228 3942 11240
rect 6080 11237 6092 11271
rect 6126 11268 6138 11271
rect 6730 11268 6736 11280
rect 6126 11240 6736 11268
rect 6126 11237 6138 11240
rect 6080 11231 6138 11237
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 6822 11228 6828 11280
rect 6880 11268 6886 11280
rect 6880 11240 7972 11268
rect 6880 11228 6886 11240
rect 1857 11203 1915 11209
rect 1857 11169 1869 11203
rect 1903 11169 1915 11203
rect 1857 11163 1915 11169
rect 2124 11203 2182 11209
rect 2124 11169 2136 11203
rect 2170 11200 2182 11203
rect 2682 11200 2688 11212
rect 2170 11172 2688 11200
rect 2170 11169 2182 11172
rect 2124 11163 2182 11169
rect 2682 11160 2688 11172
rect 2740 11200 2746 11212
rect 2740 11172 3280 11200
rect 2740 11160 2746 11172
rect 3252 11076 3280 11172
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4212 11172 4445 11200
rect 4212 11160 4218 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 5074 11200 5080 11212
rect 5035 11172 5080 11200
rect 4433 11163 4491 11169
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 7742 11209 7748 11212
rect 7469 11203 7527 11209
rect 7469 11200 7481 11203
rect 6972 11172 7481 11200
rect 6972 11160 6978 11172
rect 7469 11169 7481 11172
rect 7515 11169 7527 11203
rect 7469 11163 7527 11169
rect 7736 11163 7748 11209
rect 7800 11200 7806 11212
rect 7944 11200 7972 11240
rect 8110 11228 8116 11280
rect 8168 11268 8174 11280
rect 8386 11268 8392 11280
rect 8168 11240 8392 11268
rect 8168 11228 8174 11240
rect 8386 11228 8392 11240
rect 8444 11228 8450 11280
rect 8680 11268 8708 11308
rect 8754 11296 8760 11348
rect 8812 11336 8818 11348
rect 8849 11339 8907 11345
rect 8849 11336 8861 11339
rect 8812 11308 8861 11336
rect 8812 11296 8818 11308
rect 8849 11305 8861 11308
rect 8895 11305 8907 11339
rect 8849 11299 8907 11305
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 9674 11336 9680 11348
rect 9088 11308 9680 11336
rect 9088 11296 9094 11308
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10226 11336 10232 11348
rect 9784 11308 10232 11336
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 8680 11240 8953 11268
rect 8941 11237 8953 11240
rect 8987 11237 8999 11271
rect 8941 11231 8999 11237
rect 9125 11271 9183 11277
rect 9125 11237 9137 11271
rect 9171 11268 9183 11271
rect 9784 11268 9812 11308
rect 10226 11296 10232 11308
rect 10284 11296 10290 11348
rect 10686 11296 10692 11348
rect 10744 11336 10750 11348
rect 11698 11336 11704 11348
rect 10744 11308 11704 11336
rect 10744 11296 10750 11308
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 11977 11339 12035 11345
rect 11977 11305 11989 11339
rect 12023 11336 12035 11339
rect 12066 11336 12072 11348
rect 12023 11308 12072 11336
rect 12023 11305 12035 11308
rect 11977 11299 12035 11305
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 15657 11339 15715 11345
rect 15657 11336 15669 11339
rect 12544 11308 15669 11336
rect 9171 11240 9812 11268
rect 9876 11240 10171 11268
rect 9171 11237 9183 11240
rect 9125 11231 9183 11237
rect 9876 11200 9904 11240
rect 7800 11172 7836 11200
rect 7944 11172 9904 11200
rect 7742 11160 7748 11163
rect 7800 11160 7806 11172
rect 9950 11160 9956 11212
rect 10008 11200 10014 11212
rect 10143 11200 10171 11240
rect 10410 11228 10416 11280
rect 10468 11268 10474 11280
rect 10505 11271 10563 11277
rect 10505 11268 10517 11271
rect 10468 11240 10517 11268
rect 10468 11228 10474 11240
rect 10505 11237 10517 11240
rect 10551 11237 10563 11271
rect 10505 11231 10563 11237
rect 11514 11228 11520 11280
rect 11572 11268 11578 11280
rect 12544 11268 12572 11308
rect 15657 11305 15669 11308
rect 15703 11305 15715 11339
rect 15657 11299 15715 11305
rect 15749 11339 15807 11345
rect 15749 11305 15761 11339
rect 15795 11336 15807 11339
rect 15838 11336 15844 11348
rect 15795 11308 15844 11336
rect 15795 11305 15807 11308
rect 15749 11299 15807 11305
rect 15378 11268 15384 11280
rect 11572 11240 12572 11268
rect 12636 11240 15384 11268
rect 11572 11228 11578 11240
rect 12158 11200 12164 11212
rect 10008 11172 10101 11200
rect 10143 11172 12164 11200
rect 10008 11160 10014 11172
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 12636 11200 12664 11240
rect 15378 11228 15384 11240
rect 15436 11228 15442 11280
rect 12268 11172 12664 11200
rect 12704 11203 12762 11209
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 4304 11104 4537 11132
rect 4304 11092 4310 11104
rect 4525 11101 4537 11104
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 3234 11024 3240 11076
rect 3292 11064 3298 11076
rect 4632 11064 4660 11095
rect 5626 11092 5632 11144
rect 5684 11132 5690 11144
rect 5813 11135 5871 11141
rect 5813 11132 5825 11135
rect 5684 11104 5825 11132
rect 5684 11092 5690 11104
rect 5813 11101 5825 11104
rect 5859 11101 5871 11135
rect 5813 11095 5871 11101
rect 7006 11092 7012 11144
rect 7064 11132 7070 11144
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 7064 11104 7389 11132
rect 7064 11092 7070 11104
rect 7377 11101 7389 11104
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 3292 11036 4660 11064
rect 3292 11024 3298 11036
rect 4706 11024 4712 11076
rect 4764 11064 4770 11076
rect 5718 11064 5724 11076
rect 4764 11036 5724 11064
rect 4764 11024 4770 11036
rect 5718 11024 5724 11036
rect 5776 11024 5782 11076
rect 8941 11067 8999 11073
rect 8941 11033 8953 11067
rect 8987 11064 8999 11067
rect 9968 11064 9996 11160
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 12268 11132 12296 11172
rect 12704 11169 12716 11203
rect 12750 11200 12762 11203
rect 13722 11200 13728 11212
rect 12750 11172 13728 11200
rect 12750 11169 12762 11172
rect 12704 11163 12762 11169
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 13998 11160 14004 11212
rect 14056 11200 14062 11212
rect 14461 11203 14519 11209
rect 14461 11200 14473 11203
rect 14056 11172 14473 11200
rect 14056 11160 14062 11172
rect 14461 11169 14473 11172
rect 14507 11169 14519 11203
rect 14461 11163 14519 11169
rect 14550 11160 14556 11212
rect 14608 11200 14614 11212
rect 15672 11200 15700 11299
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 16577 11339 16635 11345
rect 16577 11305 16589 11339
rect 16623 11336 16635 11339
rect 18049 11339 18107 11345
rect 18049 11336 18061 11339
rect 16623 11308 18061 11336
rect 16623 11305 16635 11308
rect 16577 11299 16635 11305
rect 18049 11305 18061 11308
rect 18095 11305 18107 11339
rect 18049 11299 18107 11305
rect 18414 11296 18420 11348
rect 18472 11336 18478 11348
rect 18785 11339 18843 11345
rect 18472 11308 18736 11336
rect 18472 11296 18478 11308
rect 16850 11228 16856 11280
rect 16908 11268 16914 11280
rect 17037 11271 17095 11277
rect 17037 11268 17049 11271
rect 16908 11240 17049 11268
rect 16908 11228 16914 11240
rect 17037 11237 17049 11240
rect 17083 11237 17095 11271
rect 17497 11271 17555 11277
rect 17497 11268 17509 11271
rect 17037 11231 17095 11237
rect 17144 11240 17509 11268
rect 16945 11203 17003 11209
rect 14608 11172 14653 11200
rect 14752 11172 15516 11200
rect 15672 11172 16896 11200
rect 14608 11160 14614 11172
rect 12434 11132 12440 11144
rect 12032 11104 12296 11132
rect 12395 11104 12440 11132
rect 12032 11092 12038 11104
rect 12434 11092 12440 11104
rect 12492 11092 12498 11144
rect 14752 11141 14780 11172
rect 14737 11135 14795 11141
rect 14737 11132 14749 11135
rect 13832 11104 14749 11132
rect 11514 11064 11520 11076
rect 8987 11036 9996 11064
rect 10060 11036 11520 11064
rect 8987 11033 8999 11036
rect 8941 11027 8999 11033
rect 4062 10956 4068 11008
rect 4120 10996 4126 11008
rect 10060 10996 10088 11036
rect 11514 11024 11520 11036
rect 11572 11024 11578 11076
rect 11790 11024 11796 11076
rect 11848 11064 11854 11076
rect 12066 11064 12072 11076
rect 11848 11036 12072 11064
rect 11848 11024 11854 11036
rect 12066 11024 12072 11036
rect 12124 11024 12130 11076
rect 13832 11073 13860 11104
rect 14737 11101 14749 11104
rect 14783 11101 14795 11135
rect 15488 11132 15516 11172
rect 15933 11135 15991 11141
rect 15933 11132 15945 11135
rect 15488 11104 15945 11132
rect 14737 11095 14795 11101
rect 15933 11101 15945 11104
rect 15979 11132 15991 11135
rect 16390 11132 16396 11144
rect 15979 11104 16396 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 13817 11067 13875 11073
rect 13817 11064 13829 11067
rect 13372 11036 13829 11064
rect 4120 10968 10088 10996
rect 10137 10999 10195 11005
rect 4120 10956 4126 10968
rect 10137 10965 10149 10999
rect 10183 10996 10195 10999
rect 12618 10996 12624 11008
rect 10183 10968 12624 10996
rect 10183 10965 10195 10968
rect 10137 10959 10195 10965
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 12802 10956 12808 11008
rect 12860 10996 12866 11008
rect 13372 10996 13400 11036
rect 13817 11033 13829 11036
rect 13863 11033 13875 11067
rect 13817 11027 13875 11033
rect 13906 11024 13912 11076
rect 13964 11064 13970 11076
rect 15289 11067 15347 11073
rect 15289 11064 15301 11067
rect 13964 11036 15301 11064
rect 13964 11024 13970 11036
rect 15289 11033 15301 11036
rect 15335 11033 15347 11067
rect 16868 11064 16896 11172
rect 16945 11169 16957 11203
rect 16991 11200 17003 11203
rect 17144 11200 17172 11240
rect 17497 11237 17509 11240
rect 17543 11237 17555 11271
rect 17497 11231 17555 11237
rect 17770 11228 17776 11280
rect 17828 11268 17834 11280
rect 17828 11240 18644 11268
rect 17828 11228 17834 11240
rect 16991 11172 17172 11200
rect 16991 11169 17003 11172
rect 16945 11163 17003 11169
rect 17218 11160 17224 11212
rect 17276 11200 17282 11212
rect 18616 11209 18644 11240
rect 17957 11203 18015 11209
rect 17957 11200 17969 11203
rect 17276 11172 17969 11200
rect 17276 11160 17282 11172
rect 17957 11169 17969 11172
rect 18003 11169 18015 11203
rect 17957 11163 18015 11169
rect 18601 11203 18659 11209
rect 18601 11169 18613 11203
rect 18647 11169 18659 11203
rect 18708 11200 18736 11308
rect 18785 11305 18797 11339
rect 18831 11305 18843 11339
rect 18785 11299 18843 11305
rect 18800 11268 18828 11299
rect 19150 11296 19156 11348
rect 19208 11336 19214 11348
rect 20901 11339 20959 11345
rect 20901 11336 20913 11339
rect 19208 11308 20913 11336
rect 19208 11296 19214 11308
rect 20901 11305 20913 11308
rect 20947 11305 20959 11339
rect 20901 11299 20959 11305
rect 19242 11268 19248 11280
rect 18800 11240 19248 11268
rect 19242 11228 19248 11240
rect 19300 11228 19306 11280
rect 19420 11271 19478 11277
rect 19420 11237 19432 11271
rect 19466 11268 19478 11271
rect 20346 11268 20352 11280
rect 19466 11240 20352 11268
rect 19466 11237 19478 11240
rect 19420 11231 19478 11237
rect 20346 11228 20352 11240
rect 20404 11228 20410 11280
rect 20622 11200 20628 11212
rect 18708 11172 20628 11200
rect 18601 11163 18659 11169
rect 17126 11132 17132 11144
rect 17087 11104 17132 11132
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11132 18291 11135
rect 18782 11132 18788 11144
rect 18279 11104 18788 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 19153 11135 19211 11141
rect 19153 11101 19165 11135
rect 19199 11101 19211 11135
rect 19153 11095 19211 11101
rect 17310 11064 17316 11076
rect 16868 11036 17316 11064
rect 15289 11027 15347 11033
rect 17310 11024 17316 11036
rect 17368 11024 17374 11076
rect 17497 11067 17555 11073
rect 17497 11033 17509 11067
rect 17543 11064 17555 11067
rect 17954 11064 17960 11076
rect 17543 11036 17960 11064
rect 17543 11033 17555 11036
rect 17497 11027 17555 11033
rect 17954 11024 17960 11036
rect 18012 11024 18018 11076
rect 18064 11036 18644 11064
rect 14090 10996 14096 11008
rect 12860 10968 13400 10996
rect 14051 10968 14096 10996
rect 12860 10956 12866 10968
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 14182 10956 14188 11008
rect 14240 10996 14246 11008
rect 16666 10996 16672 11008
rect 14240 10968 16672 10996
rect 14240 10956 14246 10968
rect 16666 10956 16672 10968
rect 16724 10956 16730 11008
rect 17589 10999 17647 11005
rect 17589 10965 17601 10999
rect 17635 10996 17647 10999
rect 18064 10996 18092 11036
rect 17635 10968 18092 10996
rect 18616 10996 18644 11036
rect 18690 11024 18696 11076
rect 18748 11064 18754 11076
rect 19168 11064 19196 11095
rect 20548 11073 20576 11172
rect 20622 11160 20628 11172
rect 20680 11160 20686 11212
rect 18748 11036 19196 11064
rect 20533 11067 20591 11073
rect 18748 11024 18754 11036
rect 20533 11033 20545 11067
rect 20579 11033 20591 11067
rect 20533 11027 20591 11033
rect 19794 10996 19800 11008
rect 18616 10968 19800 10996
rect 17635 10965 17647 10968
rect 17589 10959 17647 10965
rect 19794 10956 19800 10968
rect 19852 10956 19858 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 3234 10792 3240 10804
rect 1820 10764 2820 10792
rect 3195 10764 3240 10792
rect 1820 10752 1826 10764
rect 2792 10724 2820 10764
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 3697 10795 3755 10801
rect 3697 10761 3709 10795
rect 3743 10792 3755 10795
rect 3786 10792 3792 10804
rect 3743 10764 3792 10792
rect 3743 10761 3755 10764
rect 3697 10755 3755 10761
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 4246 10752 4252 10804
rect 4304 10792 4310 10804
rect 4433 10795 4491 10801
rect 4433 10792 4445 10795
rect 4304 10764 4445 10792
rect 4304 10752 4310 10764
rect 4433 10761 4445 10764
rect 4479 10761 4491 10795
rect 6730 10792 6736 10804
rect 4433 10755 4491 10761
rect 5000 10764 6736 10792
rect 4338 10724 4344 10736
rect 2792 10696 4344 10724
rect 4338 10684 4344 10696
rect 4396 10684 4402 10736
rect 5000 10656 5028 10764
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 7374 10752 7380 10804
rect 7432 10792 7438 10804
rect 8570 10792 8576 10804
rect 7432 10764 8576 10792
rect 7432 10752 7438 10764
rect 8570 10752 8576 10764
rect 8628 10792 8634 10804
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 8628 10764 8861 10792
rect 8628 10752 8634 10764
rect 8849 10761 8861 10764
rect 8895 10761 8907 10795
rect 8849 10755 8907 10761
rect 8938 10752 8944 10804
rect 8996 10792 9002 10804
rect 11790 10792 11796 10804
rect 8996 10764 11796 10792
rect 8996 10752 9002 10764
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 12032 10764 12173 10792
rect 12032 10752 12038 10764
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 12161 10755 12219 10761
rect 12986 10752 12992 10804
rect 13044 10792 13050 10804
rect 13044 10764 13952 10792
rect 13044 10752 13050 10764
rect 5258 10684 5264 10736
rect 5316 10724 5322 10736
rect 7653 10727 7711 10733
rect 5316 10696 6040 10724
rect 5316 10684 5322 10696
rect 3528 10628 5028 10656
rect 5077 10659 5135 10665
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 3234 10588 3240 10600
rect 1903 10560 3240 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 3528 10597 3556 10628
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5442 10656 5448 10668
rect 5123 10628 5448 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 5902 10656 5908 10668
rect 5863 10628 5908 10656
rect 5902 10616 5908 10628
rect 5960 10616 5966 10668
rect 6012 10665 6040 10696
rect 7653 10693 7665 10727
rect 7699 10724 7711 10727
rect 8110 10724 8116 10736
rect 7699 10696 8116 10724
rect 7699 10693 7711 10696
rect 7653 10687 7711 10693
rect 8110 10684 8116 10696
rect 8168 10684 8174 10736
rect 9306 10724 9312 10736
rect 9267 10696 9312 10724
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 10778 10684 10784 10736
rect 10836 10724 10842 10736
rect 11057 10727 11115 10733
rect 11057 10724 11069 10727
rect 10836 10696 11069 10724
rect 10836 10684 10842 10696
rect 11057 10693 11069 10696
rect 11103 10693 11115 10727
rect 11057 10687 11115 10693
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 12526 10724 12532 10736
rect 11388 10696 12532 10724
rect 11388 10684 11394 10696
rect 12526 10684 12532 10696
rect 12584 10724 12590 10736
rect 13170 10724 13176 10736
rect 12584 10696 13176 10724
rect 12584 10684 12590 10696
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 13446 10724 13452 10736
rect 13407 10696 13452 10724
rect 13446 10684 13452 10696
rect 13504 10684 13510 10736
rect 13924 10724 13952 10764
rect 14366 10752 14372 10804
rect 14424 10792 14430 10804
rect 16022 10792 16028 10804
rect 14424 10764 16028 10792
rect 14424 10752 14430 10764
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 16945 10795 17003 10801
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 17218 10792 17224 10804
rect 16991 10764 17224 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 19150 10792 19156 10804
rect 17512 10764 19156 10792
rect 14737 10727 14795 10733
rect 13924 10696 14044 10724
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6362 10616 6368 10668
rect 6420 10656 6426 10668
rect 7469 10659 7527 10665
rect 6420 10628 7420 10656
rect 6420 10616 6426 10628
rect 3513 10591 3571 10597
rect 3513 10557 3525 10591
rect 3559 10557 3571 10591
rect 3513 10551 3571 10557
rect 4893 10591 4951 10597
rect 4893 10557 4905 10591
rect 4939 10588 4951 10591
rect 6822 10588 6828 10600
rect 4939 10560 6828 10588
rect 4939 10557 4951 10560
rect 4893 10551 4951 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 7392 10588 7420 10628
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 7558 10656 7564 10668
rect 7515 10628 7564 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 8202 10588 8208 10600
rect 7392 10560 8208 10588
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 8404 10532 8432 10619
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11296 10628 11713 10656
rect 11296 10616 11302 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13722 10656 13728 10668
rect 13127 10628 13728 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 13906 10656 13912 10668
rect 13867 10628 13912 10656
rect 13906 10616 13912 10628
rect 13964 10616 13970 10668
rect 14016 10665 14044 10696
rect 14737 10693 14749 10727
rect 14783 10693 14795 10727
rect 14737 10687 14795 10693
rect 15933 10727 15991 10733
rect 15933 10693 15945 10727
rect 15979 10724 15991 10727
rect 17512 10724 17540 10764
rect 19150 10752 19156 10764
rect 19208 10752 19214 10804
rect 20993 10795 21051 10801
rect 20993 10761 21005 10795
rect 21039 10792 21051 10795
rect 21174 10792 21180 10804
rect 21039 10764 21180 10792
rect 21039 10761 21051 10764
rect 20993 10755 21051 10761
rect 21174 10752 21180 10764
rect 21232 10752 21238 10804
rect 15979 10696 17540 10724
rect 15979 10693 15991 10696
rect 15933 10687 15991 10693
rect 14001 10659 14059 10665
rect 14001 10625 14013 10659
rect 14047 10625 14059 10659
rect 14752 10656 14780 10687
rect 15378 10656 15384 10668
rect 14752 10628 15240 10656
rect 15339 10628 15384 10656
rect 14001 10619 14059 10625
rect 8938 10548 8944 10600
rect 8996 10588 9002 10600
rect 9033 10591 9091 10597
rect 9033 10588 9045 10591
rect 8996 10560 9045 10588
rect 8996 10548 9002 10560
rect 9033 10557 9045 10560
rect 9079 10557 9091 10591
rect 9033 10551 9091 10557
rect 9125 10591 9183 10597
rect 9125 10557 9137 10591
rect 9171 10588 9183 10591
rect 9490 10588 9496 10600
rect 9171 10560 9496 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 9490 10548 9496 10560
rect 9548 10548 9554 10600
rect 9582 10548 9588 10600
rect 9640 10588 9646 10600
rect 9677 10591 9735 10597
rect 9677 10588 9689 10591
rect 9640 10560 9689 10588
rect 9640 10548 9646 10560
rect 9677 10557 9689 10560
rect 9723 10557 9735 10591
rect 10870 10588 10876 10600
rect 9677 10551 9735 10557
rect 9876 10560 10876 10588
rect 2124 10523 2182 10529
rect 2124 10489 2136 10523
rect 2170 10520 2182 10523
rect 2590 10520 2596 10532
rect 2170 10492 2596 10520
rect 2170 10489 2182 10492
rect 2124 10483 2182 10489
rect 2590 10480 2596 10492
rect 2648 10480 2654 10532
rect 2774 10480 2780 10532
rect 2832 10520 2838 10532
rect 3970 10520 3976 10532
rect 2832 10492 3976 10520
rect 2832 10480 2838 10492
rect 3970 10480 3976 10492
rect 4028 10480 4034 10532
rect 4801 10523 4859 10529
rect 4801 10489 4813 10523
rect 4847 10520 4859 10523
rect 4847 10492 5488 10520
rect 4847 10489 4859 10492
rect 4801 10483 4859 10489
rect 1397 10455 1455 10461
rect 1397 10421 1409 10455
rect 1443 10452 1455 10455
rect 3326 10452 3332 10464
rect 1443 10424 3332 10452
rect 1443 10421 1455 10424
rect 1397 10415 1455 10421
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 5460 10461 5488 10492
rect 5718 10480 5724 10532
rect 5776 10520 5782 10532
rect 5813 10523 5871 10529
rect 5813 10520 5825 10523
rect 5776 10492 5825 10520
rect 5776 10480 5782 10492
rect 5813 10489 5825 10492
rect 5859 10520 5871 10523
rect 6730 10520 6736 10532
rect 5859 10492 6736 10520
rect 5859 10489 5871 10492
rect 5813 10483 5871 10489
rect 6730 10480 6736 10492
rect 6788 10480 6794 10532
rect 7282 10520 7288 10532
rect 7243 10492 7288 10520
rect 7282 10480 7288 10492
rect 7340 10480 7346 10532
rect 7558 10480 7564 10532
rect 7616 10520 7622 10532
rect 8386 10520 8392 10532
rect 7616 10492 8392 10520
rect 7616 10480 7622 10492
rect 8386 10480 8392 10492
rect 8444 10480 8450 10532
rect 8754 10480 8760 10532
rect 8812 10520 8818 10532
rect 9876 10520 9904 10560
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 11112 10560 11529 10588
rect 11112 10548 11118 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 11606 10548 11612 10600
rect 11664 10588 11670 10600
rect 11974 10588 11980 10600
rect 11664 10560 11709 10588
rect 11935 10560 11980 10588
rect 11664 10548 11670 10560
rect 11974 10548 11980 10560
rect 12032 10548 12038 10600
rect 12342 10548 12348 10600
rect 12400 10588 12406 10600
rect 13817 10591 13875 10597
rect 12400 10560 13768 10588
rect 12400 10548 12406 10560
rect 8812 10492 9904 10520
rect 9944 10523 10002 10529
rect 8812 10480 8818 10492
rect 9944 10489 9956 10523
rect 9990 10520 10002 10523
rect 11238 10520 11244 10532
rect 9990 10492 11244 10520
rect 9990 10489 10002 10492
rect 9944 10483 10002 10489
rect 11238 10480 11244 10492
rect 11296 10480 11302 10532
rect 11698 10480 11704 10532
rect 11756 10520 11762 10532
rect 12897 10523 12955 10529
rect 12897 10520 12909 10523
rect 11756 10492 12909 10520
rect 11756 10480 11762 10492
rect 12897 10489 12909 10492
rect 12943 10489 12955 10523
rect 12897 10483 12955 10489
rect 5445 10455 5503 10461
rect 5445 10421 5457 10455
rect 5491 10421 5503 10455
rect 5445 10415 5503 10421
rect 6086 10412 6092 10464
rect 6144 10452 6150 10464
rect 6825 10455 6883 10461
rect 6825 10452 6837 10455
rect 6144 10424 6837 10452
rect 6144 10412 6150 10424
rect 6825 10421 6837 10424
rect 6871 10421 6883 10455
rect 6825 10415 6883 10421
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7193 10455 7251 10461
rect 7193 10452 7205 10455
rect 6972 10424 7205 10452
rect 6972 10412 6978 10424
rect 7193 10421 7205 10424
rect 7239 10452 7251 10455
rect 7653 10455 7711 10461
rect 7653 10452 7665 10455
rect 7239 10424 7665 10452
rect 7239 10421 7251 10424
rect 7193 10415 7251 10421
rect 7653 10421 7665 10424
rect 7699 10421 7711 10455
rect 7653 10415 7711 10421
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7800 10424 7849 10452
rect 7800 10412 7806 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 8202 10452 8208 10464
rect 8163 10424 8208 10452
rect 7837 10415 7895 10421
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8297 10455 8355 10461
rect 8297 10421 8309 10455
rect 8343 10452 8355 10455
rect 10318 10452 10324 10464
rect 8343 10424 10324 10452
rect 8343 10421 8355 10424
rect 8297 10415 8355 10421
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11149 10455 11207 10461
rect 11149 10452 11161 10455
rect 11112 10424 11161 10452
rect 11112 10412 11118 10424
rect 11149 10421 11161 10424
rect 11195 10421 11207 10455
rect 11149 10415 11207 10421
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12710 10452 12716 10464
rect 12483 10424 12716 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 12805 10455 12863 10461
rect 12805 10421 12817 10455
rect 12851 10452 12863 10455
rect 13170 10452 13176 10464
rect 12851 10424 13176 10452
rect 12851 10421 12863 10424
rect 12805 10415 12863 10421
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 13740 10452 13768 10560
rect 13817 10557 13829 10591
rect 13863 10588 13875 10591
rect 14090 10588 14096 10600
rect 13863 10560 14096 10588
rect 13863 10557 13875 10560
rect 13817 10551 13875 10557
rect 14090 10548 14096 10560
rect 14148 10548 14154 10600
rect 14182 10548 14188 10600
rect 14240 10588 14246 10600
rect 15105 10591 15163 10597
rect 15105 10588 15117 10591
rect 14240 10560 15117 10588
rect 14240 10548 14246 10560
rect 15105 10557 15117 10560
rect 15151 10557 15163 10591
rect 15212 10588 15240 10628
rect 15378 10616 15384 10628
rect 15436 10616 15442 10668
rect 15562 10616 15568 10668
rect 15620 10656 15626 10668
rect 16482 10656 16488 10668
rect 15620 10628 16488 10656
rect 15620 10616 15626 10628
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 16577 10659 16635 10665
rect 16577 10625 16589 10659
rect 16623 10656 16635 10659
rect 16850 10656 16856 10668
rect 16623 10628 16856 10656
rect 16623 10625 16635 10628
rect 16577 10619 16635 10625
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 17126 10616 17132 10668
rect 17184 10656 17190 10668
rect 17497 10659 17555 10665
rect 17497 10656 17509 10659
rect 17184 10628 17509 10656
rect 17184 10616 17190 10628
rect 17497 10625 17509 10628
rect 17543 10625 17555 10659
rect 17497 10619 17555 10625
rect 20162 10616 20168 10668
rect 20220 10656 20226 10668
rect 20349 10659 20407 10665
rect 20349 10656 20361 10659
rect 20220 10628 20361 10656
rect 20220 10616 20226 10628
rect 20349 10625 20361 10628
rect 20395 10656 20407 10659
rect 20622 10656 20628 10668
rect 20395 10628 20628 10656
rect 20395 10625 20407 10628
rect 20349 10619 20407 10625
rect 20622 10616 20628 10628
rect 20680 10616 20686 10668
rect 16393 10591 16451 10597
rect 16393 10588 16405 10591
rect 15212 10560 16405 10588
rect 15105 10551 15163 10557
rect 16393 10557 16405 10560
rect 16439 10557 16451 10591
rect 16393 10551 16451 10557
rect 16942 10548 16948 10600
rect 17000 10588 17006 10600
rect 17313 10591 17371 10597
rect 17313 10588 17325 10591
rect 17000 10560 17325 10588
rect 17000 10548 17006 10560
rect 17313 10557 17325 10560
rect 17359 10557 17371 10591
rect 17313 10551 17371 10557
rect 18141 10591 18199 10597
rect 18141 10557 18153 10591
rect 18187 10557 18199 10591
rect 18141 10551 18199 10557
rect 18408 10591 18466 10597
rect 18408 10557 18420 10591
rect 18454 10588 18466 10591
rect 18874 10588 18880 10600
rect 18454 10560 18880 10588
rect 18454 10557 18466 10560
rect 18408 10551 18466 10557
rect 13906 10480 13912 10532
rect 13964 10520 13970 10532
rect 13964 10492 14679 10520
rect 13964 10480 13970 10492
rect 14550 10452 14556 10464
rect 13740 10424 14556 10452
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 14651 10452 14679 10492
rect 14918 10480 14924 10532
rect 14976 10520 14982 10532
rect 18046 10520 18052 10532
rect 14976 10492 18052 10520
rect 14976 10480 14982 10492
rect 18046 10480 18052 10492
rect 18104 10480 18110 10532
rect 18156 10520 18184 10551
rect 18874 10548 18880 10560
rect 18932 10548 18938 10600
rect 18966 10548 18972 10600
rect 19024 10588 19030 10600
rect 20530 10588 20536 10600
rect 19024 10560 20536 10588
rect 19024 10548 19030 10560
rect 20530 10548 20536 10560
rect 20588 10548 20594 10600
rect 20809 10591 20867 10597
rect 20809 10557 20821 10591
rect 20855 10588 20867 10591
rect 20898 10588 20904 10600
rect 20855 10560 20904 10588
rect 20855 10557 20867 10560
rect 20809 10551 20867 10557
rect 20898 10548 20904 10560
rect 20956 10548 20962 10600
rect 18230 10520 18236 10532
rect 18143 10492 18236 10520
rect 18230 10480 18236 10492
rect 18288 10520 18294 10532
rect 18690 10520 18696 10532
rect 18288 10492 18696 10520
rect 18288 10480 18294 10492
rect 18690 10480 18696 10492
rect 18748 10480 18754 10532
rect 18782 10480 18788 10532
rect 18840 10520 18846 10532
rect 18840 10492 20300 10520
rect 18840 10480 18846 10492
rect 15197 10455 15255 10461
rect 15197 10452 15209 10455
rect 14651 10424 15209 10452
rect 15197 10421 15209 10424
rect 15243 10421 15255 10455
rect 15197 10415 15255 10421
rect 16301 10455 16359 10461
rect 16301 10421 16313 10455
rect 16347 10452 16359 10455
rect 17218 10452 17224 10464
rect 16347 10424 17224 10452
rect 16347 10421 16359 10424
rect 16301 10415 16359 10421
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 17310 10412 17316 10464
rect 17368 10452 17374 10464
rect 17405 10455 17463 10461
rect 17405 10452 17417 10455
rect 17368 10424 17417 10452
rect 17368 10412 17374 10424
rect 17405 10421 17417 10424
rect 17451 10421 17463 10455
rect 17405 10415 17463 10421
rect 17586 10412 17592 10464
rect 17644 10452 17650 10464
rect 19521 10455 19579 10461
rect 19521 10452 19533 10455
rect 17644 10424 19533 10452
rect 17644 10412 17650 10424
rect 19521 10421 19533 10424
rect 19567 10421 19579 10455
rect 19794 10452 19800 10464
rect 19755 10424 19800 10452
rect 19521 10415 19579 10421
rect 19794 10412 19800 10424
rect 19852 10412 19858 10464
rect 20070 10412 20076 10464
rect 20128 10452 20134 10464
rect 20272 10461 20300 10492
rect 20165 10455 20223 10461
rect 20165 10452 20177 10455
rect 20128 10424 20177 10452
rect 20128 10412 20134 10424
rect 20165 10421 20177 10424
rect 20211 10421 20223 10455
rect 20165 10415 20223 10421
rect 20257 10455 20315 10461
rect 20257 10421 20269 10455
rect 20303 10452 20315 10455
rect 21910 10452 21916 10464
rect 20303 10424 21916 10452
rect 20303 10421 20315 10424
rect 20257 10415 20315 10421
rect 21910 10412 21916 10424
rect 21968 10412 21974 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 1670 10248 1676 10260
rect 1631 10220 1676 10248
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 3237 10251 3295 10257
rect 3237 10248 3249 10251
rect 2924 10220 3249 10248
rect 2924 10208 2930 10220
rect 3237 10217 3249 10220
rect 3283 10217 3295 10251
rect 6362 10248 6368 10260
rect 3237 10211 3295 10217
rect 4172 10220 6368 10248
rect 2409 10183 2467 10189
rect 2409 10149 2421 10183
rect 2455 10180 2467 10183
rect 2774 10180 2780 10192
rect 2455 10152 2780 10180
rect 2455 10149 2467 10152
rect 2409 10143 2467 10149
rect 2774 10140 2780 10152
rect 2832 10140 2838 10192
rect 4172 10180 4200 10220
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 6917 10251 6975 10257
rect 6917 10217 6929 10251
rect 6963 10248 6975 10251
rect 7742 10248 7748 10260
rect 6963 10220 7748 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 8205 10251 8263 10257
rect 8205 10217 8217 10251
rect 8251 10248 8263 10251
rect 8662 10248 8668 10260
rect 8251 10220 8668 10248
rect 8251 10217 8263 10220
rect 8205 10211 8263 10217
rect 8662 10208 8668 10220
rect 8720 10248 8726 10260
rect 8846 10248 8852 10260
rect 8720 10220 8852 10248
rect 8720 10208 8726 10220
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 9214 10248 9220 10260
rect 9175 10220 9220 10248
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 11330 10248 11336 10260
rect 9548 10220 11336 10248
rect 9548 10208 9554 10220
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 11425 10251 11483 10257
rect 11425 10217 11437 10251
rect 11471 10248 11483 10251
rect 11698 10248 11704 10260
rect 11471 10220 11704 10248
rect 11471 10217 11483 10220
rect 11425 10211 11483 10217
rect 11698 10208 11704 10220
rect 11756 10208 11762 10260
rect 11885 10251 11943 10257
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 12434 10248 12440 10260
rect 11931 10220 12440 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 13538 10248 13544 10260
rect 12719 10220 13544 10248
rect 3068 10152 4200 10180
rect 1489 10115 1547 10121
rect 1489 10081 1501 10115
rect 1535 10112 1547 10115
rect 1854 10112 1860 10124
rect 1535 10084 1860 10112
rect 1535 10081 1547 10084
rect 1489 10075 1547 10081
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 2498 10112 2504 10124
rect 2459 10084 2504 10112
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 3068 10121 3096 10152
rect 4246 10140 4252 10192
rect 4304 10189 4310 10192
rect 4304 10183 4368 10189
rect 4304 10149 4322 10183
rect 4356 10149 4368 10183
rect 4304 10143 4368 10149
rect 7009 10183 7067 10189
rect 7009 10149 7021 10183
rect 7055 10180 7067 10183
rect 12618 10180 12624 10192
rect 7055 10152 12624 10180
rect 7055 10149 7067 10152
rect 7009 10143 7067 10149
rect 4304 10140 4310 10143
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 3053 10115 3111 10121
rect 3053 10081 3065 10115
rect 3099 10081 3111 10115
rect 3053 10075 3111 10081
rect 3234 10072 3240 10124
rect 3292 10112 3298 10124
rect 4062 10112 4068 10124
rect 3292 10084 4068 10112
rect 3292 10072 3298 10084
rect 4062 10072 4068 10084
rect 4120 10112 4126 10124
rect 5626 10112 5632 10124
rect 4120 10084 5632 10112
rect 4120 10072 4126 10084
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 5902 10072 5908 10124
rect 5960 10112 5966 10124
rect 6089 10115 6147 10121
rect 6089 10112 6101 10115
rect 5960 10084 6101 10112
rect 5960 10072 5966 10084
rect 6089 10081 6101 10084
rect 6135 10081 6147 10115
rect 6089 10075 6147 10081
rect 7374 10072 7380 10124
rect 7432 10112 7438 10124
rect 8110 10112 8116 10124
rect 7432 10084 8116 10112
rect 7432 10072 7438 10084
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 8570 10072 8576 10124
rect 8628 10112 8634 10124
rect 8941 10115 8999 10121
rect 8941 10112 8953 10115
rect 8628 10084 8953 10112
rect 8628 10072 8634 10084
rect 8941 10081 8953 10084
rect 8987 10081 8999 10115
rect 8941 10075 8999 10081
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 9088 10084 9133 10112
rect 9088 10072 9094 10084
rect 9398 10072 9404 10124
rect 9456 10112 9462 10124
rect 9582 10112 9588 10124
rect 9456 10084 9588 10112
rect 9456 10072 9462 10084
rect 9582 10072 9588 10084
rect 9640 10112 9646 10124
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9640 10084 9689 10112
rect 9640 10072 9646 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 9933 10115 9991 10121
rect 9933 10112 9945 10115
rect 9824 10084 9945 10112
rect 9824 10072 9830 10084
rect 9933 10081 9945 10084
rect 9979 10081 9991 10115
rect 9933 10075 9991 10081
rect 10778 10072 10784 10124
rect 10836 10112 10842 10124
rect 11698 10112 11704 10124
rect 10836 10084 11704 10112
rect 10836 10072 10842 10084
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10112 11851 10115
rect 12250 10112 12256 10124
rect 11839 10084 12256 10112
rect 11839 10081 11851 10084
rect 11793 10075 11851 10081
rect 12250 10072 12256 10084
rect 12308 10072 12314 10124
rect 12342 10072 12348 10124
rect 12400 10112 12406 10124
rect 12719 10112 12747 10220
rect 13538 10208 13544 10220
rect 13596 10248 13602 10260
rect 13817 10251 13875 10257
rect 13817 10248 13829 10251
rect 13596 10220 13829 10248
rect 13596 10208 13602 10220
rect 13817 10217 13829 10220
rect 13863 10217 13875 10251
rect 13817 10211 13875 10217
rect 14829 10251 14887 10257
rect 14829 10217 14841 10251
rect 14875 10248 14887 10251
rect 15562 10248 15568 10260
rect 14875 10220 15568 10248
rect 14875 10217 14887 10220
rect 14829 10211 14887 10217
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 15746 10208 15752 10260
rect 15804 10248 15810 10260
rect 17678 10248 17684 10260
rect 15804 10220 17684 10248
rect 15804 10208 15810 10220
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 20070 10248 20076 10260
rect 18196 10220 20076 10248
rect 18196 10208 18202 10220
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 20346 10208 20352 10260
rect 20404 10248 20410 10260
rect 20441 10251 20499 10257
rect 20441 10248 20453 10251
rect 20404 10220 20453 10248
rect 20404 10208 20410 10220
rect 20441 10217 20453 10220
rect 20487 10217 20499 10251
rect 20441 10211 20499 10217
rect 12897 10183 12955 10189
rect 12897 10149 12909 10183
rect 12943 10180 12955 10183
rect 18601 10183 18659 10189
rect 12943 10152 18451 10180
rect 12943 10149 12955 10152
rect 12897 10143 12955 10149
rect 12400 10084 12747 10112
rect 12805 10115 12863 10121
rect 12400 10072 12406 10084
rect 12805 10081 12817 10115
rect 12851 10112 12863 10115
rect 13909 10115 13967 10121
rect 12851 10084 13308 10112
rect 12851 10081 12863 10084
rect 12805 10075 12863 10081
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 6178 10044 6184 10056
rect 6139 10016 6184 10044
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10013 6331 10047
rect 6546 10044 6552 10056
rect 6273 10007 6331 10013
rect 6380 10016 6552 10044
rect 5258 9936 5264 9988
rect 5316 9976 5322 9988
rect 6288 9976 6316 10007
rect 5316 9948 6316 9976
rect 5316 9936 5322 9948
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9908 2099 9911
rect 2314 9908 2320 9920
rect 2087 9880 2320 9908
rect 2087 9877 2099 9880
rect 2041 9871 2099 9877
rect 2314 9868 2320 9880
rect 2372 9868 2378 9920
rect 5442 9908 5448 9920
rect 5403 9880 5448 9908
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 5721 9911 5779 9917
rect 5721 9908 5733 9911
rect 5592 9880 5733 9908
rect 5592 9868 5598 9880
rect 5721 9877 5733 9880
rect 5767 9877 5779 9911
rect 5721 9871 5779 9877
rect 5902 9868 5908 9920
rect 5960 9908 5966 9920
rect 6380 9908 6408 10016
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 6914 10004 6920 10056
rect 6972 10044 6978 10056
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 6972 10016 7113 10044
rect 6972 10004 6978 10016
rect 7101 10013 7113 10016
rect 7147 10013 7159 10047
rect 8386 10044 8392 10056
rect 8347 10016 8392 10044
rect 7101 10007 7159 10013
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 9140 10016 9720 10044
rect 7282 9936 7288 9988
rect 7340 9976 7346 9988
rect 9140 9976 9168 10016
rect 9692 9988 9720 10016
rect 10870 10004 10876 10056
rect 10928 10044 10934 10056
rect 12069 10047 12127 10053
rect 10928 10016 12020 10044
rect 10928 10004 10934 10016
rect 7340 9948 9168 9976
rect 7340 9936 7346 9948
rect 9674 9936 9680 9988
rect 9732 9936 9738 9988
rect 11514 9976 11520 9988
rect 10980 9948 11520 9976
rect 6546 9908 6552 9920
rect 5960 9880 6408 9908
rect 6507 9880 6552 9908
rect 5960 9868 5966 9880
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 7374 9868 7380 9920
rect 7432 9908 7438 9920
rect 7561 9911 7619 9917
rect 7561 9908 7573 9911
rect 7432 9880 7573 9908
rect 7432 9868 7438 9880
rect 7561 9877 7573 9880
rect 7607 9877 7619 9911
rect 7742 9908 7748 9920
rect 7703 9880 7748 9908
rect 7561 9871 7619 9877
rect 7742 9868 7748 9880
rect 7800 9868 7806 9920
rect 8570 9868 8576 9920
rect 8628 9908 8634 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8628 9880 8769 9908
rect 8628 9868 8634 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 9306 9868 9312 9920
rect 9364 9908 9370 9920
rect 10980 9908 11008 9948
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 9364 9880 11008 9908
rect 11057 9911 11115 9917
rect 9364 9868 9370 9880
rect 11057 9877 11069 9911
rect 11103 9908 11115 9911
rect 11146 9908 11152 9920
rect 11103 9880 11152 9908
rect 11103 9877 11115 9880
rect 11057 9871 11115 9877
rect 11146 9868 11152 9880
rect 11204 9868 11210 9920
rect 11992 9908 12020 10016
rect 12069 10013 12081 10047
rect 12115 10013 12127 10047
rect 13081 10047 13139 10053
rect 13081 10044 13093 10047
rect 12069 10007 12127 10013
rect 13004 10016 13093 10044
rect 12084 9976 12112 10007
rect 13004 9988 13032 10016
rect 13081 10013 13093 10016
rect 13127 10013 13139 10047
rect 13081 10007 13139 10013
rect 12084 9948 12940 9976
rect 12066 9908 12072 9920
rect 11992 9880 12072 9908
rect 12066 9868 12072 9880
rect 12124 9868 12130 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12912 9908 12940 9948
rect 12986 9936 12992 9988
rect 13044 9936 13050 9988
rect 13280 9976 13308 10084
rect 13909 10081 13921 10115
rect 13955 10112 13967 10115
rect 14274 10112 14280 10124
rect 13955 10084 14280 10112
rect 13955 10081 13967 10084
rect 13909 10075 13967 10081
rect 14274 10072 14280 10084
rect 14332 10072 14338 10124
rect 14550 10072 14556 10124
rect 14608 10112 14614 10124
rect 14645 10115 14703 10121
rect 14645 10112 14657 10115
rect 14608 10084 14657 10112
rect 14608 10072 14614 10084
rect 14645 10081 14657 10084
rect 14691 10081 14703 10115
rect 14645 10075 14703 10081
rect 15378 10072 15384 10124
rect 15436 10112 15442 10124
rect 15556 10115 15614 10121
rect 15556 10112 15568 10115
rect 15436 10084 15568 10112
rect 15436 10072 15442 10084
rect 15556 10081 15568 10084
rect 15602 10112 15614 10115
rect 17402 10112 17408 10124
rect 15602 10084 17408 10112
rect 15602 10081 15614 10084
rect 15556 10075 15614 10081
rect 17402 10072 17408 10084
rect 17460 10112 17466 10124
rect 17586 10112 17592 10124
rect 17460 10084 17592 10112
rect 17460 10072 17466 10084
rect 17586 10072 17592 10084
rect 17644 10072 17650 10124
rect 17681 10115 17739 10121
rect 17681 10081 17693 10115
rect 17727 10081 17739 10115
rect 17681 10075 17739 10081
rect 17773 10115 17831 10121
rect 17773 10081 17785 10115
rect 17819 10112 17831 10115
rect 18138 10112 18144 10124
rect 17819 10084 18144 10112
rect 17819 10081 17831 10084
rect 17773 10075 17831 10081
rect 13357 10047 13415 10053
rect 13357 10013 13369 10047
rect 13403 10044 13415 10047
rect 14001 10047 14059 10053
rect 14001 10044 14013 10047
rect 13403 10016 14013 10044
rect 13403 10013 13415 10016
rect 13357 10007 13415 10013
rect 14001 10013 14013 10016
rect 14047 10044 14059 10047
rect 15102 10044 15108 10056
rect 14047 10016 15108 10044
rect 14047 10013 14059 10016
rect 14001 10007 14059 10013
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15289 10047 15347 10053
rect 15289 10044 15301 10047
rect 15252 10016 15301 10044
rect 15252 10004 15258 10016
rect 15289 10013 15301 10016
rect 15335 10013 15347 10047
rect 15289 10007 15347 10013
rect 16482 10004 16488 10056
rect 16540 10044 16546 10056
rect 16850 10044 16856 10056
rect 16540 10016 16856 10044
rect 16540 10004 16546 10016
rect 16850 10004 16856 10016
rect 16908 10004 16914 10056
rect 16942 10004 16948 10056
rect 17000 10044 17006 10056
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 17000 10016 17141 10044
rect 17000 10004 17006 10016
rect 17129 10013 17141 10016
rect 17175 10044 17187 10047
rect 17696 10044 17724 10075
rect 18138 10072 18144 10084
rect 18196 10072 18202 10124
rect 18335 10115 18393 10121
rect 18335 10081 18347 10115
rect 18381 10081 18393 10115
rect 18423 10112 18451 10152
rect 18601 10149 18613 10183
rect 18647 10180 18659 10183
rect 18690 10180 18696 10192
rect 18647 10152 18696 10180
rect 18647 10149 18659 10152
rect 18601 10143 18659 10149
rect 18690 10140 18696 10152
rect 18748 10140 18754 10192
rect 18782 10140 18788 10192
rect 18840 10180 18846 10192
rect 18969 10183 19027 10189
rect 18969 10180 18981 10183
rect 18840 10152 18981 10180
rect 18840 10140 18846 10152
rect 18969 10149 18981 10152
rect 19015 10149 19027 10183
rect 18969 10143 19027 10149
rect 20254 10140 20260 10192
rect 20312 10180 20318 10192
rect 20714 10180 20720 10192
rect 20312 10152 20720 10180
rect 20312 10140 20318 10152
rect 20714 10140 20720 10152
rect 20772 10140 20778 10192
rect 19150 10112 19156 10124
rect 18423 10084 19156 10112
rect 18335 10075 18393 10081
rect 17865 10047 17923 10053
rect 17865 10044 17877 10047
rect 17175 10016 17724 10044
rect 17788 10016 17877 10044
rect 17175 10013 17187 10016
rect 17129 10007 17187 10013
rect 17788 9988 17816 10016
rect 17865 10013 17877 10016
rect 17911 10013 17923 10047
rect 18347 10044 18375 10075
rect 19150 10072 19156 10084
rect 19208 10072 19214 10124
rect 19334 10121 19340 10124
rect 19328 10112 19340 10121
rect 19295 10084 19340 10112
rect 19328 10075 19340 10084
rect 19334 10072 19340 10075
rect 19392 10072 19398 10124
rect 18782 10044 18788 10056
rect 18347 10016 18788 10044
rect 17865 10007 17923 10013
rect 18782 10004 18788 10016
rect 18840 10004 18846 10056
rect 18969 10047 19027 10053
rect 18969 10013 18981 10047
rect 19015 10044 19027 10047
rect 19061 10047 19119 10053
rect 19061 10044 19073 10047
rect 19015 10016 19073 10044
rect 19015 10013 19027 10016
rect 18969 10007 19027 10013
rect 19061 10013 19073 10016
rect 19107 10013 19119 10047
rect 20898 10044 20904 10056
rect 20859 10016 20904 10044
rect 19061 10007 19119 10013
rect 20898 10004 20904 10016
rect 20956 10004 20962 10056
rect 13280 9948 15332 9976
rect 13357 9911 13415 9917
rect 13357 9908 13369 9911
rect 12492 9880 12537 9908
rect 12912 9880 13369 9908
rect 12492 9868 12498 9880
rect 13357 9877 13369 9880
rect 13403 9877 13415 9911
rect 13357 9871 13415 9877
rect 13449 9911 13507 9917
rect 13449 9877 13461 9911
rect 13495 9908 13507 9911
rect 13722 9908 13728 9920
rect 13495 9880 13728 9908
rect 13495 9877 13507 9880
rect 13449 9871 13507 9877
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 14090 9868 14096 9920
rect 14148 9908 14154 9920
rect 14366 9908 14372 9920
rect 14148 9880 14372 9908
rect 14148 9868 14154 9880
rect 14366 9868 14372 9880
rect 14424 9868 14430 9920
rect 15304 9908 15332 9948
rect 16408 9948 17724 9976
rect 16408 9908 16436 9948
rect 15304 9880 16436 9908
rect 16482 9868 16488 9920
rect 16540 9908 16546 9920
rect 16669 9911 16727 9917
rect 16669 9908 16681 9911
rect 16540 9880 16681 9908
rect 16540 9868 16546 9880
rect 16669 9877 16681 9880
rect 16715 9877 16727 9911
rect 16669 9871 16727 9877
rect 17126 9868 17132 9920
rect 17184 9908 17190 9920
rect 17313 9911 17371 9917
rect 17313 9908 17325 9911
rect 17184 9880 17325 9908
rect 17184 9868 17190 9880
rect 17313 9877 17325 9880
rect 17359 9877 17371 9911
rect 17696 9908 17724 9948
rect 17770 9936 17776 9988
rect 17828 9936 17834 9988
rect 17880 9948 19012 9976
rect 17880 9908 17908 9948
rect 18984 9920 19012 9948
rect 17696 9880 17908 9908
rect 17313 9871 17371 9877
rect 18966 9868 18972 9920
rect 19024 9868 19030 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 3145 9707 3203 9713
rect 3145 9704 3157 9707
rect 2556 9676 3157 9704
rect 2556 9664 2562 9676
rect 3145 9673 3157 9676
rect 3191 9673 3203 9707
rect 3145 9667 3203 9673
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 8754 9704 8760 9716
rect 5776 9676 8760 9704
rect 5776 9664 5782 9676
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 9217 9707 9275 9713
rect 9217 9673 9229 9707
rect 9263 9704 9275 9707
rect 9398 9704 9404 9716
rect 9263 9676 9404 9704
rect 9263 9673 9275 9676
rect 9217 9667 9275 9673
rect 9398 9664 9404 9676
rect 9456 9704 9462 9716
rect 9766 9704 9772 9716
rect 9456 9676 9772 9704
rect 9456 9664 9462 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 10410 9664 10416 9716
rect 10468 9704 10474 9716
rect 12342 9704 12348 9716
rect 10468 9676 12348 9704
rect 10468 9664 10474 9676
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 17586 9704 17592 9716
rect 13136 9676 16795 9704
rect 17547 9676 17592 9704
rect 13136 9664 13142 9676
rect 1765 9639 1823 9645
rect 1765 9605 1777 9639
rect 1811 9636 1823 9639
rect 3050 9636 3056 9648
rect 1811 9608 3056 9636
rect 1811 9605 1823 9608
rect 1765 9599 1823 9605
rect 3050 9596 3056 9608
rect 3108 9596 3114 9648
rect 3510 9596 3516 9648
rect 3568 9636 3574 9648
rect 3786 9636 3792 9648
rect 3568 9608 3792 9636
rect 3568 9596 3574 9608
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 4154 9636 4160 9648
rect 4115 9608 4160 9636
rect 4154 9596 4160 9608
rect 4212 9596 4218 9648
rect 5258 9636 5264 9648
rect 4264 9608 5264 9636
rect 4264 9580 4292 9608
rect 5258 9596 5264 9608
rect 5316 9636 5322 9648
rect 6362 9636 6368 9648
rect 5316 9608 5764 9636
rect 6323 9608 6368 9636
rect 5316 9596 5322 9608
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2464 9540 2697 9568
rect 2464 9528 2470 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9500 1639 9503
rect 1854 9500 1860 9512
rect 1627 9472 1860 9500
rect 1627 9469 1639 9472
rect 1581 9463 1639 9469
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 2700 9500 2728 9531
rect 3234 9528 3240 9580
rect 3292 9568 3298 9580
rect 3697 9571 3755 9577
rect 3697 9568 3709 9571
rect 3292 9540 3709 9568
rect 3292 9528 3298 9540
rect 3697 9537 3709 9540
rect 3743 9568 3755 9571
rect 4246 9568 4252 9580
rect 3743 9540 4252 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 4709 9571 4767 9577
rect 4709 9568 4721 9571
rect 4540 9540 4721 9568
rect 4540 9500 4568 9540
rect 4709 9537 4721 9540
rect 4755 9568 4767 9571
rect 5442 9568 5448 9580
rect 4755 9540 5448 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5736 9577 5764 9608
rect 6362 9596 6368 9608
rect 6420 9596 6426 9648
rect 6822 9636 6828 9648
rect 6783 9608 6828 9636
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 7190 9596 7196 9648
rect 7248 9636 7254 9648
rect 7650 9636 7656 9648
rect 7248 9608 7656 9636
rect 7248 9596 7254 9608
rect 7650 9596 7656 9608
rect 7708 9596 7714 9648
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 10870 9636 10876 9648
rect 9732 9608 10876 9636
rect 9732 9596 9738 9608
rect 10870 9596 10876 9608
rect 10928 9636 10934 9648
rect 11333 9639 11391 9645
rect 10928 9608 11100 9636
rect 10928 9596 10934 9608
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9568 5779 9571
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 5767 9540 7389 9568
rect 5767 9537 5779 9540
rect 5721 9531 5779 9537
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7558 9528 7564 9580
rect 7616 9568 7622 9580
rect 7616 9540 7880 9568
rect 7616 9528 7622 9540
rect 2700 9472 4568 9500
rect 4617 9503 4675 9509
rect 4617 9469 4629 9503
rect 4663 9500 4675 9503
rect 5534 9500 5540 9512
rect 4663 9472 5540 9500
rect 4663 9469 4675 9472
rect 4617 9463 4675 9469
rect 5534 9460 5540 9472
rect 5592 9460 5598 9512
rect 7852 9509 7880 9540
rect 8938 9528 8944 9580
rect 8996 9568 9002 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 8996 9540 10149 9568
rect 8996 9528 9002 9540
rect 10137 9537 10149 9540
rect 10183 9568 10195 9571
rect 10226 9568 10232 9580
rect 10183 9540 10232 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 10226 9528 10232 9540
rect 10284 9528 10290 9580
rect 11072 9577 11100 9608
rect 11333 9605 11345 9639
rect 11379 9636 11391 9639
rect 11379 9608 12480 9636
rect 11379 9605 11391 9608
rect 11333 9599 11391 9605
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9537 11115 9571
rect 11882 9568 11888 9580
rect 11843 9540 11888 9568
rect 11057 9531 11115 9537
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 12452 9568 12480 9608
rect 13814 9596 13820 9648
rect 13872 9636 13878 9648
rect 14369 9639 14427 9645
rect 13872 9608 14320 9636
rect 13872 9596 13878 9608
rect 12452 9540 12572 9568
rect 12544 9512 12572 9540
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9500 6239 9503
rect 7837 9503 7895 9509
rect 6227 9472 7788 9500
rect 6227 9469 6239 9472
rect 6181 9463 6239 9469
rect 2590 9432 2596 9444
rect 2551 9404 2596 9432
rect 2590 9392 2596 9404
rect 2648 9392 2654 9444
rect 3878 9432 3884 9444
rect 3528 9404 3884 9432
rect 2133 9367 2191 9373
rect 2133 9333 2145 9367
rect 2179 9364 2191 9367
rect 2406 9364 2412 9376
rect 2179 9336 2412 9364
rect 2179 9333 2191 9336
rect 2133 9327 2191 9333
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 2498 9324 2504 9376
rect 2556 9364 2562 9376
rect 2556 9336 2601 9364
rect 2556 9324 2562 9336
rect 2958 9324 2964 9376
rect 3016 9364 3022 9376
rect 3528 9373 3556 9404
rect 3878 9392 3884 9404
rect 3936 9392 3942 9444
rect 4525 9435 4583 9441
rect 4525 9401 4537 9435
rect 4571 9432 4583 9435
rect 4571 9404 5212 9432
rect 4571 9401 4583 9404
rect 4525 9395 4583 9401
rect 3513 9367 3571 9373
rect 3513 9364 3525 9367
rect 3016 9336 3525 9364
rect 3016 9324 3022 9336
rect 3513 9333 3525 9336
rect 3559 9333 3571 9367
rect 3513 9327 3571 9333
rect 3605 9367 3663 9373
rect 3605 9333 3617 9367
rect 3651 9364 3663 9367
rect 3694 9364 3700 9376
rect 3651 9336 3700 9364
rect 3651 9333 3663 9336
rect 3605 9327 3663 9333
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 5184 9373 5212 9404
rect 5718 9392 5724 9444
rect 5776 9432 5782 9444
rect 7285 9435 7343 9441
rect 7285 9432 7297 9435
rect 5776 9404 7297 9432
rect 5776 9392 5782 9404
rect 7285 9401 7297 9404
rect 7331 9401 7343 9435
rect 7760 9432 7788 9472
rect 7837 9469 7849 9503
rect 7883 9500 7895 9503
rect 9490 9500 9496 9512
rect 7883 9472 9496 9500
rect 7883 9469 7895 9472
rect 7837 9463 7895 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9500 9919 9503
rect 9907 9472 12204 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 7926 9432 7932 9444
rect 7760 9404 7932 9432
rect 7285 9395 7343 9401
rect 7926 9392 7932 9404
rect 7984 9392 7990 9444
rect 8104 9435 8162 9441
rect 8104 9401 8116 9435
rect 8150 9432 8162 9435
rect 8754 9432 8760 9444
rect 8150 9404 8760 9432
rect 8150 9401 8162 9404
rect 8104 9395 8162 9401
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 8846 9392 8852 9444
rect 8904 9432 8910 9444
rect 8904 9404 10548 9432
rect 8904 9392 8910 9404
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9333 5227 9367
rect 5169 9327 5227 9333
rect 5258 9324 5264 9376
rect 5316 9364 5322 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 5316 9336 5549 9364
rect 5316 9324 5322 9336
rect 5537 9333 5549 9336
rect 5583 9333 5595 9367
rect 5537 9327 5595 9333
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 5902 9364 5908 9376
rect 5684 9336 5908 9364
rect 5684 9324 5690 9336
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 7193 9367 7251 9373
rect 7193 9333 7205 9367
rect 7239 9364 7251 9367
rect 9306 9364 9312 9376
rect 7239 9336 9312 9364
rect 7239 9333 7251 9336
rect 7193 9327 7251 9333
rect 9306 9324 9312 9336
rect 9364 9324 9370 9376
rect 9490 9364 9496 9376
rect 9451 9336 9496 9364
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 9950 9364 9956 9376
rect 9911 9336 9956 9364
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 10520 9373 10548 9404
rect 10962 9392 10968 9444
rect 11020 9432 11026 9444
rect 11514 9432 11520 9444
rect 11020 9404 11520 9432
rect 11020 9392 11026 9404
rect 11514 9392 11520 9404
rect 11572 9392 11578 9444
rect 11698 9432 11704 9444
rect 11659 9404 11704 9432
rect 11698 9392 11704 9404
rect 11756 9392 11762 9444
rect 11790 9392 11796 9444
rect 11848 9432 11854 9444
rect 12176 9432 12204 9472
rect 12342 9460 12348 9512
rect 12400 9500 12406 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12400 9472 12449 9500
rect 12400 9460 12406 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 12526 9460 12532 9512
rect 12584 9460 12590 9512
rect 14090 9500 14096 9512
rect 12636 9472 14096 9500
rect 12636 9432 12664 9472
rect 14090 9460 14096 9472
rect 14148 9460 14154 9512
rect 14292 9509 14320 9608
rect 14369 9605 14381 9639
rect 14415 9605 14427 9639
rect 14369 9599 14427 9605
rect 14384 9568 14412 9599
rect 14458 9596 14464 9648
rect 14516 9636 14522 9648
rect 14516 9608 15056 9636
rect 14516 9596 14522 9608
rect 14918 9568 14924 9580
rect 14384 9540 14495 9568
rect 14879 9540 14924 9568
rect 14269 9503 14327 9509
rect 14269 9469 14281 9503
rect 14315 9469 14327 9503
rect 14269 9463 14327 9469
rect 14366 9460 14372 9512
rect 14424 9500 14430 9512
rect 14467 9500 14495 9540
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 15028 9568 15056 9608
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 15746 9636 15752 9648
rect 15252 9608 15752 9636
rect 15252 9596 15258 9608
rect 15746 9596 15752 9608
rect 15804 9596 15810 9648
rect 16767 9568 16795 9676
rect 17586 9664 17592 9676
rect 17644 9664 17650 9716
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18049 9707 18107 9713
rect 18049 9704 18061 9707
rect 18012 9676 18061 9704
rect 18012 9664 18018 9676
rect 18049 9673 18061 9676
rect 18095 9673 18107 9707
rect 20714 9704 20720 9716
rect 18049 9667 18107 9673
rect 18156 9676 20720 9704
rect 17126 9636 17132 9648
rect 17087 9608 17132 9636
rect 17126 9596 17132 9608
rect 17184 9596 17190 9648
rect 17313 9639 17371 9645
rect 17313 9605 17325 9639
rect 17359 9636 17371 9639
rect 18156 9636 18184 9676
rect 20714 9664 20720 9676
rect 20772 9664 20778 9716
rect 17359 9608 18184 9636
rect 17359 9605 17371 9608
rect 17313 9599 17371 9605
rect 19058 9596 19064 9648
rect 19116 9636 19122 9648
rect 19116 9608 19161 9636
rect 19116 9596 19122 9608
rect 19242 9596 19248 9648
rect 19300 9636 19306 9648
rect 20073 9639 20131 9645
rect 20073 9636 20085 9639
rect 19300 9608 20085 9636
rect 19300 9596 19306 9608
rect 20073 9605 20085 9608
rect 20119 9605 20131 9639
rect 20073 9599 20131 9605
rect 17770 9568 17776 9580
rect 15028 9540 15884 9568
rect 16767 9540 17776 9568
rect 15562 9500 15568 9512
rect 14424 9472 14495 9500
rect 14660 9472 15568 9500
rect 14424 9460 14430 9472
rect 11848 9404 11893 9432
rect 12176 9404 12664 9432
rect 12704 9435 12762 9441
rect 11848 9392 11854 9404
rect 12704 9401 12716 9435
rect 12750 9432 12762 9435
rect 12802 9432 12808 9444
rect 12750 9404 12808 9432
rect 12750 9401 12762 9404
rect 12704 9395 12762 9401
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 14660 9432 14688 9472
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 15746 9500 15752 9512
rect 15707 9472 15752 9500
rect 15746 9460 15752 9472
rect 15804 9460 15810 9512
rect 15856 9500 15884 9540
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 17862 9528 17868 9580
rect 17920 9568 17926 9580
rect 18601 9571 18659 9577
rect 18601 9568 18613 9571
rect 17920 9540 18613 9568
rect 17920 9528 17926 9540
rect 18601 9537 18613 9540
rect 18647 9537 18659 9571
rect 19610 9568 19616 9580
rect 18601 9531 18659 9537
rect 19067 9540 19616 9568
rect 17313 9503 17371 9509
rect 17313 9500 17325 9503
rect 15856 9472 17325 9500
rect 17313 9469 17325 9472
rect 17359 9469 17371 9503
rect 17313 9463 17371 9469
rect 17405 9503 17463 9509
rect 17405 9469 17417 9503
rect 17451 9500 17463 9503
rect 17494 9500 17500 9512
rect 17451 9472 17500 9500
rect 17451 9469 17463 9472
rect 17405 9463 17463 9469
rect 17494 9460 17500 9472
rect 17552 9460 17558 9512
rect 18417 9503 18475 9509
rect 18417 9469 18429 9503
rect 18463 9500 18475 9503
rect 19067 9500 19095 9540
rect 19610 9528 19616 9540
rect 19668 9528 19674 9580
rect 19702 9528 19708 9580
rect 19760 9568 19766 9580
rect 19981 9571 20039 9577
rect 19760 9540 19805 9568
rect 19760 9528 19766 9540
rect 19981 9537 19993 9571
rect 20027 9568 20039 9571
rect 20625 9571 20683 9577
rect 20625 9568 20637 9571
rect 20027 9540 20637 9568
rect 20027 9537 20039 9540
rect 19981 9531 20039 9537
rect 20625 9537 20637 9540
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 19150 9500 19156 9512
rect 18463 9472 19156 9500
rect 18463 9469 18475 9472
rect 18417 9463 18475 9469
rect 19150 9460 19156 9472
rect 19208 9460 19214 9512
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9500 19487 9503
rect 19475 9472 19748 9500
rect 19475 9469 19487 9472
rect 19429 9463 19487 9469
rect 12912 9404 14688 9432
rect 14737 9435 14795 9441
rect 10505 9367 10563 9373
rect 10505 9333 10517 9367
rect 10551 9333 10563 9367
rect 10505 9327 10563 9333
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 10873 9367 10931 9373
rect 10873 9364 10885 9367
rect 10744 9336 10885 9364
rect 10744 9324 10750 9336
rect 10873 9333 10885 9336
rect 10919 9333 10931 9367
rect 10873 9327 10931 9333
rect 11974 9324 11980 9376
rect 12032 9364 12038 9376
rect 12912 9364 12940 9404
rect 14737 9401 14749 9435
rect 14783 9432 14795 9435
rect 15286 9432 15292 9444
rect 14783 9404 15292 9432
rect 14783 9401 14795 9404
rect 14737 9395 14795 9401
rect 15286 9392 15292 9404
rect 15344 9392 15350 9444
rect 16016 9435 16074 9441
rect 16016 9401 16028 9435
rect 16062 9432 16074 9435
rect 16482 9432 16488 9444
rect 16062 9404 16488 9432
rect 16062 9401 16074 9404
rect 16016 9395 16074 9401
rect 16482 9392 16488 9404
rect 16540 9392 16546 9444
rect 16666 9392 16672 9444
rect 16724 9432 16730 9444
rect 17586 9432 17592 9444
rect 16724 9404 17592 9432
rect 16724 9392 16730 9404
rect 17586 9392 17592 9404
rect 17644 9432 17650 9444
rect 18509 9435 18567 9441
rect 18509 9432 18521 9435
rect 17644 9404 18521 9432
rect 17644 9392 17650 9404
rect 18509 9401 18521 9404
rect 18555 9432 18567 9435
rect 18555 9404 19196 9432
rect 18555 9401 18567 9404
rect 18509 9395 18567 9401
rect 12032 9336 12940 9364
rect 12032 9324 12038 9336
rect 12986 9324 12992 9376
rect 13044 9364 13050 9376
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 13044 9336 13829 9364
rect 13044 9324 13050 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 14090 9364 14096 9376
rect 14051 9336 14096 9364
rect 13817 9327 13875 9333
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14829 9367 14887 9373
rect 14829 9333 14841 9367
rect 14875 9364 14887 9367
rect 16298 9364 16304 9376
rect 14875 9336 16304 9364
rect 14875 9333 14887 9336
rect 14829 9327 14887 9333
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 19168 9364 19196 9404
rect 19242 9392 19248 9444
rect 19300 9432 19306 9444
rect 19610 9432 19616 9444
rect 19300 9404 19616 9432
rect 19300 9392 19306 9404
rect 19610 9392 19616 9404
rect 19668 9392 19674 9444
rect 19720 9432 19748 9472
rect 19794 9460 19800 9512
rect 19852 9500 19858 9512
rect 20441 9503 20499 9509
rect 20441 9500 20453 9503
rect 19852 9472 20453 9500
rect 19852 9460 19858 9472
rect 20441 9469 20453 9472
rect 20487 9469 20499 9503
rect 20441 9463 20499 9469
rect 20898 9432 20904 9444
rect 19720 9404 20904 9432
rect 20898 9392 20904 9404
rect 20956 9392 20962 9444
rect 19426 9364 19432 9376
rect 19168 9336 19432 9364
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 19521 9367 19579 9373
rect 19521 9333 19533 9367
rect 19567 9364 19579 9367
rect 19702 9364 19708 9376
rect 19567 9336 19708 9364
rect 19567 9333 19579 9336
rect 19521 9327 19579 9333
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 19794 9324 19800 9376
rect 19852 9364 19858 9376
rect 19981 9367 20039 9373
rect 19981 9364 19993 9367
rect 19852 9336 19993 9364
rect 19852 9324 19858 9336
rect 19981 9333 19993 9336
rect 20027 9333 20039 9367
rect 20530 9364 20536 9376
rect 20491 9336 20536 9364
rect 19981 9327 20039 9333
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2222 9160 2228 9172
rect 1995 9132 2228 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 2406 9160 2412 9172
rect 2367 9132 2412 9160
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 2590 9120 2596 9172
rect 2648 9160 2654 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 2648 9132 4077 9160
rect 2648 9120 2654 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 7009 9163 7067 9169
rect 4764 9132 6592 9160
rect 4764 9120 4770 9132
rect 2314 9092 2320 9104
rect 2275 9064 2320 9092
rect 2314 9052 2320 9064
rect 2372 9052 2378 9104
rect 3326 9092 3332 9104
rect 3287 9064 3332 9092
rect 3326 9052 3332 9064
rect 3384 9052 3390 9104
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 5534 9092 5540 9104
rect 4212 9064 5540 9092
rect 4212 9052 4218 9064
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 2406 8984 2412 9036
rect 2464 9024 2470 9036
rect 2958 9024 2964 9036
rect 2464 8996 2964 9024
rect 2464 8984 2470 8996
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 3050 8984 3056 9036
rect 3108 9024 3114 9036
rect 4433 9027 4491 9033
rect 3108 8996 3648 9024
rect 3108 8984 3114 8996
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 2682 8956 2688 8968
rect 2639 8928 2688 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 3421 8959 3479 8965
rect 3421 8956 3433 8959
rect 3252 8928 3433 8956
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 3142 8888 3148 8900
rect 1627 8860 3148 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 3252 8832 3280 8928
rect 3421 8925 3433 8928
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8925 3571 8959
rect 3620 8956 3648 8996
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4890 9024 4896 9036
rect 4479 8996 4896 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 5092 9033 5120 9064
rect 5534 9052 5540 9064
rect 5592 9052 5598 9104
rect 5350 9033 5356 9036
rect 5077 9027 5135 9033
rect 5077 8993 5089 9027
rect 5123 8993 5135 9027
rect 5077 8987 5135 8993
rect 5344 8987 5356 9033
rect 5408 9024 5414 9036
rect 5408 8996 5444 9024
rect 5350 8984 5356 8987
rect 5408 8984 5414 8996
rect 4525 8959 4583 8965
rect 4525 8956 4537 8959
rect 3620 8928 4537 8956
rect 3513 8919 3571 8925
rect 4525 8925 4537 8928
rect 4571 8925 4583 8959
rect 4525 8919 4583 8925
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 3326 8848 3332 8900
rect 3384 8888 3390 8900
rect 3528 8888 3556 8919
rect 4632 8888 4660 8919
rect 3384 8860 4660 8888
rect 3384 8848 3390 8860
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 2961 8823 3019 8829
rect 2961 8820 2973 8823
rect 2832 8792 2973 8820
rect 2832 8780 2838 8792
rect 2961 8789 2973 8792
rect 3007 8789 3019 8823
rect 2961 8783 3019 8789
rect 3234 8780 3240 8832
rect 3292 8780 3298 8832
rect 4632 8820 4660 8860
rect 6457 8823 6515 8829
rect 6457 8820 6469 8823
rect 4632 8792 6469 8820
rect 6457 8789 6469 8792
rect 6503 8789 6515 8823
rect 6564 8820 6592 9132
rect 7009 9129 7021 9163
rect 7055 9160 7067 9163
rect 8202 9160 8208 9172
rect 7055 9132 8208 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 8754 9160 8760 9172
rect 8715 9132 8760 9160
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 9214 9160 9220 9172
rect 9175 9132 9220 9160
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 9548 9132 10057 9160
rect 9548 9120 9554 9132
rect 10045 9129 10057 9132
rect 10091 9129 10103 9163
rect 10045 9123 10103 9129
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10318 9160 10324 9172
rect 10192 9132 10324 9160
rect 10192 9120 10198 9132
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 10502 9120 10508 9172
rect 10560 9160 10566 9172
rect 10686 9160 10692 9172
rect 10560 9132 10692 9160
rect 10560 9120 10566 9132
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 12342 9160 12348 9172
rect 10836 9132 12348 9160
rect 10836 9120 10842 9132
rect 12342 9120 12348 9132
rect 12400 9160 12406 9172
rect 12894 9160 12900 9172
rect 12400 9132 12900 9160
rect 12400 9120 12406 9132
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 12989 9163 13047 9169
rect 12989 9129 13001 9163
rect 13035 9160 13047 9163
rect 13446 9160 13452 9172
rect 13035 9132 13452 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 13541 9163 13599 9169
rect 13541 9129 13553 9163
rect 13587 9160 13599 9163
rect 13906 9160 13912 9172
rect 13587 9132 13912 9160
rect 13587 9129 13599 9132
rect 13541 9123 13599 9129
rect 13906 9120 13912 9132
rect 13964 9120 13970 9172
rect 14182 9120 14188 9172
rect 14240 9160 14246 9172
rect 14829 9163 14887 9169
rect 14829 9160 14841 9163
rect 14240 9132 14841 9160
rect 14240 9120 14246 9132
rect 14829 9129 14841 9132
rect 14875 9129 14887 9163
rect 15286 9160 15292 9172
rect 15247 9132 15292 9160
rect 14829 9123 14887 9129
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15654 9160 15660 9172
rect 15488 9132 15660 9160
rect 7558 9092 7564 9104
rect 7392 9064 7564 9092
rect 6822 9024 6828 9036
rect 6783 8996 6828 9024
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7392 9033 7420 9064
rect 7558 9052 7564 9064
rect 7616 9092 7622 9104
rect 8110 9092 8116 9104
rect 7616 9064 8116 9092
rect 7616 9052 7622 9064
rect 8110 9052 8116 9064
rect 8168 9052 8174 9104
rect 8772 9092 8800 9120
rect 12066 9092 12072 9104
rect 8772 9064 10079 9092
rect 7650 9033 7656 9036
rect 7377 9027 7435 9033
rect 7377 8993 7389 9027
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 7644 8987 7656 9033
rect 7708 9024 7714 9036
rect 8938 9024 8944 9036
rect 7708 8996 8944 9024
rect 6822 8848 6828 8900
rect 6880 8888 6886 8900
rect 7392 8888 7420 8987
rect 7650 8984 7656 8987
rect 7708 8984 7714 8996
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 9033 9027 9091 9033
rect 9033 8993 9045 9027
rect 9079 8993 9091 9027
rect 9033 8987 9091 8993
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 9048 8956 9076 8987
rect 9306 8984 9312 9036
rect 9364 9024 9370 9036
rect 9401 9027 9459 9033
rect 9401 9024 9413 9027
rect 9364 8996 9413 9024
rect 9364 8984 9370 8996
rect 9401 8993 9413 8996
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 9950 8984 9956 9036
rect 10008 8984 10014 9036
rect 9766 8956 9772 8968
rect 8812 8928 9076 8956
rect 9140 8928 9772 8956
rect 8812 8916 8818 8928
rect 6880 8860 7420 8888
rect 6880 8848 6886 8860
rect 8386 8848 8392 8900
rect 8444 8888 8450 8900
rect 9140 8888 9168 8928
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 9968 8888 9996 8984
rect 10051 8956 10079 9064
rect 10612 9064 12072 9092
rect 10612 9033 10640 9064
rect 12066 9052 12072 9064
rect 12124 9052 12130 9104
rect 12434 9052 12440 9104
rect 12492 9092 12498 9104
rect 13081 9095 13139 9101
rect 13081 9092 13093 9095
rect 12492 9064 13093 9092
rect 12492 9052 12498 9064
rect 13081 9061 13093 9064
rect 13127 9061 13139 9095
rect 13081 9055 13139 9061
rect 13170 9052 13176 9104
rect 13228 9092 13234 9104
rect 14001 9095 14059 9101
rect 13228 9064 13952 9092
rect 13228 9052 13234 9064
rect 10137 9027 10195 9033
rect 10137 8993 10149 9027
rect 10183 9024 10195 9027
rect 10597 9027 10655 9033
rect 10183 8996 10550 9024
rect 10183 8993 10195 8996
rect 10137 8987 10195 8993
rect 10226 8956 10232 8968
rect 10051 8928 10232 8956
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 8444 8860 9168 8888
rect 9324 8860 9996 8888
rect 10522 8888 10550 8996
rect 10597 8993 10609 9027
rect 10643 8993 10655 9027
rect 10597 8987 10655 8993
rect 11232 9027 11290 9033
rect 11232 8993 11244 9027
rect 11278 9024 11290 9027
rect 12986 9024 12992 9036
rect 11278 8996 12992 9024
rect 11278 8993 11290 8996
rect 11232 8987 11290 8993
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 10778 8916 10784 8968
rect 10836 8956 10842 8968
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10836 8928 10977 8956
rect 10836 8916 10842 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 13078 8956 13084 8968
rect 12584 8928 13084 8956
rect 12584 8916 12590 8928
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 13188 8888 13216 8919
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 13814 8956 13820 8968
rect 13688 8928 13820 8956
rect 13688 8916 13694 8928
rect 13814 8916 13820 8928
rect 13872 8916 13878 8968
rect 10522 8860 11008 8888
rect 8444 8848 8450 8860
rect 9324 8820 9352 8860
rect 10980 8832 11008 8860
rect 12360 8860 13216 8888
rect 12360 8832 12388 8860
rect 6564 8792 9352 8820
rect 9401 8823 9459 8829
rect 6457 8783 6515 8789
rect 9401 8789 9413 8823
rect 9447 8820 9459 8823
rect 9677 8823 9735 8829
rect 9677 8820 9689 8823
rect 9447 8792 9689 8820
rect 9447 8789 9459 8792
rect 9401 8783 9459 8789
rect 9677 8789 9689 8792
rect 9723 8789 9735 8823
rect 10778 8820 10784 8832
rect 10739 8792 10784 8820
rect 9677 8783 9735 8789
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 10962 8780 10968 8832
rect 11020 8780 11026 8832
rect 12342 8820 12348 8832
rect 12303 8792 12348 8820
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 12621 8823 12679 8829
rect 12621 8789 12633 8823
rect 12667 8820 12679 8823
rect 12710 8820 12716 8832
rect 12667 8792 12716 8820
rect 12667 8789 12679 8792
rect 12621 8783 12679 8789
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 13538 8820 13544 8832
rect 13499 8792 13544 8820
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 13633 8823 13691 8829
rect 13633 8789 13645 8823
rect 13679 8820 13691 8823
rect 13814 8820 13820 8832
rect 13679 8792 13820 8820
rect 13679 8789 13691 8792
rect 13633 8783 13691 8789
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 13924 8820 13952 9064
rect 14001 9061 14013 9095
rect 14047 9092 14059 9095
rect 15194 9092 15200 9104
rect 14047 9064 15200 9092
rect 14047 9061 14059 9064
rect 14001 9055 14059 9061
rect 15194 9052 15200 9064
rect 15252 9052 15258 9104
rect 14642 8984 14648 9036
rect 14700 9024 14706 9036
rect 14700 8996 14745 9024
rect 14700 8984 14706 8996
rect 15286 8984 15292 9036
rect 15344 9024 15350 9036
rect 15488 9024 15516 9132
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 16298 9160 16304 9172
rect 16259 9132 16304 9160
rect 16298 9120 16304 9132
rect 16356 9120 16362 9172
rect 16390 9120 16396 9172
rect 16448 9160 16454 9172
rect 17221 9163 17279 9169
rect 17221 9160 17233 9163
rect 16448 9132 17233 9160
rect 16448 9120 16454 9132
rect 17221 9129 17233 9132
rect 17267 9129 17279 9163
rect 17221 9123 17279 9129
rect 17402 9120 17408 9172
rect 17460 9160 17466 9172
rect 18141 9163 18199 9169
rect 18141 9160 18153 9163
rect 17460 9132 18153 9160
rect 17460 9120 17466 9132
rect 18141 9129 18153 9132
rect 18187 9160 18199 9163
rect 19242 9160 19248 9172
rect 18187 9132 19248 9160
rect 18187 9129 18199 9132
rect 18141 9123 18199 9129
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 19334 9120 19340 9172
rect 19392 9160 19398 9172
rect 19705 9163 19763 9169
rect 19705 9160 19717 9163
rect 19392 9132 19717 9160
rect 19392 9120 19398 9132
rect 19705 9129 19717 9132
rect 19751 9129 19763 9163
rect 19705 9123 19763 9129
rect 20714 9120 20720 9172
rect 20772 9160 20778 9172
rect 20901 9163 20959 9169
rect 20901 9160 20913 9163
rect 20772 9132 20913 9160
rect 20772 9120 20778 9132
rect 20901 9129 20913 9132
rect 20947 9129 20959 9163
rect 20901 9123 20959 9129
rect 15562 9052 15568 9104
rect 15620 9092 15626 9104
rect 20257 9095 20315 9101
rect 20257 9092 20269 9095
rect 15620 9064 18828 9092
rect 15620 9052 15626 9064
rect 15654 9024 15660 9036
rect 15344 8996 15516 9024
rect 15615 8996 15660 9024
rect 15344 8984 15350 8996
rect 15654 8984 15660 8996
rect 15712 8984 15718 9036
rect 15749 9027 15807 9033
rect 15749 8993 15761 9027
rect 15795 9024 15807 9027
rect 15930 9024 15936 9036
rect 15795 8996 15936 9024
rect 15795 8993 15807 8996
rect 15749 8987 15807 8993
rect 15930 8984 15936 8996
rect 15988 9024 15994 9036
rect 16390 9024 16396 9036
rect 15988 8996 16396 9024
rect 15988 8984 15994 8996
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 16669 9027 16727 9033
rect 16669 9024 16681 9027
rect 16632 8996 16681 9024
rect 16632 8984 16638 8996
rect 16669 8993 16681 8996
rect 16715 8993 16727 9027
rect 16669 8987 16727 8993
rect 16761 9027 16819 9033
rect 16761 8993 16773 9027
rect 16807 9024 16819 9027
rect 16942 9024 16948 9036
rect 16807 8996 16948 9024
rect 16807 8993 16819 8996
rect 16761 8987 16819 8993
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17586 8984 17592 9036
rect 17644 9024 17650 9036
rect 17681 9027 17739 9033
rect 17681 9024 17693 9027
rect 17644 8996 17693 9024
rect 17644 8984 17650 8996
rect 17681 8993 17693 8996
rect 17727 8993 17739 9027
rect 17681 8987 17739 8993
rect 17770 8984 17776 9036
rect 17828 9024 17834 9036
rect 17828 8996 17873 9024
rect 17828 8984 17834 8996
rect 18046 8984 18052 9036
rect 18104 9024 18110 9036
rect 18598 9033 18604 9036
rect 18325 9027 18383 9033
rect 18325 9024 18337 9027
rect 18104 8996 18337 9024
rect 18104 8984 18110 8996
rect 18325 8993 18337 8996
rect 18371 8993 18383 9027
rect 18592 9024 18604 9033
rect 18559 8996 18604 9024
rect 18325 8987 18383 8993
rect 18592 8987 18604 8996
rect 18598 8984 18604 8987
rect 18656 8984 18662 9036
rect 18800 9024 18828 9064
rect 18984 9064 20269 9092
rect 18984 9024 19012 9064
rect 20257 9061 20269 9064
rect 20303 9061 20315 9095
rect 20257 9055 20315 9061
rect 19978 9024 19984 9036
rect 18800 8996 19012 9024
rect 19939 8996 19984 9024
rect 19978 8984 19984 8996
rect 20036 8984 20042 9036
rect 14093 8959 14151 8965
rect 14093 8925 14105 8959
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8956 14335 8959
rect 14734 8956 14740 8968
rect 14323 8928 14740 8956
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 14108 8888 14136 8919
rect 14734 8916 14740 8928
rect 14792 8916 14798 8968
rect 14826 8916 14832 8968
rect 14884 8956 14890 8968
rect 15013 8959 15071 8965
rect 15013 8956 15025 8959
rect 14884 8928 15025 8956
rect 14884 8916 14890 8928
rect 15013 8925 15025 8928
rect 15059 8925 15071 8959
rect 15013 8919 15071 8925
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 15160 8928 15853 8956
rect 15160 8916 15166 8928
rect 15841 8925 15853 8928
rect 15887 8956 15899 8959
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 15887 8928 16865 8956
rect 15887 8925 15899 8928
rect 15841 8919 15899 8925
rect 16853 8925 16865 8928
rect 16899 8956 16911 8959
rect 17034 8956 17040 8968
rect 16899 8928 17040 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 17034 8916 17040 8928
rect 17092 8916 17098 8968
rect 17954 8916 17960 8968
rect 18012 8956 18018 8968
rect 18141 8959 18199 8965
rect 18141 8956 18153 8959
rect 18012 8928 18153 8956
rect 18012 8916 18018 8928
rect 18141 8925 18153 8928
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 19886 8956 19892 8968
rect 19392 8928 19892 8956
rect 19392 8916 19398 8928
rect 19886 8916 19892 8928
rect 19944 8916 19950 8968
rect 16390 8888 16396 8900
rect 14108 8860 14780 8888
rect 14090 8820 14096 8832
rect 13924 8792 14096 8820
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 14274 8780 14280 8832
rect 14332 8820 14338 8832
rect 14642 8820 14648 8832
rect 14332 8792 14648 8820
rect 14332 8780 14338 8792
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 14752 8820 14780 8860
rect 14936 8860 16396 8888
rect 14936 8820 14964 8860
rect 16390 8848 16396 8860
rect 16448 8848 16454 8900
rect 17221 8891 17279 8897
rect 17221 8857 17233 8891
rect 17267 8888 17279 8891
rect 17267 8860 17724 8888
rect 17267 8857 17279 8860
rect 17221 8851 17279 8857
rect 14752 8792 14964 8820
rect 15013 8823 15071 8829
rect 15013 8789 15025 8823
rect 15059 8820 15071 8823
rect 15562 8820 15568 8832
rect 15059 8792 15568 8820
rect 15059 8789 15071 8792
rect 15013 8783 15071 8789
rect 15562 8780 15568 8792
rect 15620 8780 15626 8832
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 17313 8823 17371 8829
rect 17313 8820 17325 8823
rect 16724 8792 17325 8820
rect 16724 8780 16730 8792
rect 17313 8789 17325 8792
rect 17359 8789 17371 8823
rect 17696 8820 17724 8860
rect 19426 8848 19432 8900
rect 19484 8888 19490 8900
rect 19610 8888 19616 8900
rect 19484 8860 19616 8888
rect 19484 8848 19490 8860
rect 19610 8848 19616 8860
rect 19668 8848 19674 8900
rect 19794 8820 19800 8832
rect 17696 8792 19800 8820
rect 17313 8783 17371 8789
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 19978 8780 19984 8832
rect 20036 8820 20042 8832
rect 21266 8820 21272 8832
rect 20036 8792 21272 8820
rect 20036 8780 20042 8792
rect 21266 8780 21272 8792
rect 21324 8780 21330 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2409 8619 2467 8625
rect 2409 8585 2421 8619
rect 2455 8616 2467 8619
rect 2498 8616 2504 8628
rect 2455 8588 2504 8616
rect 2455 8585 2467 8588
rect 2409 8579 2467 8585
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 3602 8616 3608 8628
rect 3563 8588 3608 8616
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 5350 8616 5356 8628
rect 5311 8588 5356 8616
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 5718 8616 5724 8628
rect 5679 8588 5724 8616
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 6104 8588 6561 8616
rect 3234 8548 3240 8560
rect 1872 8520 3240 8548
rect 1872 8489 1900 8520
rect 3234 8508 3240 8520
rect 3292 8508 3298 8560
rect 5368 8548 5396 8576
rect 6104 8548 6132 8588
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 8389 8619 8447 8625
rect 8389 8616 8401 8619
rect 6549 8579 6607 8585
rect 6656 8588 8401 8616
rect 5368 8520 6132 8548
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8449 1915 8483
rect 2038 8480 2044 8492
rect 1951 8452 2044 8480
rect 1857 8443 1915 8449
rect 2038 8440 2044 8452
rect 2096 8480 2102 8492
rect 2866 8480 2872 8492
rect 2096 8452 2728 8480
rect 2827 8452 2872 8480
rect 2096 8440 2102 8452
rect 1762 8344 1768 8356
rect 1723 8316 1768 8344
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 1394 8276 1400 8288
rect 1355 8248 1400 8276
rect 1394 8236 1400 8248
rect 1452 8236 1458 8288
rect 2700 8276 2728 8452
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3326 8480 3332 8492
rect 3099 8452 3332 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 3970 8480 3976 8492
rect 3931 8452 3976 8480
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 6181 8483 6239 8489
rect 6181 8480 6193 8483
rect 5684 8452 6193 8480
rect 5684 8440 5690 8452
rect 6181 8449 6193 8452
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8480 6423 8483
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6411 8452 6561 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 3418 8412 3424 8424
rect 3379 8384 3424 8412
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 6656 8412 6684 8588
rect 8389 8585 8401 8588
rect 8435 8585 8447 8619
rect 9306 8616 9312 8628
rect 9267 8588 9312 8616
rect 8389 8579 8447 8585
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 10505 8619 10563 8625
rect 10505 8585 10517 8619
rect 10551 8616 10563 8619
rect 10962 8616 10968 8628
rect 10551 8588 10968 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 12986 8576 12992 8628
rect 13044 8616 13050 8628
rect 18506 8616 18512 8628
rect 13044 8588 18512 8616
rect 13044 8576 13050 8588
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 18877 8619 18935 8625
rect 18877 8585 18889 8619
rect 18923 8585 18935 8619
rect 18877 8579 18935 8585
rect 11422 8548 11428 8560
rect 8220 8520 11428 8548
rect 6822 8480 6828 8492
rect 6783 8452 6828 8480
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 4356 8384 6684 8412
rect 6932 8384 7236 8412
rect 4356 8356 4384 8384
rect 2777 8347 2835 8353
rect 2777 8313 2789 8347
rect 2823 8344 2835 8347
rect 3510 8344 3516 8356
rect 2823 8316 3516 8344
rect 2823 8313 2835 8316
rect 2777 8307 2835 8313
rect 3510 8304 3516 8316
rect 3568 8304 3574 8356
rect 4154 8304 4160 8356
rect 4212 8353 4218 8356
rect 4212 8347 4276 8353
rect 4212 8313 4230 8347
rect 4264 8313 4276 8347
rect 4212 8307 4276 8313
rect 4212 8304 4218 8307
rect 4338 8304 4344 8356
rect 4396 8304 4402 8356
rect 4706 8304 4712 8356
rect 4764 8344 4770 8356
rect 6932 8344 6960 8384
rect 7098 8353 7104 8356
rect 7092 8344 7104 8353
rect 4764 8316 6960 8344
rect 7059 8316 7104 8344
rect 4764 8304 4770 8316
rect 7092 8307 7104 8316
rect 7098 8304 7104 8307
rect 7156 8304 7162 8356
rect 7208 8344 7236 8384
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 8018 8412 8024 8424
rect 7432 8384 8024 8412
rect 7432 8372 7438 8384
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8220 8344 8248 8520
rect 11422 8508 11428 8520
rect 11480 8508 11486 8560
rect 12802 8508 12808 8560
rect 12860 8548 12866 8560
rect 13078 8548 13084 8560
rect 12860 8520 13084 8548
rect 12860 8508 12866 8520
rect 13078 8508 13084 8520
rect 13136 8508 13142 8560
rect 13906 8508 13912 8560
rect 13964 8548 13970 8560
rect 14734 8548 14740 8560
rect 13964 8520 14740 8548
rect 13964 8508 13970 8520
rect 14734 8508 14740 8520
rect 14792 8548 14798 8560
rect 15749 8551 15807 8557
rect 14792 8520 15148 8548
rect 14792 8508 14798 8520
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8480 9183 8483
rect 9306 8480 9312 8492
rect 9171 8452 9312 8480
rect 9171 8449 9183 8452
rect 9125 8443 9183 8449
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8480 10195 8483
rect 10226 8480 10232 8492
rect 10183 8452 10232 8480
rect 10183 8449 10195 8452
rect 10137 8443 10195 8449
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 10410 8440 10416 8492
rect 10468 8480 10474 8492
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10468 8452 11069 8480
rect 10468 8440 10474 8452
rect 11057 8449 11069 8452
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 11330 8440 11336 8492
rect 11388 8480 11394 8492
rect 12342 8480 12348 8492
rect 11388 8452 12348 8480
rect 11388 8440 11394 8452
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 12986 8480 12992 8492
rect 12947 8452 12992 8480
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 13998 8440 14004 8492
rect 14056 8480 14062 8492
rect 14056 8452 14101 8480
rect 14056 8440 14062 8452
rect 14366 8440 14372 8492
rect 14424 8480 14430 8492
rect 15120 8489 15148 8520
rect 15749 8517 15761 8551
rect 15795 8548 15807 8551
rect 15930 8548 15936 8560
rect 15795 8520 15936 8548
rect 15795 8517 15807 8520
rect 15749 8511 15807 8517
rect 15930 8508 15936 8520
rect 15988 8508 15994 8560
rect 17218 8508 17224 8560
rect 17276 8548 17282 8560
rect 18049 8551 18107 8557
rect 18049 8548 18061 8551
rect 17276 8520 18061 8548
rect 17276 8508 17282 8520
rect 18049 8517 18061 8520
rect 18095 8517 18107 8551
rect 18049 8511 18107 8517
rect 18322 8508 18328 8560
rect 18380 8548 18386 8560
rect 18892 8548 18920 8579
rect 18966 8576 18972 8628
rect 19024 8616 19030 8628
rect 19061 8619 19119 8625
rect 19061 8616 19073 8619
rect 19024 8588 19073 8616
rect 19024 8576 19030 8588
rect 19061 8585 19073 8588
rect 19107 8585 19119 8619
rect 19061 8579 19119 8585
rect 19242 8576 19248 8628
rect 19300 8616 19306 8628
rect 19978 8616 19984 8628
rect 19300 8588 19984 8616
rect 19300 8576 19306 8588
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 20073 8619 20131 8625
rect 20073 8585 20085 8619
rect 20119 8616 20131 8619
rect 20530 8616 20536 8628
rect 20119 8588 20536 8616
rect 20119 8585 20131 8588
rect 20073 8579 20131 8585
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 20162 8548 20168 8560
rect 18380 8520 18920 8548
rect 19444 8520 20168 8548
rect 18380 8508 18386 8520
rect 14921 8483 14979 8489
rect 14921 8480 14933 8483
rect 14424 8452 14933 8480
rect 14424 8440 14430 8452
rect 14921 8449 14933 8452
rect 14967 8449 14979 8483
rect 14921 8443 14979 8449
rect 15105 8483 15163 8489
rect 15105 8449 15117 8483
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 18601 8483 18659 8489
rect 18601 8480 18613 8483
rect 17920 8452 18613 8480
rect 17920 8440 17926 8452
rect 18601 8449 18613 8452
rect 18647 8449 18659 8483
rect 18601 8443 18659 8449
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8480 18935 8483
rect 19334 8480 19340 8492
rect 18923 8452 19340 8480
rect 18923 8449 18935 8452
rect 18877 8443 18935 8449
rect 19334 8440 19340 8452
rect 19392 8440 19398 8492
rect 8294 8372 8300 8424
rect 8352 8412 8358 8424
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 8352 8384 11805 8412
rect 8352 8372 8358 8384
rect 11793 8381 11805 8384
rect 11839 8412 11851 8415
rect 12434 8412 12440 8424
rect 11839 8384 12440 8412
rect 11839 8381 11851 8384
rect 11793 8375 11851 8381
rect 12434 8372 12440 8384
rect 12492 8372 12498 8424
rect 12802 8372 12808 8424
rect 12860 8412 12866 8424
rect 13630 8412 13636 8424
rect 12860 8384 13636 8412
rect 12860 8372 12866 8384
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 13814 8412 13820 8424
rect 13775 8384 13820 8412
rect 13814 8372 13820 8384
rect 13872 8372 13878 8424
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 14608 8384 14964 8412
rect 14608 8372 14614 8384
rect 7208 8316 8248 8344
rect 8389 8347 8447 8353
rect 8389 8313 8401 8347
rect 8435 8344 8447 8347
rect 8662 8344 8668 8356
rect 8435 8316 8668 8344
rect 8435 8313 8447 8316
rect 8389 8307 8447 8313
rect 8662 8304 8668 8316
rect 8720 8304 8726 8356
rect 8849 8347 8907 8353
rect 8849 8313 8861 8347
rect 8895 8344 8907 8347
rect 9309 8347 9367 8353
rect 9309 8344 9321 8347
rect 8895 8316 9321 8344
rect 8895 8313 8907 8316
rect 8849 8307 8907 8313
rect 9309 8313 9321 8316
rect 9355 8313 9367 8347
rect 9309 8307 9367 8313
rect 9861 8347 9919 8353
rect 9861 8313 9873 8347
rect 9907 8344 9919 8347
rect 10042 8344 10048 8356
rect 9907 8316 10048 8344
rect 9907 8313 9919 8316
rect 9861 8307 9919 8313
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 10226 8304 10232 8356
rect 10284 8304 10290 8356
rect 10410 8304 10416 8356
rect 10468 8344 10474 8356
rect 10965 8347 11023 8353
rect 10965 8344 10977 8347
rect 10468 8316 10977 8344
rect 10468 8304 10474 8316
rect 10965 8313 10977 8316
rect 11011 8313 11023 8347
rect 10965 8307 11023 8313
rect 12526 8304 12532 8356
rect 12584 8344 12590 8356
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 12584 8316 12909 8344
rect 12584 8304 12590 8316
rect 12897 8313 12909 8316
rect 12943 8313 12955 8347
rect 12897 8307 12955 8313
rect 13078 8304 13084 8356
rect 13136 8344 13142 8356
rect 14829 8347 14887 8353
rect 14829 8344 14841 8347
rect 13136 8316 14841 8344
rect 13136 8304 13142 8316
rect 14829 8313 14841 8316
rect 14875 8313 14887 8347
rect 14936 8344 14964 8384
rect 15010 8372 15016 8424
rect 15068 8412 15074 8424
rect 15565 8415 15623 8421
rect 15565 8412 15577 8415
rect 15068 8384 15577 8412
rect 15068 8372 15074 8384
rect 15565 8381 15577 8384
rect 15611 8381 15623 8415
rect 15565 8375 15623 8381
rect 15746 8372 15752 8424
rect 15804 8412 15810 8424
rect 15930 8412 15936 8424
rect 15804 8384 15936 8412
rect 15804 8372 15810 8384
rect 15930 8372 15936 8384
rect 15988 8412 15994 8424
rect 16117 8415 16175 8421
rect 16117 8412 16129 8415
rect 15988 8384 16129 8412
rect 15988 8372 15994 8384
rect 16117 8381 16129 8384
rect 16163 8381 16175 8415
rect 16117 8375 16175 8381
rect 16384 8415 16442 8421
rect 16384 8381 16396 8415
rect 16430 8412 16442 8415
rect 17126 8412 17132 8424
rect 16430 8384 17132 8412
rect 16430 8381 16442 8384
rect 16384 8375 16442 8381
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 18509 8415 18567 8421
rect 18509 8381 18521 8415
rect 18555 8412 18567 8415
rect 18966 8412 18972 8424
rect 18555 8384 18972 8412
rect 18555 8381 18567 8384
rect 18509 8375 18567 8381
rect 18966 8372 18972 8384
rect 19024 8412 19030 8424
rect 19444 8412 19472 8520
rect 20162 8508 20168 8520
rect 20220 8508 20226 8560
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 19024 8384 19472 8412
rect 19024 8372 19030 8384
rect 16298 8344 16304 8356
rect 14936 8316 16304 8344
rect 14829 8307 14887 8313
rect 16298 8304 16304 8316
rect 16356 8304 16362 8356
rect 17034 8304 17040 8356
rect 17092 8344 17098 8356
rect 18417 8347 18475 8353
rect 17092 8316 17540 8344
rect 17092 8304 17098 8316
rect 5166 8276 5172 8288
rect 2700 8248 5172 8276
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 6089 8279 6147 8285
rect 6089 8245 6101 8279
rect 6135 8276 6147 8279
rect 7374 8276 7380 8288
rect 6135 8248 7380 8276
rect 6135 8245 6147 8248
rect 6089 8239 6147 8245
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 7558 8236 7564 8288
rect 7616 8276 7622 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 7616 8248 8217 8276
rect 7616 8236 7622 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 8478 8276 8484 8288
rect 8439 8248 8484 8276
rect 8205 8239 8263 8245
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 8941 8279 8999 8285
rect 8941 8245 8953 8279
rect 8987 8276 8999 8279
rect 9493 8279 9551 8285
rect 9493 8276 9505 8279
rect 8987 8248 9505 8276
rect 8987 8245 8999 8248
rect 8941 8239 8999 8245
rect 9493 8245 9505 8248
rect 9539 8245 9551 8279
rect 9493 8239 9551 8245
rect 9953 8279 10011 8285
rect 9953 8245 9965 8279
rect 9999 8276 10011 8279
rect 10244 8276 10272 8304
rect 9999 8248 10272 8276
rect 9999 8245 10011 8248
rect 9953 8239 10011 8245
rect 10594 8236 10600 8288
rect 10652 8276 10658 8288
rect 10873 8279 10931 8285
rect 10873 8276 10885 8279
rect 10652 8248 10885 8276
rect 10652 8236 10658 8248
rect 10873 8245 10885 8248
rect 10919 8245 10931 8279
rect 10873 8239 10931 8245
rect 11977 8279 12035 8285
rect 11977 8245 11989 8279
rect 12023 8276 12035 8279
rect 12158 8276 12164 8288
rect 12023 8248 12164 8276
rect 12023 8245 12035 8248
rect 11977 8239 12035 8245
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 12805 8279 12863 8285
rect 12492 8248 12537 8276
rect 12492 8236 12498 8248
rect 12805 8245 12817 8279
rect 12851 8276 12863 8279
rect 13262 8276 13268 8288
rect 12851 8248 13268 8276
rect 12851 8245 12863 8248
rect 12805 8239 12863 8245
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 13446 8276 13452 8288
rect 13407 8248 13452 8276
rect 13446 8236 13452 8248
rect 13504 8236 13510 8288
rect 17512 8285 17540 8316
rect 18417 8313 18429 8347
rect 18463 8344 18475 8347
rect 18877 8347 18935 8353
rect 18877 8344 18889 8347
rect 18463 8316 18889 8344
rect 18463 8313 18475 8316
rect 18417 8307 18475 8313
rect 18877 8313 18889 8316
rect 18923 8313 18935 8347
rect 19521 8347 19579 8353
rect 19521 8344 19533 8347
rect 18877 8307 18935 8313
rect 18984 8316 19533 8344
rect 18984 8285 19012 8316
rect 19521 8313 19533 8316
rect 19567 8313 19579 8347
rect 19628 8344 19656 8443
rect 19978 8440 19984 8492
rect 20036 8480 20042 8492
rect 20622 8480 20628 8492
rect 20036 8452 20628 8480
rect 20036 8440 20042 8452
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 20438 8372 20444 8424
rect 20496 8412 20502 8424
rect 20533 8415 20591 8421
rect 20533 8412 20545 8415
rect 20496 8384 20545 8412
rect 20496 8372 20502 8384
rect 20533 8381 20545 8384
rect 20579 8381 20591 8415
rect 20533 8375 20591 8381
rect 19794 8344 19800 8356
rect 19628 8316 19800 8344
rect 19521 8307 19579 8313
rect 19794 8304 19800 8316
rect 19852 8304 19858 8356
rect 13909 8279 13967 8285
rect 13909 8245 13921 8279
rect 13955 8276 13967 8279
rect 14461 8279 14519 8285
rect 14461 8276 14473 8279
rect 13955 8248 14473 8276
rect 13955 8245 13967 8248
rect 13909 8239 13967 8245
rect 14461 8245 14473 8248
rect 14507 8245 14519 8279
rect 14461 8239 14519 8245
rect 17497 8279 17555 8285
rect 17497 8245 17509 8279
rect 17543 8245 17555 8279
rect 17497 8239 17555 8245
rect 18969 8279 19027 8285
rect 18969 8245 18981 8279
rect 19015 8245 19027 8279
rect 19426 8276 19432 8288
rect 19387 8248 19432 8276
rect 18969 8239 19027 8245
rect 19426 8236 19432 8248
rect 19484 8236 19490 8288
rect 19610 8236 19616 8288
rect 19668 8276 19674 8288
rect 20441 8279 20499 8285
rect 20441 8276 20453 8279
rect 19668 8248 20453 8276
rect 19668 8236 19674 8248
rect 20441 8245 20453 8248
rect 20487 8245 20499 8279
rect 20441 8239 20499 8245
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 3418 8072 3424 8084
rect 2179 8044 3424 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 4065 8075 4123 8081
rect 4065 8041 4077 8075
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 4571 8044 5089 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 5077 8041 5089 8044
rect 5123 8041 5135 8075
rect 5077 8035 5135 8041
rect 5537 8075 5595 8081
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 6546 8072 6552 8084
rect 5583 8044 6552 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 4080 8004 4108 8035
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 6917 8075 6975 8081
rect 6917 8041 6929 8075
rect 6963 8041 6975 8075
rect 6917 8035 6975 8041
rect 7377 8075 7435 8081
rect 7377 8041 7389 8075
rect 7423 8072 7435 8075
rect 12434 8072 12440 8084
rect 7423 8044 12440 8072
rect 7423 8041 7435 8044
rect 7377 8035 7435 8041
rect 1596 7976 4108 8004
rect 6932 8004 6960 8035
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 14921 8075 14979 8081
rect 14921 8072 14933 8075
rect 14424 8044 14933 8072
rect 14424 8032 14430 8044
rect 14921 8041 14933 8044
rect 14967 8072 14979 8075
rect 15010 8072 15016 8084
rect 14967 8044 15016 8072
rect 14967 8041 14979 8044
rect 14921 8035 14979 8041
rect 15010 8032 15016 8044
rect 15068 8032 15074 8084
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 15289 8075 15347 8081
rect 15289 8072 15301 8075
rect 15252 8044 15301 8072
rect 15252 8032 15258 8044
rect 15289 8041 15301 8044
rect 15335 8041 15347 8075
rect 17862 8072 17868 8084
rect 15289 8035 15347 8041
rect 17144 8044 17868 8072
rect 10226 8004 10232 8016
rect 6932 7976 10232 8004
rect 1596 7945 1624 7976
rect 10226 7964 10232 7976
rect 10284 7964 10290 8016
rect 10864 8007 10922 8013
rect 10864 7973 10876 8007
rect 10910 8004 10922 8007
rect 11054 8004 11060 8016
rect 10910 7976 11060 8004
rect 10910 7973 10922 7976
rect 10864 7967 10922 7973
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 11422 7964 11428 8016
rect 11480 8004 11486 8016
rect 12250 8004 12256 8016
rect 11480 7976 12256 8004
rect 11480 7964 11486 7976
rect 12250 7964 12256 7976
rect 12308 8004 12314 8016
rect 12621 8007 12679 8013
rect 12621 8004 12633 8007
rect 12308 7976 12633 8004
rect 12308 7964 12314 7976
rect 12621 7973 12633 7976
rect 12667 7973 12679 8007
rect 12621 7967 12679 7973
rect 12713 8007 12771 8013
rect 12713 7973 12725 8007
rect 12759 8004 12771 8007
rect 13354 8004 13360 8016
rect 12759 7976 13360 8004
rect 12759 7973 12771 7976
rect 12713 7967 12771 7973
rect 13354 7964 13360 7976
rect 13412 7964 13418 8016
rect 14090 8004 14096 8016
rect 13464 7976 14096 8004
rect 2590 7945 2596 7948
rect 1581 7939 1639 7945
rect 1581 7905 1593 7939
rect 1627 7905 1639 7939
rect 1581 7899 1639 7905
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7936 1915 7939
rect 2133 7939 2191 7945
rect 2133 7936 2145 7939
rect 1903 7908 2145 7936
rect 1903 7905 1915 7908
rect 1857 7899 1915 7905
rect 2133 7905 2145 7908
rect 2179 7905 2191 7939
rect 2133 7899 2191 7905
rect 2584 7899 2596 7945
rect 2648 7936 2654 7948
rect 2648 7908 2684 7936
rect 2590 7896 2596 7899
rect 2648 7896 2654 7908
rect 2958 7896 2964 7948
rect 3016 7936 3022 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 3016 7908 4445 7936
rect 3016 7896 3022 7908
rect 4433 7905 4445 7908
rect 4479 7905 4491 7939
rect 5442 7936 5448 7948
rect 5403 7908 5448 7936
rect 4433 7899 4491 7905
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 6270 7936 6276 7948
rect 6231 7908 6276 7936
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6365 7939 6423 7945
rect 6365 7905 6377 7939
rect 6411 7905 6423 7939
rect 6365 7899 6423 7905
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7936 7343 7939
rect 7929 7939 7987 7945
rect 7331 7908 7880 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 1854 7692 1860 7744
rect 1912 7732 1918 7744
rect 2332 7732 2360 7831
rect 3697 7803 3755 7809
rect 3697 7769 3709 7803
rect 3743 7800 3755 7803
rect 4154 7800 4160 7812
rect 3743 7772 4160 7800
rect 3743 7769 3755 7772
rect 3697 7763 3755 7769
rect 4154 7760 4160 7772
rect 4212 7800 4218 7812
rect 4632 7800 4660 7831
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 5629 7871 5687 7877
rect 5629 7868 5641 7871
rect 4764 7840 5641 7868
rect 4764 7828 4770 7840
rect 5629 7837 5641 7840
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 6380 7868 6408 7899
rect 5960 7840 6408 7868
rect 7561 7871 7619 7877
rect 5960 7828 5966 7840
rect 7561 7837 7573 7871
rect 7607 7868 7619 7871
rect 7650 7868 7656 7880
rect 7607 7840 7656 7868
rect 7607 7837 7619 7840
rect 7561 7831 7619 7837
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 4212 7772 4660 7800
rect 4212 7760 4218 7772
rect 5534 7760 5540 7812
rect 5592 7800 5598 7812
rect 6089 7803 6147 7809
rect 6089 7800 6101 7803
rect 5592 7772 6101 7800
rect 5592 7760 5598 7772
rect 6089 7769 6101 7772
rect 6135 7769 6147 7803
rect 6089 7763 6147 7769
rect 6380 7772 7696 7800
rect 3970 7732 3976 7744
rect 1912 7704 3976 7732
rect 1912 7692 1918 7704
rect 3970 7692 3976 7704
rect 4028 7692 4034 7744
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 6380 7732 6408 7772
rect 7668 7744 7696 7772
rect 6546 7732 6552 7744
rect 4120 7704 6408 7732
rect 6507 7704 6552 7732
rect 4120 7692 4126 7704
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 7650 7692 7656 7744
rect 7708 7692 7714 7744
rect 7852 7732 7880 7908
rect 7929 7905 7941 7939
rect 7975 7936 7987 7939
rect 8018 7936 8024 7948
rect 7975 7908 8024 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 8018 7896 8024 7908
rect 8076 7896 8082 7948
rect 8202 7945 8208 7948
rect 8196 7936 8208 7945
rect 8163 7908 8208 7936
rect 8196 7899 8208 7908
rect 8202 7896 8208 7899
rect 8260 7896 8266 7948
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 9953 7939 10011 7945
rect 9953 7936 9965 7939
rect 9180 7908 9965 7936
rect 9180 7896 9186 7908
rect 9953 7905 9965 7908
rect 9999 7905 10011 7939
rect 9953 7899 10011 7905
rect 10597 7939 10655 7945
rect 10597 7905 10609 7939
rect 10643 7936 10655 7939
rect 10686 7936 10692 7948
rect 10643 7908 10692 7936
rect 10643 7905 10655 7908
rect 10597 7899 10655 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 13464 7945 13492 7976
rect 14090 7964 14096 7976
rect 14148 8004 14154 8016
rect 14148 7976 16528 8004
rect 14148 7964 14154 7976
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7905 13507 7939
rect 13630 7936 13636 7948
rect 13449 7899 13507 7905
rect 13556 7908 13636 7936
rect 9214 7828 9220 7880
rect 9272 7868 9278 7880
rect 10410 7868 10416 7880
rect 9272 7840 10416 7868
rect 9272 7828 9278 7840
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7868 12955 7871
rect 12986 7868 12992 7880
rect 12943 7840 12992 7868
rect 12943 7837 12955 7840
rect 12897 7831 12955 7837
rect 8938 7760 8944 7812
rect 8996 7800 9002 7812
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 8996 7772 9321 7800
rect 8996 7760 9002 7772
rect 9309 7769 9321 7772
rect 9355 7800 9367 7803
rect 9398 7800 9404 7812
rect 9355 7772 9404 7800
rect 9355 7769 9367 7772
rect 9309 7763 9367 7769
rect 9398 7760 9404 7772
rect 9456 7760 9462 7812
rect 10042 7760 10048 7812
rect 10100 7800 10106 7812
rect 10226 7800 10232 7812
rect 10100 7772 10232 7800
rect 10100 7760 10106 7772
rect 10226 7760 10232 7772
rect 10284 7760 10290 7812
rect 12912 7800 12940 7831
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 13556 7877 13584 7908
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 13808 7939 13866 7945
rect 13808 7905 13820 7939
rect 13854 7936 13866 7939
rect 14642 7936 14648 7948
rect 13854 7908 14648 7936
rect 13854 7905 13866 7908
rect 13808 7899 13866 7905
rect 14642 7896 14648 7908
rect 14700 7896 14706 7948
rect 15010 7896 15016 7948
rect 15068 7936 15074 7948
rect 16500 7945 16528 7976
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 15068 7908 15669 7936
rect 15068 7896 15074 7908
rect 15657 7905 15669 7908
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 16485 7939 16543 7945
rect 16485 7905 16497 7939
rect 16531 7905 16543 7939
rect 16485 7899 16543 7905
rect 16577 7939 16635 7945
rect 16577 7905 16589 7939
rect 16623 7936 16635 7939
rect 17034 7936 17040 7948
rect 16623 7908 17040 7936
rect 16623 7905 16635 7908
rect 16577 7899 16635 7905
rect 17034 7896 17040 7908
rect 17092 7896 17098 7948
rect 17144 7945 17172 8044
rect 17862 8032 17868 8044
rect 17920 8072 17926 8084
rect 18046 8072 18052 8084
rect 17920 8044 18052 8072
rect 17920 8032 17926 8044
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 18322 8032 18328 8084
rect 18380 8072 18386 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 18380 8044 18613 8072
rect 18380 8032 18386 8044
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 19797 8075 19855 8081
rect 18601 8035 18659 8041
rect 19067 8044 19564 8072
rect 17954 7964 17960 8016
rect 18012 8004 18018 8016
rect 19067 8004 19095 8044
rect 19334 8004 19340 8016
rect 18012 7976 19095 8004
rect 19168 7976 19340 8004
rect 18012 7964 18018 7976
rect 17129 7939 17187 7945
rect 17129 7905 17141 7939
rect 17175 7905 17187 7939
rect 17129 7899 17187 7905
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7868 13231 7871
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13219 7840 13553 7868
rect 13219 7837 13231 7840
rect 13173 7831 13231 7837
rect 13541 7837 13553 7840
rect 13587 7837 13599 7871
rect 15746 7868 15752 7880
rect 15707 7840 15752 7868
rect 13541 7831 13599 7837
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7837 15899 7871
rect 17144 7868 17172 7899
rect 17218 7896 17224 7948
rect 17276 7936 17282 7948
rect 17385 7939 17443 7945
rect 17385 7936 17397 7939
rect 17276 7908 17397 7936
rect 17276 7896 17282 7908
rect 17385 7905 17397 7908
rect 17431 7905 17443 7939
rect 17385 7899 17443 7905
rect 17678 7896 17684 7948
rect 17736 7936 17742 7948
rect 18969 7939 19027 7945
rect 18969 7936 18981 7939
rect 17736 7908 18981 7936
rect 17736 7896 17742 7908
rect 18969 7905 18981 7908
rect 19015 7905 19027 7939
rect 18969 7899 19027 7905
rect 19061 7939 19119 7945
rect 19061 7905 19073 7939
rect 19107 7936 19119 7939
rect 19168 7936 19196 7976
rect 19334 7964 19340 7976
rect 19392 7964 19398 8016
rect 19536 8004 19564 8044
rect 19797 8041 19809 8075
rect 19843 8072 19855 8075
rect 19886 8072 19892 8084
rect 19843 8044 19892 8072
rect 19843 8041 19855 8044
rect 19797 8035 19855 8041
rect 19886 8032 19892 8044
rect 19944 8032 19950 8084
rect 20162 8032 20168 8084
rect 20220 8072 20226 8084
rect 21821 8075 21879 8081
rect 21821 8072 21833 8075
rect 20220 8044 21833 8072
rect 20220 8032 20226 8044
rect 21821 8041 21833 8044
rect 21867 8041 21879 8075
rect 21821 8035 21879 8041
rect 19536 7976 20208 8004
rect 19978 7936 19984 7948
rect 19107 7908 19196 7936
rect 19536 7908 19984 7936
rect 19107 7905 19119 7908
rect 19061 7899 19119 7905
rect 15841 7831 15899 7837
rect 16316 7840 17172 7868
rect 19245 7871 19303 7877
rect 11808 7772 12940 7800
rect 8846 7732 8852 7744
rect 7852 7704 8852 7732
rect 8846 7692 8852 7704
rect 8904 7692 8910 7744
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 9674 7732 9680 7744
rect 9272 7704 9680 7732
rect 9272 7692 9278 7704
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 10137 7735 10195 7741
rect 10137 7701 10149 7735
rect 10183 7732 10195 7735
rect 10594 7732 10600 7744
rect 10183 7704 10600 7732
rect 10183 7701 10195 7704
rect 10137 7695 10195 7701
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 10870 7692 10876 7744
rect 10928 7732 10934 7744
rect 11808 7732 11836 7772
rect 13078 7760 13084 7812
rect 13136 7800 13142 7812
rect 15013 7803 15071 7809
rect 13136 7772 13400 7800
rect 13136 7760 13142 7772
rect 11974 7732 11980 7744
rect 10928 7704 11836 7732
rect 11935 7704 11980 7732
rect 10928 7692 10934 7704
rect 11974 7692 11980 7704
rect 12032 7692 12038 7744
rect 12250 7732 12256 7744
rect 12211 7704 12256 7732
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 12434 7692 12440 7744
rect 12492 7732 12498 7744
rect 12894 7732 12900 7744
rect 12492 7704 12900 7732
rect 12492 7692 12498 7704
rect 12894 7692 12900 7704
rect 12952 7732 12958 7744
rect 13173 7735 13231 7741
rect 13173 7732 13185 7735
rect 12952 7704 13185 7732
rect 12952 7692 12958 7704
rect 13173 7701 13185 7704
rect 13219 7732 13231 7735
rect 13265 7735 13323 7741
rect 13265 7732 13277 7735
rect 13219 7704 13277 7732
rect 13219 7701 13231 7704
rect 13173 7695 13231 7701
rect 13265 7701 13277 7704
rect 13311 7701 13323 7735
rect 13372 7732 13400 7772
rect 15013 7769 15025 7803
rect 15059 7800 15071 7803
rect 15856 7800 15884 7831
rect 16206 7800 16212 7812
rect 15059 7772 16212 7800
rect 15059 7769 15071 7772
rect 15013 7763 15071 7769
rect 16206 7760 16212 7772
rect 16264 7760 16270 7812
rect 14734 7732 14740 7744
rect 13372 7704 14740 7732
rect 13265 7695 13323 7701
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 15930 7692 15936 7744
rect 15988 7732 15994 7744
rect 16316 7741 16344 7840
rect 19245 7837 19257 7871
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 18690 7800 18696 7812
rect 18432 7772 18696 7800
rect 16301 7735 16359 7741
rect 16301 7732 16313 7735
rect 15988 7704 16313 7732
rect 15988 7692 15994 7704
rect 16301 7701 16313 7704
rect 16347 7701 16359 7735
rect 16301 7695 16359 7701
rect 16761 7735 16819 7741
rect 16761 7701 16773 7735
rect 16807 7732 16819 7735
rect 18432 7732 18460 7772
rect 18690 7760 18696 7772
rect 18748 7760 18754 7812
rect 19260 7800 19288 7831
rect 19536 7800 19564 7908
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 20180 7945 20208 7976
rect 20346 7964 20352 8016
rect 20404 8004 20410 8016
rect 21082 8004 21088 8016
rect 20404 7976 21088 8004
rect 20404 7964 20410 7976
rect 21082 7964 21088 7976
rect 21140 7964 21146 8016
rect 20165 7939 20223 7945
rect 20165 7905 20177 7939
rect 20211 7936 20223 7939
rect 20530 7936 20536 7948
rect 20211 7908 20536 7936
rect 20211 7905 20223 7908
rect 20165 7899 20223 7905
rect 20530 7896 20536 7908
rect 20588 7896 20594 7948
rect 20257 7871 20315 7877
rect 20257 7868 20269 7871
rect 19720 7840 20269 7868
rect 19720 7809 19748 7840
rect 20257 7837 20269 7840
rect 20303 7837 20315 7871
rect 20257 7831 20315 7837
rect 19260 7772 19564 7800
rect 19705 7803 19763 7809
rect 19705 7769 19717 7803
rect 19751 7769 19763 7803
rect 20272 7800 20300 7831
rect 20346 7828 20352 7880
rect 20404 7868 20410 7880
rect 20404 7840 20449 7868
rect 20404 7828 20410 7840
rect 20714 7800 20720 7812
rect 20272 7772 20720 7800
rect 19705 7763 19763 7769
rect 20714 7760 20720 7772
rect 20772 7760 20778 7812
rect 16807 7704 18460 7732
rect 18509 7735 18567 7741
rect 16807 7701 16819 7704
rect 16761 7695 16819 7701
rect 18509 7701 18521 7735
rect 18555 7732 18567 7735
rect 18598 7732 18604 7744
rect 18555 7704 18604 7732
rect 18555 7701 18567 7704
rect 18509 7695 18567 7701
rect 18598 7692 18604 7704
rect 18656 7692 18662 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 2740 7500 3157 7528
rect 2740 7488 2746 7500
rect 3145 7497 3157 7500
rect 3191 7528 3203 7531
rect 4706 7528 4712 7540
rect 3191 7500 4712 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 5166 7528 5172 7540
rect 5127 7500 5172 7528
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 5442 7528 5448 7540
rect 5403 7500 5448 7528
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 6270 7488 6276 7540
rect 6328 7528 6334 7540
rect 8570 7528 8576 7540
rect 6328 7500 8576 7528
rect 6328 7488 6334 7500
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 8849 7531 8907 7537
rect 8849 7497 8861 7531
rect 8895 7528 8907 7531
rect 8895 7500 9352 7528
rect 8895 7497 8907 7500
rect 8849 7491 8907 7497
rect 6638 7420 6644 7472
rect 6696 7460 6702 7472
rect 7098 7460 7104 7472
rect 6696 7432 7104 7460
rect 6696 7420 6702 7432
rect 7098 7420 7104 7432
rect 7156 7420 7162 7472
rect 8202 7420 8208 7472
rect 8260 7460 8266 7472
rect 8481 7463 8539 7469
rect 8481 7460 8493 7463
rect 8260 7432 8493 7460
rect 8260 7420 8266 7432
rect 8481 7429 8493 7432
rect 8527 7460 8539 7463
rect 9214 7460 9220 7472
rect 8527 7432 9220 7460
rect 8527 7429 8539 7432
rect 8481 7423 8539 7429
rect 9214 7420 9220 7432
rect 9272 7420 9278 7472
rect 9324 7460 9352 7500
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 16390 7528 16396 7540
rect 9640 7500 14504 7528
rect 16351 7500 16396 7528
rect 9640 7488 9646 7500
rect 10226 7460 10232 7472
rect 9324 7432 10232 7460
rect 10226 7420 10232 7432
rect 10284 7420 10290 7472
rect 10962 7420 10968 7472
rect 11020 7460 11026 7472
rect 12250 7460 12256 7472
rect 11020 7432 12256 7460
rect 11020 7420 11026 7432
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 14093 7463 14151 7469
rect 14093 7429 14105 7463
rect 14139 7460 14151 7463
rect 14182 7460 14188 7472
rect 14139 7432 14188 7460
rect 14139 7429 14151 7432
rect 14093 7423 14151 7429
rect 14182 7420 14188 7432
rect 14240 7420 14246 7472
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 5224 7364 6009 7392
rect 5224 7352 5230 7364
rect 5997 7361 6009 7364
rect 6043 7392 6055 7395
rect 6914 7392 6920 7404
rect 6043 7364 6920 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 9398 7392 9404 7404
rect 9359 7364 9404 7392
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 10502 7392 10508 7404
rect 10463 7364 10508 7392
rect 10502 7352 10508 7364
rect 10560 7392 10566 7404
rect 11425 7395 11483 7401
rect 11425 7392 11437 7395
rect 10560 7364 11437 7392
rect 10560 7352 10566 7364
rect 11425 7361 11437 7364
rect 11471 7361 11483 7395
rect 11425 7355 11483 7361
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 14366 7392 14372 7404
rect 11664 7364 12572 7392
rect 11664 7352 11670 7364
rect 12544 7336 12572 7364
rect 13648 7364 14372 7392
rect 1765 7327 1823 7333
rect 1765 7293 1777 7327
rect 1811 7324 1823 7327
rect 1854 7324 1860 7336
rect 1811 7296 1860 7324
rect 1811 7293 1823 7296
rect 1765 7287 1823 7293
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 2038 7333 2044 7336
rect 2032 7287 2044 7333
rect 2096 7324 2102 7336
rect 3789 7327 3847 7333
rect 2096 7296 2132 7324
rect 2038 7284 2044 7287
rect 2096 7284 2102 7296
rect 3789 7293 3801 7327
rect 3835 7324 3847 7327
rect 3878 7324 3884 7336
rect 3835 7296 3884 7324
rect 3835 7293 3847 7296
rect 3789 7287 3847 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7324 5871 7327
rect 6086 7324 6092 7336
rect 5859 7296 6092 7324
rect 5859 7293 5871 7296
rect 5813 7287 5871 7293
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7324 7159 7327
rect 7926 7324 7932 7336
rect 7147 7296 7932 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7926 7284 7932 7296
rect 7984 7324 7990 7336
rect 8294 7324 8300 7336
rect 7984 7296 8300 7324
rect 7984 7284 7990 7296
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 9309 7327 9367 7333
rect 9309 7293 9321 7327
rect 9355 7324 9367 7327
rect 10962 7324 10968 7336
rect 9355 7296 10968 7324
rect 9355 7293 9367 7296
rect 9309 7287 9367 7293
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11514 7324 11520 7336
rect 11072 7296 11520 7324
rect 3326 7216 3332 7268
rect 3384 7256 3390 7268
rect 4034 7259 4092 7265
rect 4034 7256 4046 7259
rect 3384 7228 4046 7256
rect 3384 7216 3390 7228
rect 3804 7200 3832 7228
rect 4034 7225 4046 7228
rect 4080 7225 4092 7259
rect 4034 7219 4092 7225
rect 4706 7216 4712 7268
rect 4764 7256 4770 7268
rect 4890 7256 4896 7268
rect 4764 7228 4896 7256
rect 4764 7216 4770 7228
rect 4890 7216 4896 7228
rect 4948 7216 4954 7268
rect 7368 7259 7426 7265
rect 7368 7225 7380 7259
rect 7414 7256 7426 7259
rect 8202 7256 8208 7268
rect 7414 7228 8208 7256
rect 7414 7225 7426 7228
rect 7368 7219 7426 7225
rect 8202 7216 8208 7228
rect 8260 7216 8266 7268
rect 8938 7216 8944 7268
rect 8996 7256 9002 7268
rect 9490 7256 9496 7268
rect 8996 7228 9496 7256
rect 8996 7216 9002 7228
rect 9490 7216 9496 7228
rect 9548 7216 9554 7268
rect 9674 7216 9680 7268
rect 9732 7256 9738 7268
rect 10321 7259 10379 7265
rect 10321 7256 10333 7259
rect 9732 7228 10333 7256
rect 9732 7216 9738 7228
rect 10321 7225 10333 7228
rect 10367 7225 10379 7259
rect 10321 7219 10379 7225
rect 10410 7216 10416 7268
rect 10468 7256 10474 7268
rect 11072 7256 11100 7296
rect 11514 7284 11520 7296
rect 11572 7284 11578 7336
rect 12434 7324 12440 7336
rect 12395 7296 12440 7324
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 12526 7284 12532 7336
rect 12584 7284 12590 7336
rect 12704 7327 12762 7333
rect 12704 7293 12716 7327
rect 12750 7324 12762 7327
rect 13648 7324 13676 7364
rect 14366 7352 14372 7364
rect 14424 7352 14430 7404
rect 12750 7296 13676 7324
rect 12750 7293 12762 7296
rect 12704 7287 12762 7293
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 14476 7333 14504 7500
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 17589 7531 17647 7537
rect 17589 7497 17601 7531
rect 17635 7528 17647 7531
rect 17954 7528 17960 7540
rect 17635 7500 17960 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 18877 7531 18935 7537
rect 18877 7497 18889 7531
rect 18923 7528 18935 7531
rect 19150 7528 19156 7540
rect 18923 7500 19156 7528
rect 18923 7497 18935 7500
rect 18877 7491 18935 7497
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 19610 7488 19616 7540
rect 19668 7528 19674 7540
rect 20073 7531 20131 7537
rect 20073 7528 20085 7531
rect 19668 7500 20085 7528
rect 19668 7488 19674 7500
rect 20073 7497 20085 7500
rect 20119 7497 20131 7531
rect 20073 7491 20131 7497
rect 14734 7420 14740 7472
rect 14792 7460 14798 7472
rect 20346 7460 20352 7472
rect 14792 7432 20352 7460
rect 14792 7420 14798 7432
rect 14642 7392 14648 7404
rect 14603 7364 14648 7392
rect 14642 7352 14648 7364
rect 14700 7392 14706 7404
rect 15102 7392 15108 7404
rect 14700 7364 15108 7392
rect 14700 7352 14706 7364
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 15838 7392 15844 7404
rect 15799 7364 15844 7392
rect 15838 7352 15844 7364
rect 15896 7352 15902 7404
rect 16022 7392 16028 7404
rect 15983 7364 16028 7392
rect 16022 7352 16028 7364
rect 16080 7352 16086 7404
rect 16206 7352 16212 7404
rect 16264 7392 16270 7404
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 16264 7364 16957 7392
rect 16264 7352 16270 7364
rect 16945 7361 16957 7364
rect 16991 7361 17003 7395
rect 17678 7392 17684 7404
rect 16945 7355 17003 7361
rect 17328 7364 17684 7392
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 13780 7296 14013 7324
rect 13780 7284 13786 7296
rect 14001 7293 14013 7296
rect 14047 7293 14059 7327
rect 14001 7287 14059 7293
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7293 14519 7327
rect 17328 7324 17356 7364
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 17788 7364 18613 7392
rect 14461 7287 14519 7293
rect 14568 7296 17356 7324
rect 17405 7327 17463 7333
rect 10468 7228 11100 7256
rect 11241 7259 11299 7265
rect 10468 7216 10474 7228
rect 11241 7225 11253 7259
rect 11287 7256 11299 7259
rect 11606 7256 11612 7268
rect 11287 7228 11612 7256
rect 11287 7225 11299 7228
rect 11241 7219 11299 7225
rect 11606 7216 11612 7228
rect 11664 7216 11670 7268
rect 11885 7259 11943 7265
rect 11885 7225 11897 7259
rect 11931 7256 11943 7259
rect 13538 7256 13544 7268
rect 11931 7228 13544 7256
rect 11931 7225 11943 7228
rect 11885 7219 11943 7225
rect 13538 7216 13544 7228
rect 13596 7216 13602 7268
rect 14568 7265 14596 7296
rect 17405 7293 17417 7327
rect 17451 7293 17463 7327
rect 17405 7287 17463 7293
rect 14553 7259 14611 7265
rect 14553 7256 14565 7259
rect 13648 7228 14565 7256
rect 2038 7148 2044 7200
rect 2096 7188 2102 7200
rect 2406 7188 2412 7200
rect 2096 7160 2412 7188
rect 2096 7148 2102 7160
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 3786 7148 3792 7200
rect 3844 7148 3850 7200
rect 5905 7191 5963 7197
rect 5905 7157 5917 7191
rect 5951 7188 5963 7191
rect 7742 7188 7748 7200
rect 5951 7160 7748 7188
rect 5951 7157 5963 7160
rect 5905 7151 5963 7157
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 8846 7148 8852 7200
rect 8904 7188 8910 7200
rect 9217 7191 9275 7197
rect 9217 7188 9229 7191
rect 8904 7160 9229 7188
rect 8904 7148 8910 7160
rect 9217 7157 9229 7160
rect 9263 7188 9275 7191
rect 9582 7188 9588 7200
rect 9263 7160 9588 7188
rect 9263 7157 9275 7160
rect 9217 7151 9275 7157
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 9858 7188 9864 7200
rect 9819 7160 9864 7188
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 10226 7188 10232 7200
rect 10187 7160 10232 7188
rect 10226 7148 10232 7160
rect 10284 7148 10290 7200
rect 10870 7188 10876 7200
rect 10831 7160 10876 7188
rect 10870 7148 10876 7160
rect 10928 7148 10934 7200
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 11020 7160 11345 7188
rect 11020 7148 11026 7160
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 11333 7151 11391 7157
rect 11422 7148 11428 7200
rect 11480 7188 11486 7200
rect 13648 7188 13676 7228
rect 14553 7225 14565 7228
rect 14599 7225 14611 7259
rect 16853 7259 16911 7265
rect 16853 7256 16865 7259
rect 14553 7219 14611 7225
rect 15304 7228 16865 7256
rect 13814 7188 13820 7200
rect 11480 7160 13676 7188
rect 13775 7160 13820 7188
rect 11480 7148 11486 7160
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 14001 7191 14059 7197
rect 14001 7157 14013 7191
rect 14047 7188 14059 7191
rect 15304 7188 15332 7228
rect 16853 7225 16865 7228
rect 16899 7225 16911 7259
rect 17420 7256 17448 7287
rect 17494 7284 17500 7336
rect 17552 7324 17558 7336
rect 17788 7324 17816 7364
rect 18601 7361 18613 7364
rect 18647 7392 18659 7395
rect 19334 7392 19340 7404
rect 18647 7364 19340 7392
rect 18647 7361 18659 7364
rect 18601 7355 18659 7361
rect 19334 7352 19340 7364
rect 19392 7352 19398 7404
rect 19426 7352 19432 7404
rect 19484 7352 19490 7404
rect 19720 7401 19748 7432
rect 20346 7420 20352 7432
rect 20404 7420 20410 7472
rect 19705 7395 19763 7401
rect 19705 7361 19717 7395
rect 19751 7361 19763 7395
rect 19705 7355 19763 7361
rect 19794 7352 19800 7404
rect 19852 7392 19858 7404
rect 20625 7395 20683 7401
rect 20625 7392 20637 7395
rect 19852 7364 20637 7392
rect 19852 7352 19858 7364
rect 20625 7361 20637 7364
rect 20671 7361 20683 7395
rect 20625 7355 20683 7361
rect 17552 7296 17816 7324
rect 18417 7327 18475 7333
rect 17552 7284 17558 7296
rect 18417 7293 18429 7327
rect 18463 7324 18475 7327
rect 18506 7324 18512 7336
rect 18463 7296 18512 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 18506 7284 18512 7296
rect 18564 7284 18570 7336
rect 18969 7327 19027 7333
rect 18969 7293 18981 7327
rect 19015 7324 19027 7327
rect 19444 7324 19472 7352
rect 19015 7296 19472 7324
rect 19521 7327 19579 7333
rect 19015 7293 19027 7296
rect 18969 7287 19027 7293
rect 19521 7293 19533 7327
rect 19567 7324 19579 7327
rect 21082 7324 21088 7336
rect 19567 7296 21088 7324
rect 19567 7293 19579 7296
rect 19521 7287 19579 7293
rect 21082 7284 21088 7296
rect 21140 7284 21146 7336
rect 19794 7256 19800 7268
rect 17420 7228 19800 7256
rect 16853 7219 16911 7225
rect 19794 7216 19800 7228
rect 19852 7216 19858 7268
rect 14047 7160 15332 7188
rect 15381 7191 15439 7197
rect 14047 7157 14059 7160
rect 14001 7151 14059 7157
rect 15381 7157 15393 7191
rect 15427 7188 15439 7191
rect 15654 7188 15660 7200
rect 15427 7160 15660 7188
rect 15427 7157 15439 7160
rect 15381 7151 15439 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 15749 7191 15807 7197
rect 15749 7157 15761 7191
rect 15795 7188 15807 7191
rect 15930 7188 15936 7200
rect 15795 7160 15936 7188
rect 15795 7157 15807 7160
rect 15749 7151 15807 7157
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 16206 7148 16212 7200
rect 16264 7188 16270 7200
rect 16761 7191 16819 7197
rect 16761 7188 16773 7191
rect 16264 7160 16773 7188
rect 16264 7148 16270 7160
rect 16761 7157 16773 7160
rect 16807 7157 16819 7191
rect 18046 7188 18052 7200
rect 18007 7160 18052 7188
rect 16761 7151 16819 7157
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 18509 7191 18567 7197
rect 18509 7157 18521 7191
rect 18555 7188 18567 7191
rect 18877 7191 18935 7197
rect 18877 7188 18889 7191
rect 18555 7160 18889 7188
rect 18555 7157 18567 7160
rect 18509 7151 18567 7157
rect 18877 7157 18889 7160
rect 18923 7157 18935 7191
rect 18877 7151 18935 7157
rect 18969 7191 19027 7197
rect 18969 7157 18981 7191
rect 19015 7188 19027 7191
rect 19061 7191 19119 7197
rect 19061 7188 19073 7191
rect 19015 7160 19073 7188
rect 19015 7157 19027 7160
rect 18969 7151 19027 7157
rect 19061 7157 19073 7160
rect 19107 7157 19119 7191
rect 19061 7151 19119 7157
rect 19242 7148 19248 7200
rect 19300 7188 19306 7200
rect 19429 7191 19487 7197
rect 19429 7188 19441 7191
rect 19300 7160 19441 7188
rect 19300 7148 19306 7160
rect 19429 7157 19441 7160
rect 19475 7157 19487 7191
rect 19429 7151 19487 7157
rect 19610 7148 19616 7200
rect 19668 7188 19674 7200
rect 20441 7191 20499 7197
rect 20441 7188 20453 7191
rect 19668 7160 20453 7188
rect 19668 7148 19674 7160
rect 20441 7157 20453 7160
rect 20487 7157 20499 7191
rect 20441 7151 20499 7157
rect 20533 7191 20591 7197
rect 20533 7157 20545 7191
rect 20579 7188 20591 7191
rect 21634 7188 21640 7200
rect 20579 7160 21640 7188
rect 20579 7157 20591 7160
rect 20533 7151 20591 7157
rect 21634 7148 21640 7160
rect 21692 7148 21698 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 2501 6987 2559 6993
rect 2501 6984 2513 6987
rect 1452 6956 2513 6984
rect 1452 6944 1458 6956
rect 2501 6953 2513 6956
rect 2547 6953 2559 6987
rect 3602 6984 3608 6996
rect 3563 6956 3608 6984
rect 2501 6947 2559 6953
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 5810 6944 5816 6996
rect 5868 6984 5874 6996
rect 8941 6987 8999 6993
rect 5868 6956 8791 6984
rect 5868 6944 5874 6956
rect 2593 6919 2651 6925
rect 2593 6916 2605 6919
rect 2424 6888 2605 6916
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6848 1639 6851
rect 1670 6848 1676 6860
rect 1627 6820 1676 6848
rect 1627 6817 1639 6820
rect 1581 6811 1639 6817
rect 1670 6808 1676 6820
rect 1728 6808 1734 6860
rect 1765 6715 1823 6721
rect 1765 6681 1777 6715
rect 1811 6712 1823 6715
rect 2222 6712 2228 6724
rect 1811 6684 2228 6712
rect 1811 6681 1823 6684
rect 1765 6675 1823 6681
rect 2222 6672 2228 6684
rect 2280 6672 2286 6724
rect 2424 6712 2452 6888
rect 2593 6885 2605 6888
rect 2639 6885 2651 6919
rect 2593 6879 2651 6885
rect 3694 6876 3700 6928
rect 3752 6916 3758 6928
rect 4433 6919 4491 6925
rect 4433 6916 4445 6919
rect 3752 6888 4445 6916
rect 3752 6876 3758 6888
rect 4433 6885 4445 6888
rect 4479 6885 4491 6919
rect 4433 6879 4491 6885
rect 5629 6919 5687 6925
rect 5629 6885 5641 6919
rect 5675 6916 5687 6919
rect 7190 6916 7196 6928
rect 5675 6888 7196 6916
rect 5675 6885 5687 6888
rect 5629 6879 5687 6885
rect 7190 6876 7196 6888
rect 7248 6876 7254 6928
rect 7282 6876 7288 6928
rect 7340 6916 7346 6928
rect 7653 6919 7711 6925
rect 7653 6916 7665 6919
rect 7340 6888 7665 6916
rect 7340 6876 7346 6888
rect 7653 6885 7665 6888
rect 7699 6885 7711 6919
rect 7653 6879 7711 6885
rect 7742 6876 7748 6928
rect 7800 6916 7806 6928
rect 8205 6919 8263 6925
rect 8205 6916 8217 6919
rect 7800 6888 8217 6916
rect 7800 6876 7806 6888
rect 8205 6885 8217 6888
rect 8251 6885 8263 6919
rect 8205 6879 8263 6885
rect 2498 6808 2504 6860
rect 2556 6848 2562 6860
rect 3421 6851 3479 6857
rect 2556 6820 3372 6848
rect 2556 6808 2562 6820
rect 2590 6740 2596 6792
rect 2648 6780 2654 6792
rect 2685 6783 2743 6789
rect 2685 6780 2697 6783
rect 2648 6752 2697 6780
rect 2648 6740 2654 6752
rect 2685 6749 2697 6752
rect 2731 6749 2743 6783
rect 3344 6780 3372 6820
rect 3421 6817 3433 6851
rect 3467 6848 3479 6851
rect 4246 6848 4252 6860
rect 3467 6820 4252 6848
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 5534 6808 5540 6860
rect 5592 6848 5598 6860
rect 6362 6848 6368 6860
rect 5592 6820 6368 6848
rect 5592 6808 5598 6820
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 6457 6851 6515 6857
rect 6457 6817 6469 6851
rect 6503 6848 6515 6851
rect 8481 6851 8539 6857
rect 6503 6820 8156 6848
rect 6503 6817 6515 6820
rect 6457 6811 6515 6817
rect 8128 6792 8156 6820
rect 8481 6817 8493 6851
rect 8527 6848 8539 6851
rect 8570 6848 8576 6860
rect 8527 6820 8576 6848
rect 8527 6817 8539 6820
rect 8481 6811 8539 6817
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 8763 6848 8791 6956
rect 8941 6953 8953 6987
rect 8987 6984 8999 6987
rect 9214 6984 9220 6996
rect 8987 6956 9220 6984
rect 8987 6953 8999 6956
rect 8941 6947 8999 6953
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 10229 6987 10287 6993
rect 10229 6984 10241 6987
rect 9916 6956 10241 6984
rect 9916 6944 9922 6956
rect 10229 6953 10241 6956
rect 10275 6953 10287 6987
rect 10229 6947 10287 6953
rect 10321 6987 10379 6993
rect 10321 6953 10333 6987
rect 10367 6984 10379 6987
rect 10870 6984 10876 6996
rect 10367 6956 10876 6984
rect 10367 6953 10379 6956
rect 10321 6947 10379 6953
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 11238 6984 11244 6996
rect 11199 6956 11244 6984
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 11333 6987 11391 6993
rect 11333 6953 11345 6987
rect 11379 6984 11391 6987
rect 11514 6984 11520 6996
rect 11379 6956 11520 6984
rect 11379 6953 11391 6956
rect 11333 6947 11391 6953
rect 11514 6944 11520 6956
rect 11572 6944 11578 6996
rect 11606 6944 11612 6996
rect 11664 6984 11670 6996
rect 11885 6987 11943 6993
rect 11885 6984 11897 6987
rect 11664 6956 11897 6984
rect 11664 6944 11670 6956
rect 11885 6953 11897 6956
rect 11931 6953 11943 6987
rect 12802 6984 12808 6996
rect 11885 6947 11943 6953
rect 12084 6956 12808 6984
rect 11146 6916 11152 6928
rect 9048 6888 11152 6916
rect 9048 6857 9076 6888
rect 11146 6876 11152 6888
rect 11204 6876 11210 6928
rect 11532 6916 11560 6944
rect 12084 6916 12112 6956
rect 12802 6944 12808 6956
rect 12860 6944 12866 6996
rect 13265 6987 13323 6993
rect 13265 6953 13277 6987
rect 13311 6984 13323 6987
rect 13354 6984 13360 6996
rect 13311 6956 13360 6984
rect 13311 6953 13323 6956
rect 13265 6947 13323 6953
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 13722 6944 13728 6996
rect 13780 6984 13786 6996
rect 13909 6987 13967 6993
rect 13909 6984 13921 6987
rect 13780 6956 13921 6984
rect 13780 6944 13786 6956
rect 13909 6953 13921 6956
rect 13955 6953 13967 6987
rect 13909 6947 13967 6953
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 15102 6984 15108 6996
rect 14516 6956 15108 6984
rect 14516 6944 14522 6956
rect 15102 6944 15108 6956
rect 15160 6944 15166 6996
rect 15654 6984 15660 6996
rect 15615 6956 15660 6984
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 16485 6987 16543 6993
rect 16485 6953 16497 6987
rect 16531 6953 16543 6987
rect 16485 6947 16543 6953
rect 17221 6987 17279 6993
rect 17221 6953 17233 6987
rect 17267 6984 17279 6987
rect 17865 6987 17923 6993
rect 17865 6984 17877 6987
rect 17267 6956 17877 6984
rect 17267 6953 17279 6956
rect 17221 6947 17279 6953
rect 17865 6953 17877 6956
rect 17911 6953 17923 6987
rect 17865 6947 17923 6953
rect 11532 6888 12112 6916
rect 12158 6876 12164 6928
rect 12216 6916 12222 6928
rect 12253 6919 12311 6925
rect 12253 6916 12265 6919
rect 12216 6888 12265 6916
rect 12216 6876 12222 6888
rect 12253 6885 12265 6888
rect 12299 6885 12311 6919
rect 13372 6916 13400 6944
rect 15470 6916 15476 6928
rect 13372 6888 15476 6916
rect 12253 6879 12311 6885
rect 15470 6876 15476 6888
rect 15528 6876 15534 6928
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 8763 6820 9045 6848
rect 9033 6817 9045 6820
rect 9079 6817 9091 6851
rect 11882 6848 11888 6860
rect 9033 6811 9091 6817
rect 9416 6820 11888 6848
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 3344 6752 4537 6780
rect 2685 6743 2743 6749
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 5166 6780 5172 6792
rect 4755 6752 5172 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 4065 6715 4123 6721
rect 4065 6712 4077 6715
rect 2424 6684 4077 6712
rect 4065 6681 4077 6684
rect 4111 6681 4123 6715
rect 5736 6712 5764 6743
rect 5810 6740 5816 6792
rect 5868 6780 5874 6792
rect 5868 6752 5913 6780
rect 5868 6740 5874 6752
rect 6546 6740 6552 6792
rect 6604 6780 6610 6792
rect 6730 6780 6736 6792
rect 6604 6752 6649 6780
rect 6691 6752 6736 6780
rect 6604 6740 6610 6752
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 7466 6780 7472 6792
rect 7116 6752 7472 6780
rect 7116 6712 7144 6752
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6749 7803 6783
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7745 6743 7803 6749
rect 7852 6752 7941 6780
rect 7282 6712 7288 6724
rect 5736 6684 7144 6712
rect 7243 6684 7288 6712
rect 4065 6675 4123 6681
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6644 2191 6647
rect 2958 6644 2964 6656
rect 2179 6616 2964 6644
rect 2179 6613 2191 6616
rect 2133 6607 2191 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5534 6644 5540 6656
rect 5307 6616 5540 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 5626 6604 5632 6656
rect 5684 6644 5690 6656
rect 6089 6647 6147 6653
rect 6089 6644 6101 6647
rect 5684 6616 6101 6644
rect 5684 6604 5690 6616
rect 6089 6613 6101 6616
rect 6135 6613 6147 6647
rect 6089 6607 6147 6613
rect 6362 6604 6368 6656
rect 6420 6644 6426 6656
rect 6914 6644 6920 6656
rect 6420 6616 6920 6644
rect 6420 6604 6426 6616
rect 6914 6604 6920 6616
rect 6972 6644 6978 6656
rect 7101 6647 7159 6653
rect 7101 6644 7113 6647
rect 6972 6616 7113 6644
rect 6972 6604 6978 6616
rect 7101 6613 7113 6616
rect 7147 6644 7159 6647
rect 7760 6644 7788 6743
rect 7852 6724 7880 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 8938 6780 8944 6792
rect 8168 6752 8944 6780
rect 8168 6740 8174 6752
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6780 9275 6783
rect 9306 6780 9312 6792
rect 9263 6752 9312 6780
rect 9263 6749 9275 6752
rect 9217 6743 9275 6749
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 7834 6672 7840 6724
rect 7892 6672 7898 6724
rect 8205 6715 8263 6721
rect 8205 6681 8217 6715
rect 8251 6712 8263 6715
rect 9416 6712 9444 6820
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 14274 6848 14280 6860
rect 12452 6820 13584 6848
rect 14235 6820 14280 6848
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 10376 6752 10425 6780
rect 10376 6740 10382 6752
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6780 10839 6783
rect 11422 6780 11428 6792
rect 10827 6752 11428 6780
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 11606 6780 11612 6792
rect 11563 6752 11612 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 11606 6740 11612 6752
rect 11664 6780 11670 6792
rect 11974 6780 11980 6792
rect 11664 6752 11980 6780
rect 11664 6740 11670 6752
rect 11974 6740 11980 6752
rect 12032 6780 12038 6792
rect 12345 6783 12403 6789
rect 12032 6752 12204 6780
rect 12032 6740 12038 6752
rect 8251 6684 9444 6712
rect 9861 6715 9919 6721
rect 8251 6681 8263 6684
rect 8205 6675 8263 6681
rect 9861 6681 9873 6715
rect 9907 6712 9919 6715
rect 12176 6712 12204 6752
rect 12345 6749 12357 6783
rect 12391 6780 12403 6783
rect 12452 6780 12480 6820
rect 12391 6752 12480 6780
rect 12529 6783 12587 6789
rect 12391 6749 12403 6752
rect 12345 6743 12403 6749
rect 12529 6749 12541 6783
rect 12575 6749 12587 6783
rect 13354 6780 13360 6792
rect 13315 6752 13360 6780
rect 12529 6743 12587 6749
rect 12544 6712 12572 6743
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6749 13507 6783
rect 13449 6743 13507 6749
rect 9907 6684 12112 6712
rect 12176 6684 12572 6712
rect 9907 6681 9919 6684
rect 9861 6675 9919 6681
rect 8294 6644 8300 6656
rect 7147 6616 7788 6644
rect 8255 6616 8300 6644
rect 7147 6613 7159 6616
rect 7101 6607 7159 6613
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 10226 6644 10232 6656
rect 8619 6616 10232 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 10781 6647 10839 6653
rect 10781 6644 10793 6647
rect 10468 6616 10793 6644
rect 10468 6604 10474 6616
rect 10781 6613 10793 6616
rect 10827 6613 10839 6647
rect 10781 6607 10839 6613
rect 10873 6647 10931 6653
rect 10873 6613 10885 6647
rect 10919 6644 10931 6647
rect 10962 6644 10968 6656
rect 10919 6616 10968 6644
rect 10919 6613 10931 6616
rect 10873 6607 10931 6613
rect 10962 6604 10968 6616
rect 11020 6604 11026 6656
rect 12084 6644 12112 6684
rect 12618 6672 12624 6724
rect 12676 6712 12682 6724
rect 12897 6715 12955 6721
rect 12897 6712 12909 6715
rect 12676 6684 12909 6712
rect 12676 6672 12682 6684
rect 12897 6681 12909 6684
rect 12943 6681 12955 6715
rect 12897 6675 12955 6681
rect 12986 6672 12992 6724
rect 13044 6712 13050 6724
rect 13464 6712 13492 6743
rect 13044 6684 13492 6712
rect 13556 6712 13584 6820
rect 14274 6808 14280 6820
rect 14332 6808 14338 6860
rect 14752 6820 16151 6848
rect 14366 6780 14372 6792
rect 14327 6752 14372 6780
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 14516 6752 14561 6780
rect 14516 6740 14522 6752
rect 14752 6712 14780 6820
rect 15746 6780 15752 6792
rect 15707 6752 15752 6780
rect 15746 6740 15752 6752
rect 15804 6740 15810 6792
rect 15933 6783 15991 6789
rect 15933 6749 15945 6783
rect 15979 6780 15991 6783
rect 16022 6780 16028 6792
rect 15979 6752 16028 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 16123 6780 16151 6820
rect 16298 6808 16304 6860
rect 16356 6848 16362 6860
rect 16500 6848 16528 6947
rect 18046 6944 18052 6996
rect 18104 6984 18110 6996
rect 18325 6987 18383 6993
rect 18325 6984 18337 6987
rect 18104 6956 18337 6984
rect 18104 6944 18110 6956
rect 18325 6953 18337 6956
rect 18371 6953 18383 6987
rect 18325 6947 18383 6953
rect 19334 6944 19340 6996
rect 19392 6944 19398 6996
rect 18233 6919 18291 6925
rect 18233 6885 18245 6919
rect 18279 6916 18291 6919
rect 19352 6916 19380 6944
rect 18279 6888 19380 6916
rect 18279 6885 18291 6888
rect 18233 6879 18291 6885
rect 19242 6848 19248 6860
rect 16356 6820 16401 6848
rect 16500 6820 19248 6848
rect 16356 6808 16362 6820
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 19426 6857 19432 6860
rect 19420 6848 19432 6857
rect 19387 6820 19432 6848
rect 19420 6811 19432 6820
rect 19426 6808 19432 6811
rect 19484 6808 19490 6860
rect 17034 6780 17040 6792
rect 16123 6752 17040 6780
rect 17034 6740 17040 6752
rect 17092 6740 17098 6792
rect 17313 6783 17371 6789
rect 17313 6749 17325 6783
rect 17359 6749 17371 6783
rect 17494 6780 17500 6792
rect 17455 6752 17500 6780
rect 17313 6743 17371 6749
rect 13556 6684 14780 6712
rect 15289 6715 15347 6721
rect 13044 6672 13050 6684
rect 15289 6681 15301 6715
rect 15335 6712 15347 6715
rect 17328 6712 17356 6743
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6780 18567 6783
rect 18598 6780 18604 6792
rect 18555 6752 18604 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 19061 6783 19119 6789
rect 19061 6749 19073 6783
rect 19107 6780 19119 6783
rect 19150 6780 19156 6792
rect 19107 6752 19156 6780
rect 19107 6749 19119 6752
rect 19061 6743 19119 6749
rect 19150 6740 19156 6752
rect 19208 6740 19214 6792
rect 20898 6780 20904 6792
rect 20859 6752 20904 6780
rect 20898 6740 20904 6752
rect 20956 6740 20962 6792
rect 15335 6684 17356 6712
rect 15335 6681 15347 6684
rect 15289 6675 15347 6681
rect 17678 6672 17684 6724
rect 17736 6712 17742 6724
rect 17736 6684 19196 6712
rect 17736 6672 17742 6684
rect 15194 6644 15200 6656
rect 12084 6616 15200 6644
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 15378 6604 15384 6656
rect 15436 6644 15442 6656
rect 16298 6644 16304 6656
rect 15436 6616 16304 6644
rect 15436 6604 15442 6616
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 16853 6647 16911 6653
rect 16853 6613 16865 6647
rect 16899 6644 16911 6647
rect 17402 6644 17408 6656
rect 16899 6616 17408 6644
rect 16899 6613 16911 6616
rect 16853 6607 16911 6613
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 17862 6604 17868 6656
rect 17920 6644 17926 6656
rect 19061 6647 19119 6653
rect 19061 6644 19073 6647
rect 17920 6616 19073 6644
rect 17920 6604 17926 6616
rect 19061 6613 19073 6616
rect 19107 6613 19119 6647
rect 19168 6644 19196 6684
rect 20162 6672 20168 6724
rect 20220 6712 20226 6724
rect 20533 6715 20591 6721
rect 20533 6712 20545 6715
rect 20220 6684 20545 6712
rect 20220 6672 20226 6684
rect 20533 6681 20545 6684
rect 20579 6681 20591 6715
rect 20533 6675 20591 6681
rect 19426 6644 19432 6656
rect 19168 6616 19432 6644
rect 19061 6607 19119 6613
rect 19426 6604 19432 6616
rect 19484 6644 19490 6656
rect 20438 6644 20444 6656
rect 19484 6616 20444 6644
rect 19484 6604 19490 6616
rect 20438 6604 20444 6616
rect 20496 6604 20502 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 1946 6400 1952 6452
rect 2004 6440 2010 6452
rect 3605 6443 3663 6449
rect 3605 6440 3617 6443
rect 2004 6412 3617 6440
rect 2004 6400 2010 6412
rect 3605 6409 3617 6412
rect 3651 6409 3663 6443
rect 3605 6403 3663 6409
rect 5074 6400 5080 6452
rect 5132 6440 5138 6452
rect 6638 6440 6644 6452
rect 5132 6412 6644 6440
rect 5132 6400 5138 6412
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 8662 6440 8668 6452
rect 8312 6412 8668 6440
rect 3326 6372 3332 6384
rect 3287 6344 3332 6372
rect 3326 6332 3332 6344
rect 3384 6332 3390 6384
rect 4890 6372 4896 6384
rect 4851 6344 4896 6372
rect 4890 6332 4896 6344
rect 4948 6332 4954 6384
rect 5169 6375 5227 6381
rect 5169 6341 5181 6375
rect 5215 6372 5227 6375
rect 5261 6375 5319 6381
rect 5261 6372 5273 6375
rect 5215 6344 5273 6372
rect 5215 6341 5227 6344
rect 5169 6335 5227 6341
rect 5261 6341 5273 6344
rect 5307 6341 5319 6375
rect 7469 6375 7527 6381
rect 7469 6372 7481 6375
rect 5261 6335 5319 6341
rect 5368 6344 7481 6372
rect 3510 6264 3516 6316
rect 3568 6304 3574 6316
rect 4157 6307 4215 6313
rect 4157 6304 4169 6307
rect 3568 6276 4169 6304
rect 3568 6264 3574 6276
rect 4157 6273 4169 6276
rect 4203 6273 4215 6307
rect 4157 6267 4215 6273
rect 4614 6264 4620 6316
rect 4672 6304 4678 6316
rect 5368 6304 5396 6344
rect 7469 6341 7481 6344
rect 7515 6372 7527 6375
rect 7561 6375 7619 6381
rect 7561 6372 7573 6375
rect 7515 6344 7573 6372
rect 7515 6341 7527 6344
rect 7469 6335 7527 6341
rect 7561 6341 7573 6344
rect 7607 6341 7619 6375
rect 7561 6335 7619 6341
rect 4672 6276 5396 6304
rect 4672 6264 4678 6276
rect 5442 6264 5448 6316
rect 5500 6304 5506 6316
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5500 6276 5825 6304
rect 5500 6264 5506 6276
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6304 6331 6307
rect 6362 6304 6368 6316
rect 6319 6276 6368 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 6362 6264 6368 6276
rect 6420 6264 6426 6316
rect 8312 6304 8340 6412
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 8757 6443 8815 6449
rect 8757 6409 8769 6443
rect 8803 6440 8815 6443
rect 9674 6440 9680 6452
rect 8803 6412 9680 6440
rect 8803 6409 8815 6412
rect 8757 6403 8815 6409
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 9784 6412 10815 6440
rect 8478 6332 8484 6384
rect 8536 6372 8542 6384
rect 8536 6344 8708 6372
rect 8536 6332 8542 6344
rect 8680 6316 8708 6344
rect 9122 6332 9128 6384
rect 9180 6372 9186 6384
rect 9306 6372 9312 6384
rect 9180 6344 9312 6372
rect 9180 6332 9186 6344
rect 9306 6332 9312 6344
rect 9364 6372 9370 6384
rect 9784 6372 9812 6412
rect 9364 6344 9812 6372
rect 9364 6332 9370 6344
rect 7024 6276 8340 6304
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 1578 6236 1584 6248
rect 1443 6208 1584 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 1578 6196 1584 6208
rect 1636 6196 1642 6248
rect 1854 6196 1860 6248
rect 1912 6236 1918 6248
rect 1949 6239 2007 6245
rect 1949 6236 1961 6239
rect 1912 6208 1961 6236
rect 1912 6196 1918 6208
rect 1949 6205 1961 6208
rect 1995 6205 2007 6239
rect 1949 6199 2007 6205
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 4798 6236 4804 6248
rect 4755 6208 4804 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 4890 6196 4896 6248
rect 4948 6236 4954 6248
rect 5258 6236 5264 6248
rect 4948 6208 5264 6236
rect 4948 6196 4954 6208
rect 5258 6196 5264 6208
rect 5316 6196 5322 6248
rect 5626 6236 5632 6248
rect 5587 6208 5632 6236
rect 5626 6196 5632 6208
rect 5684 6196 5690 6248
rect 5721 6239 5779 6245
rect 5721 6205 5733 6239
rect 5767 6236 5779 6239
rect 6454 6236 6460 6248
rect 5767 6208 6460 6236
rect 5767 6205 5779 6208
rect 5721 6199 5779 6205
rect 6454 6196 6460 6208
rect 6512 6196 6518 6248
rect 7024 6245 7052 6276
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 8662 6304 8668 6316
rect 8444 6276 8489 6304
rect 8575 6276 8668 6304
rect 8444 6264 8450 6276
rect 8662 6264 8668 6276
rect 8720 6304 8726 6316
rect 8720 6276 9352 6304
rect 8720 6264 8726 6276
rect 7009 6239 7067 6245
rect 7009 6205 7021 6239
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6236 7527 6239
rect 8205 6239 8263 6245
rect 8205 6236 8217 6239
rect 7515 6208 8217 6236
rect 7515 6205 7527 6208
rect 7469 6199 7527 6205
rect 8205 6205 8217 6208
rect 8251 6236 8263 6239
rect 8294 6236 8300 6248
rect 8251 6208 8300 6236
rect 8251 6205 8263 6208
rect 8205 6199 8263 6205
rect 8294 6196 8300 6208
rect 8352 6196 8358 6248
rect 9214 6236 9220 6248
rect 9175 6208 9220 6236
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9324 6236 9352 6276
rect 9398 6264 9404 6316
rect 9456 6304 9462 6316
rect 9585 6307 9643 6313
rect 9585 6304 9597 6307
rect 9456 6276 9597 6304
rect 9456 6264 9462 6276
rect 9585 6273 9597 6276
rect 9631 6273 9643 6307
rect 10787 6304 10815 6412
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 12158 6440 12164 6452
rect 12032 6412 12164 6440
rect 12032 6400 12038 6412
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 14458 6440 14464 6452
rect 12268 6412 14464 6440
rect 10870 6332 10876 6384
rect 10928 6372 10934 6384
rect 12268 6372 12296 6412
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 14645 6443 14703 6449
rect 14645 6409 14657 6443
rect 14691 6440 14703 6443
rect 16853 6443 16911 6449
rect 16853 6440 16865 6443
rect 14691 6412 16865 6440
rect 14691 6409 14703 6412
rect 14645 6403 14703 6409
rect 16853 6409 16865 6412
rect 16899 6409 16911 6443
rect 16853 6403 16911 6409
rect 16945 6443 17003 6449
rect 16945 6409 16957 6443
rect 16991 6440 17003 6443
rect 18782 6440 18788 6452
rect 16991 6412 18788 6440
rect 16991 6409 17003 6412
rect 16945 6403 17003 6409
rect 18782 6400 18788 6412
rect 18840 6400 18846 6452
rect 19245 6443 19303 6449
rect 19245 6409 19257 6443
rect 19291 6440 19303 6443
rect 19518 6440 19524 6452
rect 19291 6412 19524 6440
rect 19291 6409 19303 6412
rect 19245 6403 19303 6409
rect 19518 6400 19524 6412
rect 19576 6400 19582 6452
rect 20438 6400 20444 6452
rect 20496 6440 20502 6452
rect 20717 6443 20775 6449
rect 20717 6440 20729 6443
rect 20496 6412 20729 6440
rect 20496 6400 20502 6412
rect 20717 6409 20729 6412
rect 20763 6409 20775 6443
rect 20717 6403 20775 6409
rect 13998 6372 14004 6384
rect 10928 6344 12296 6372
rect 13959 6344 14004 6372
rect 10928 6332 10934 6344
rect 13998 6332 14004 6344
rect 14056 6332 14062 6384
rect 16022 6332 16028 6384
rect 16080 6372 16086 6384
rect 16393 6375 16451 6381
rect 16393 6372 16405 6375
rect 16080 6344 16405 6372
rect 16080 6332 16086 6344
rect 16393 6341 16405 6344
rect 16439 6372 16451 6375
rect 16439 6344 18644 6372
rect 16439 6341 16451 6344
rect 16393 6335 16451 6341
rect 18616 6316 18644 6344
rect 10787 6276 12747 6304
rect 9585 6267 9643 6273
rect 9674 6236 9680 6248
rect 9324 6208 9680 6236
rect 9674 6196 9680 6208
rect 9732 6236 9738 6248
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 9732 6208 9781 6236
rect 9732 6196 9738 6208
rect 9769 6205 9781 6208
rect 9815 6205 9827 6239
rect 9769 6199 9827 6205
rect 11793 6239 11851 6245
rect 11793 6205 11805 6239
rect 11839 6236 11851 6239
rect 12342 6236 12348 6248
rect 11839 6208 12348 6236
rect 11839 6205 11851 6208
rect 11793 6199 11851 6205
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 12618 6236 12624 6248
rect 12492 6208 12624 6236
rect 12492 6196 12498 6208
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 12719 6236 12747 6276
rect 13722 6264 13728 6316
rect 13780 6304 13786 6316
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 13780 6276 15025 6304
rect 13780 6264 13786 6276
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 17402 6304 17408 6316
rect 17363 6276 17408 6304
rect 15013 6267 15071 6273
rect 17402 6264 17408 6276
rect 17460 6264 17466 6316
rect 17589 6307 17647 6313
rect 17589 6273 17601 6307
rect 17635 6304 17647 6307
rect 17678 6304 17684 6316
rect 17635 6276 17684 6304
rect 17635 6273 17647 6276
rect 17589 6267 17647 6273
rect 17678 6264 17684 6276
rect 17736 6264 17742 6316
rect 18414 6264 18420 6316
rect 18472 6304 18478 6316
rect 18509 6307 18567 6313
rect 18509 6304 18521 6307
rect 18472 6276 18521 6304
rect 18472 6264 18478 6276
rect 18509 6273 18521 6276
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 18598 6264 18604 6316
rect 18656 6304 18662 6316
rect 18656 6276 18701 6304
rect 18656 6264 18662 6276
rect 18782 6264 18788 6316
rect 18840 6304 18846 6316
rect 19150 6304 19156 6316
rect 18840 6276 19156 6304
rect 18840 6264 18846 6276
rect 19150 6264 19156 6276
rect 19208 6304 19214 6316
rect 19337 6307 19395 6313
rect 19337 6304 19349 6307
rect 19208 6276 19349 6304
rect 19208 6264 19214 6276
rect 19337 6273 19349 6276
rect 19383 6273 19395 6307
rect 19337 6267 19395 6273
rect 14274 6236 14280 6248
rect 12719 6208 14280 6236
rect 14274 6196 14280 6208
rect 14332 6196 14338 6248
rect 14458 6236 14464 6248
rect 14371 6208 14464 6236
rect 2216 6171 2274 6177
rect 2216 6137 2228 6171
rect 2262 6168 2274 6171
rect 2406 6168 2412 6180
rect 2262 6140 2412 6168
rect 2262 6137 2274 6140
rect 2216 6131 2274 6137
rect 2406 6128 2412 6140
rect 2464 6128 2470 6180
rect 4065 6171 4123 6177
rect 4065 6137 4077 6171
rect 4111 6168 4123 6171
rect 5169 6171 5227 6177
rect 5169 6168 5181 6171
rect 4111 6140 5181 6168
rect 4111 6137 4123 6140
rect 4065 6131 4123 6137
rect 5169 6137 5181 6140
rect 5215 6137 5227 6171
rect 5169 6131 5227 6137
rect 7098 6128 7104 6180
rect 7156 6168 7162 6180
rect 8113 6171 8171 6177
rect 8113 6168 8125 6171
rect 7156 6140 8125 6168
rect 7156 6128 7162 6140
rect 8113 6137 8125 6140
rect 8159 6137 8171 6171
rect 8113 6131 8171 6137
rect 10036 6171 10094 6177
rect 10036 6137 10048 6171
rect 10082 6168 10094 6171
rect 11606 6168 11612 6180
rect 10082 6140 11612 6168
rect 10082 6137 10094 6140
rect 10036 6131 10094 6137
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 3973 6103 4031 6109
rect 3973 6100 3985 6103
rect 3384 6072 3985 6100
rect 3384 6060 3390 6072
rect 3973 6069 3985 6072
rect 4019 6069 4031 6103
rect 3973 6063 4031 6069
rect 5626 6060 5632 6112
rect 5684 6100 5690 6112
rect 6178 6100 6184 6112
rect 5684 6072 6184 6100
rect 5684 6060 5690 6072
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 7193 6103 7251 6109
rect 7193 6069 7205 6103
rect 7239 6100 7251 6103
rect 7282 6100 7288 6112
rect 7239 6072 7288 6100
rect 7239 6069 7251 6072
rect 7193 6063 7251 6069
rect 7282 6060 7288 6072
rect 7340 6060 7346 6112
rect 7742 6100 7748 6112
rect 7703 6072 7748 6100
rect 7742 6060 7748 6072
rect 7800 6060 7806 6112
rect 9122 6100 9128 6112
rect 9083 6072 9128 6100
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9585 6103 9643 6109
rect 9585 6069 9597 6103
rect 9631 6100 9643 6103
rect 10051 6100 10079 6131
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 12888 6171 12946 6177
rect 12888 6137 12900 6171
rect 12934 6168 12946 6171
rect 13814 6168 13820 6180
rect 12934 6140 13820 6168
rect 12934 6137 12946 6140
rect 12888 6131 12946 6137
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 14182 6128 14188 6180
rect 14240 6168 14246 6180
rect 14384 6168 14412 6208
rect 14458 6196 14464 6208
rect 14516 6196 14522 6248
rect 15838 6196 15844 6248
rect 15896 6236 15902 6248
rect 19245 6239 19303 6245
rect 19245 6236 19257 6239
rect 15896 6208 19257 6236
rect 15896 6196 15902 6208
rect 19245 6205 19257 6208
rect 19291 6205 19303 6239
rect 19245 6199 19303 6205
rect 14240 6140 14412 6168
rect 15280 6171 15338 6177
rect 14240 6128 14246 6140
rect 15280 6137 15292 6171
rect 15326 6168 15338 6171
rect 15378 6168 15384 6180
rect 15326 6140 15384 6168
rect 15326 6137 15338 6140
rect 15280 6131 15338 6137
rect 15378 6128 15384 6140
rect 15436 6168 15442 6180
rect 15930 6168 15936 6180
rect 15436 6140 15936 6168
rect 15436 6128 15442 6140
rect 15930 6128 15936 6140
rect 15988 6128 15994 6180
rect 16853 6171 16911 6177
rect 16853 6137 16865 6171
rect 16899 6168 16911 6171
rect 18417 6171 18475 6177
rect 16899 6140 18368 6168
rect 16899 6137 16911 6140
rect 16853 6131 16911 6137
rect 9631 6072 10079 6100
rect 9631 6069 9643 6072
rect 9585 6063 9643 6069
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 11020 6072 11161 6100
rect 11020 6060 11026 6072
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 11149 6063 11207 6069
rect 11977 6103 12035 6109
rect 11977 6069 11989 6103
rect 12023 6100 12035 6103
rect 12526 6100 12532 6112
rect 12023 6072 12532 6100
rect 12023 6069 12035 6072
rect 11977 6063 12035 6069
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 12802 6060 12808 6112
rect 12860 6100 12866 6112
rect 15654 6100 15660 6112
rect 12860 6072 15660 6100
rect 12860 6060 12866 6072
rect 15654 6060 15660 6072
rect 15712 6060 15718 6112
rect 17313 6103 17371 6109
rect 17313 6069 17325 6103
rect 17359 6100 17371 6103
rect 17862 6100 17868 6112
rect 17359 6072 17868 6100
rect 17359 6069 17371 6072
rect 17313 6063 17371 6069
rect 17862 6060 17868 6072
rect 17920 6060 17926 6112
rect 18046 6100 18052 6112
rect 18007 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 18340 6100 18368 6140
rect 18417 6137 18429 6171
rect 18463 6168 18475 6171
rect 19426 6168 19432 6180
rect 18463 6140 19432 6168
rect 18463 6137 18475 6140
rect 18417 6131 18475 6137
rect 19426 6128 19432 6140
rect 19484 6128 19490 6180
rect 19604 6171 19662 6177
rect 19604 6137 19616 6171
rect 19650 6168 19662 6171
rect 20162 6168 20168 6180
rect 19650 6140 20168 6168
rect 19650 6137 19662 6140
rect 19604 6131 19662 6137
rect 20162 6128 20168 6140
rect 20220 6128 20226 6180
rect 21818 6100 21824 6112
rect 18340 6072 21824 6100
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 1762 5896 1768 5908
rect 1723 5868 1768 5896
rect 1762 5856 1768 5868
rect 1820 5856 1826 5908
rect 3970 5896 3976 5908
rect 2507 5868 3976 5896
rect 2507 5837 2535 5868
rect 3970 5856 3976 5868
rect 4028 5896 4034 5908
rect 5442 5896 5448 5908
rect 4028 5868 5448 5896
rect 4028 5856 4034 5868
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 5644 5868 7021 5896
rect 2492 5831 2550 5837
rect 2492 5797 2504 5831
rect 2538 5797 2550 5831
rect 2492 5791 2550 5797
rect 4246 5788 4252 5840
rect 4304 5828 4310 5840
rect 5644 5828 5672 5868
rect 7009 5865 7021 5868
rect 7055 5865 7067 5899
rect 7190 5896 7196 5908
rect 7151 5868 7196 5896
rect 7009 5859 7067 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 7466 5856 7472 5908
rect 7524 5896 7530 5908
rect 8205 5899 8263 5905
rect 8205 5896 8217 5899
rect 7524 5868 8217 5896
rect 7524 5856 7530 5868
rect 8205 5865 8217 5868
rect 8251 5865 8263 5899
rect 12342 5896 12348 5908
rect 8205 5859 8263 5865
rect 8404 5868 12348 5896
rect 4304 5800 5672 5828
rect 5721 5831 5779 5837
rect 4304 5788 4310 5800
rect 5721 5797 5733 5831
rect 5767 5828 5779 5831
rect 7561 5831 7619 5837
rect 7561 5828 7573 5831
rect 5767 5800 7573 5828
rect 5767 5797 5779 5800
rect 5721 5791 5779 5797
rect 7561 5797 7573 5800
rect 7607 5797 7619 5831
rect 7561 5791 7619 5797
rect 8113 5831 8171 5837
rect 8113 5797 8125 5831
rect 8159 5828 8171 5831
rect 8404 5828 8432 5868
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 14090 5896 14096 5908
rect 12492 5868 14096 5896
rect 12492 5856 12498 5868
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 14182 5856 14188 5908
rect 14240 5896 14246 5908
rect 14461 5899 14519 5905
rect 14461 5896 14473 5899
rect 14240 5868 14473 5896
rect 14240 5856 14246 5868
rect 14461 5865 14473 5868
rect 14507 5865 14519 5899
rect 14461 5859 14519 5865
rect 14737 5899 14795 5905
rect 14737 5865 14749 5899
rect 14783 5896 14795 5899
rect 15010 5896 15016 5908
rect 14783 5868 15016 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 15841 5899 15899 5905
rect 15841 5865 15853 5899
rect 15887 5896 15899 5899
rect 16206 5896 16212 5908
rect 15887 5868 16212 5896
rect 15887 5865 15899 5868
rect 15841 5859 15899 5865
rect 16206 5856 16212 5868
rect 16264 5856 16270 5908
rect 17954 5896 17960 5908
rect 16684 5868 17960 5896
rect 8570 5828 8576 5840
rect 8159 5800 8432 5828
rect 8531 5800 8576 5828
rect 8159 5797 8171 5800
rect 8113 5791 8171 5797
rect 8570 5788 8576 5800
rect 8628 5788 8634 5840
rect 8665 5831 8723 5837
rect 8665 5797 8677 5831
rect 8711 5797 8723 5831
rect 8665 5791 8723 5797
rect 9944 5831 10002 5837
rect 9944 5797 9956 5831
rect 9990 5828 10002 5831
rect 10502 5828 10508 5840
rect 9990 5800 10508 5828
rect 9990 5797 10002 5800
rect 9944 5791 10002 5797
rect 4332 5763 4390 5769
rect 4332 5729 4344 5763
rect 4378 5760 4390 5763
rect 5074 5760 5080 5772
rect 4378 5732 5080 5760
rect 4378 5729 4390 5732
rect 4332 5723 4390 5729
rect 5074 5720 5080 5732
rect 5132 5720 5138 5772
rect 6546 5760 6552 5772
rect 6507 5732 6552 5760
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 6641 5763 6699 5769
rect 6641 5729 6653 5763
rect 6687 5760 6699 5763
rect 7282 5760 7288 5772
rect 6687 5732 7288 5760
rect 6687 5729 6699 5732
rect 6641 5723 6699 5729
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 8680 5760 8708 5791
rect 10502 5788 10508 5800
rect 10560 5828 10566 5840
rect 10962 5828 10968 5840
rect 10560 5800 10968 5828
rect 10560 5788 10566 5800
rect 10962 5788 10968 5800
rect 11020 5788 11026 5840
rect 11793 5831 11851 5837
rect 11793 5797 11805 5831
rect 11839 5828 11851 5831
rect 11882 5828 11888 5840
rect 11839 5800 11888 5828
rect 11839 5797 11851 5800
rect 11793 5791 11851 5797
rect 11882 5788 11888 5800
rect 11940 5788 11946 5840
rect 12986 5828 12992 5840
rect 11992 5800 12992 5828
rect 8938 5760 8944 5772
rect 7383 5732 8944 5760
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 6822 5692 6828 5704
rect 6783 5664 6828 5692
rect 4065 5655 4123 5661
rect 1854 5516 1860 5568
rect 1912 5556 1918 5568
rect 2240 5556 2268 5655
rect 4080 5624 4108 5655
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 7383 5692 7411 5732
rect 8938 5720 8944 5732
rect 8996 5720 9002 5772
rect 9674 5760 9680 5772
rect 9635 5732 9680 5760
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 9766 5720 9772 5772
rect 9824 5760 9830 5772
rect 11698 5760 11704 5772
rect 9824 5732 11275 5760
rect 11659 5732 11704 5760
rect 9824 5720 9830 5732
rect 6932 5664 7411 5692
rect 7653 5695 7711 5701
rect 3436 5596 4108 5624
rect 3436 5556 3464 5596
rect 6730 5584 6736 5636
rect 6788 5624 6794 5636
rect 6932 5624 6960 5664
rect 7653 5661 7665 5695
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5692 7895 5695
rect 8386 5692 8392 5704
rect 7883 5664 8392 5692
rect 7883 5661 7895 5664
rect 7837 5655 7895 5661
rect 6788 5596 6960 5624
rect 6788 5584 6794 5596
rect 7466 5584 7472 5636
rect 7524 5624 7530 5636
rect 7668 5624 7696 5655
rect 8386 5652 8392 5664
rect 8444 5692 8450 5704
rect 8757 5695 8815 5701
rect 8757 5692 8769 5695
rect 8444 5664 8769 5692
rect 8444 5652 8450 5664
rect 8757 5661 8769 5664
rect 8803 5661 8815 5695
rect 9306 5692 9312 5704
rect 8757 5655 8815 5661
rect 8864 5664 9312 5692
rect 7524 5596 7696 5624
rect 7524 5584 7530 5596
rect 7742 5584 7748 5636
rect 7800 5624 7806 5636
rect 8113 5627 8171 5633
rect 8113 5624 8125 5627
rect 7800 5596 8125 5624
rect 7800 5584 7806 5596
rect 8113 5593 8125 5596
rect 8159 5593 8171 5627
rect 8113 5587 8171 5593
rect 8294 5584 8300 5636
rect 8352 5624 8358 5636
rect 8864 5624 8892 5664
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 10962 5652 10968 5704
rect 11020 5692 11026 5704
rect 11146 5692 11152 5704
rect 11020 5664 11152 5692
rect 11020 5652 11026 5664
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 11247 5692 11275 5732
rect 11698 5720 11704 5732
rect 11756 5720 11762 5772
rect 11992 5760 12020 5800
rect 12986 5788 12992 5800
rect 13044 5788 13050 5840
rect 13348 5831 13406 5837
rect 13348 5797 13360 5831
rect 13394 5828 13406 5831
rect 13998 5828 14004 5840
rect 13394 5800 14004 5828
rect 13394 5797 13406 5800
rect 13348 5791 13406 5797
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 11808 5732 12020 5760
rect 11808 5692 11836 5732
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12529 5763 12587 5769
rect 12529 5760 12541 5763
rect 12492 5732 12541 5760
rect 12492 5720 12498 5732
rect 12529 5729 12541 5732
rect 12575 5729 12587 5763
rect 12529 5723 12587 5729
rect 16390 5720 16396 5772
rect 16448 5760 16454 5772
rect 16684 5769 16712 5868
rect 17954 5856 17960 5868
rect 18012 5856 18018 5908
rect 18046 5856 18052 5908
rect 18104 5896 18110 5908
rect 18509 5899 18567 5905
rect 18509 5896 18521 5899
rect 18104 5868 18521 5896
rect 18104 5856 18110 5868
rect 18509 5865 18521 5868
rect 18555 5865 18567 5899
rect 19334 5896 19340 5908
rect 19295 5868 19340 5896
rect 18509 5859 18567 5865
rect 19334 5856 19340 5868
rect 19392 5856 19398 5908
rect 19426 5856 19432 5908
rect 19484 5896 19490 5908
rect 20349 5899 20407 5905
rect 20349 5896 20361 5899
rect 19484 5868 20361 5896
rect 19484 5856 19490 5868
rect 20349 5865 20361 5868
rect 20395 5865 20407 5899
rect 20349 5859 20407 5865
rect 18601 5831 18659 5837
rect 18601 5828 18613 5831
rect 16776 5800 18613 5828
rect 16669 5763 16727 5769
rect 16669 5760 16681 5763
rect 16448 5732 16681 5760
rect 16448 5720 16454 5732
rect 16669 5729 16681 5732
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 11247 5664 11836 5692
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5692 12035 5695
rect 12250 5692 12256 5704
rect 12023 5664 12256 5692
rect 12023 5661 12035 5664
rect 11977 5655 12035 5661
rect 12250 5652 12256 5664
rect 12308 5652 12314 5704
rect 13081 5695 13139 5701
rect 13081 5692 13093 5695
rect 12544 5664 13093 5692
rect 12544 5636 12572 5664
rect 13081 5661 13093 5664
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 14826 5652 14832 5704
rect 14884 5692 14890 5704
rect 15933 5695 15991 5701
rect 15933 5692 15945 5695
rect 14884 5664 15945 5692
rect 14884 5652 14890 5664
rect 15933 5661 15945 5664
rect 15979 5661 15991 5695
rect 15933 5655 15991 5661
rect 16022 5652 16028 5704
rect 16080 5692 16086 5704
rect 16776 5692 16804 5800
rect 18601 5797 18613 5800
rect 18647 5797 18659 5831
rect 18601 5791 18659 5797
rect 16936 5763 16994 5769
rect 16936 5729 16948 5763
rect 16982 5760 16994 5763
rect 17494 5760 17500 5772
rect 16982 5732 17500 5760
rect 16982 5729 16994 5732
rect 16936 5723 16994 5729
rect 17494 5720 17500 5732
rect 17552 5760 17558 5772
rect 17552 5732 18092 5760
rect 17552 5720 17558 5732
rect 17954 5692 17960 5704
rect 16080 5664 16125 5692
rect 16684 5664 16804 5692
rect 17696 5664 17960 5692
rect 16080 5652 16086 5664
rect 9674 5624 9680 5636
rect 8352 5596 8892 5624
rect 8956 5596 9680 5624
rect 8352 5584 8358 5596
rect 1912 5528 3464 5556
rect 1912 5516 1918 5528
rect 3510 5516 3516 5568
rect 3568 5556 3574 5568
rect 3605 5559 3663 5565
rect 3605 5556 3617 5559
rect 3568 5528 3617 5556
rect 3568 5516 3574 5528
rect 3605 5525 3617 5528
rect 3651 5525 3663 5559
rect 3605 5519 3663 5525
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 6086 5556 6092 5568
rect 4120 5528 6092 5556
rect 4120 5516 4126 5528
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 6181 5559 6239 5565
rect 6181 5525 6193 5559
rect 6227 5556 6239 5559
rect 6914 5556 6920 5568
rect 6227 5528 6920 5556
rect 6227 5525 6239 5528
rect 6181 5519 6239 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 7009 5559 7067 5565
rect 7009 5525 7021 5559
rect 7055 5556 7067 5559
rect 8956 5556 8984 5596
rect 9674 5584 9680 5596
rect 9732 5584 9738 5636
rect 10686 5584 10692 5636
rect 10744 5624 10750 5636
rect 12434 5624 12440 5636
rect 10744 5596 12440 5624
rect 10744 5584 10750 5596
rect 12434 5584 12440 5596
rect 12492 5584 12498 5636
rect 12526 5584 12532 5636
rect 12584 5584 12590 5636
rect 15473 5627 15531 5633
rect 12636 5596 13124 5624
rect 7055 5528 8984 5556
rect 7055 5525 7067 5528
rect 7009 5519 7067 5525
rect 9582 5516 9588 5568
rect 9640 5556 9646 5568
rect 10318 5556 10324 5568
rect 9640 5528 10324 5556
rect 9640 5516 9646 5528
rect 10318 5516 10324 5528
rect 10376 5556 10382 5568
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 10376 5528 11069 5556
rect 10376 5516 10382 5528
rect 11057 5525 11069 5528
rect 11103 5525 11115 5559
rect 11057 5519 11115 5525
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 11204 5528 11345 5556
rect 11204 5516 11210 5528
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 11333 5519 11391 5525
rect 12342 5516 12348 5568
rect 12400 5556 12406 5568
rect 12636 5556 12664 5596
rect 12400 5528 12664 5556
rect 12713 5559 12771 5565
rect 12400 5516 12406 5528
rect 12713 5525 12725 5559
rect 12759 5556 12771 5559
rect 12802 5556 12808 5568
rect 12759 5528 12808 5556
rect 12759 5525 12771 5528
rect 12713 5519 12771 5525
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 13096 5556 13124 5596
rect 15473 5593 15485 5627
rect 15519 5624 15531 5627
rect 16684 5624 16712 5664
rect 17696 5624 17724 5664
rect 17954 5652 17960 5664
rect 18012 5652 18018 5704
rect 18064 5692 18092 5732
rect 18138 5720 18144 5772
rect 18196 5760 18202 5772
rect 19153 5763 19211 5769
rect 19153 5760 19165 5763
rect 18196 5732 19165 5760
rect 18196 5720 18202 5732
rect 19153 5729 19165 5732
rect 19199 5760 19211 5763
rect 19705 5763 19763 5769
rect 19705 5760 19717 5763
rect 19199 5732 19717 5760
rect 19199 5729 19211 5732
rect 19153 5723 19211 5729
rect 19705 5729 19717 5732
rect 19751 5729 19763 5763
rect 19705 5723 19763 5729
rect 19797 5763 19855 5769
rect 19797 5729 19809 5763
rect 19843 5760 19855 5763
rect 20990 5760 20996 5772
rect 19843 5732 20996 5760
rect 19843 5729 19855 5732
rect 19797 5723 19855 5729
rect 18693 5695 18751 5701
rect 18693 5692 18705 5695
rect 18064 5664 18705 5692
rect 18693 5661 18705 5664
rect 18739 5661 18751 5695
rect 18693 5655 18751 5661
rect 15519 5596 16712 5624
rect 17604 5596 17724 5624
rect 15519 5593 15531 5596
rect 15473 5587 15531 5593
rect 14550 5556 14556 5568
rect 13096 5528 14556 5556
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 14642 5516 14648 5568
rect 14700 5556 14706 5568
rect 17604 5556 17632 5596
rect 17862 5584 17868 5636
rect 17920 5624 17926 5636
rect 18141 5627 18199 5633
rect 18141 5624 18153 5627
rect 17920 5596 18153 5624
rect 17920 5584 17926 5596
rect 18141 5593 18153 5596
rect 18187 5593 18199 5627
rect 18141 5587 18199 5593
rect 19702 5584 19708 5636
rect 19760 5624 19766 5636
rect 19812 5624 19840 5723
rect 20990 5720 20996 5732
rect 21048 5720 21054 5772
rect 19978 5692 19984 5704
rect 19939 5664 19984 5692
rect 19978 5652 19984 5664
rect 20036 5652 20042 5704
rect 19760 5596 19840 5624
rect 19760 5584 19766 5596
rect 14700 5528 17632 5556
rect 14700 5516 14706 5528
rect 17678 5516 17684 5568
rect 17736 5556 17742 5568
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 17736 5528 18061 5556
rect 17736 5516 17742 5528
rect 18049 5525 18061 5528
rect 18095 5525 18107 5559
rect 18049 5519 18107 5525
rect 18690 5516 18696 5568
rect 18748 5556 18754 5568
rect 20070 5556 20076 5568
rect 18748 5528 20076 5556
rect 18748 5516 18754 5528
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 3326 5352 3332 5364
rect 3287 5324 3332 5352
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 7190 5352 7196 5364
rect 5767 5324 7196 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 8202 5352 8208 5364
rect 8163 5324 8208 5352
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 9490 5312 9496 5364
rect 9548 5352 9554 5364
rect 9548 5324 9720 5352
rect 9548 5312 9554 5324
rect 6641 5287 6699 5293
rect 6641 5284 6653 5287
rect 6380 5256 6653 5284
rect 1578 5216 1584 5228
rect 1539 5188 1584 5216
rect 1578 5176 1584 5188
rect 1636 5176 1642 5228
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 2958 5216 2964 5228
rect 2731 5188 2964 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 3970 5216 3976 5228
rect 3931 5188 3976 5216
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4614 5176 4620 5228
rect 4672 5216 4678 5228
rect 4985 5219 5043 5225
rect 4985 5216 4997 5219
rect 4672 5188 4997 5216
rect 4672 5176 4678 5188
rect 4985 5185 4997 5188
rect 5031 5216 5043 5219
rect 5074 5216 5080 5228
rect 5031 5188 5080 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 6380 5225 6408 5256
rect 6641 5253 6653 5256
rect 6687 5284 6699 5287
rect 6822 5284 6828 5296
rect 6687 5256 6828 5284
rect 6687 5253 6699 5256
rect 6641 5247 6699 5253
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 9692 5284 9720 5324
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 10134 5352 10140 5364
rect 9824 5324 10140 5352
rect 9824 5312 9830 5324
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10321 5355 10379 5361
rect 10321 5321 10333 5355
rect 10367 5352 10379 5355
rect 13538 5352 13544 5364
rect 10367 5324 13544 5352
rect 10367 5321 10379 5324
rect 10321 5315 10379 5321
rect 13538 5312 13544 5324
rect 13596 5312 13602 5364
rect 14737 5355 14795 5361
rect 14737 5321 14749 5355
rect 14783 5352 14795 5355
rect 14826 5352 14832 5364
rect 14783 5324 14832 5352
rect 14783 5321 14795 5324
rect 14737 5315 14795 5321
rect 14826 5312 14832 5324
rect 14884 5312 14890 5364
rect 15930 5352 15936 5364
rect 15764 5324 15936 5352
rect 10597 5287 10655 5293
rect 9692 5256 9996 5284
rect 9968 5228 9996 5256
rect 10597 5253 10609 5287
rect 10643 5284 10655 5287
rect 10643 5256 11652 5284
rect 10643 5253 10655 5256
rect 10597 5247 10655 5253
rect 6365 5219 6423 5225
rect 5316 5188 6316 5216
rect 5316 5176 5322 5188
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5108 1458 5160
rect 3234 5108 3240 5160
rect 3292 5148 3298 5160
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 3292 5120 4813 5148
rect 3292 5108 3298 5120
rect 4801 5117 4813 5120
rect 4847 5117 4859 5151
rect 4801 5111 4859 5117
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 6089 5151 6147 5157
rect 6089 5148 6101 5151
rect 5592 5120 6101 5148
rect 5592 5108 5598 5120
rect 6089 5117 6101 5120
rect 6135 5117 6147 5151
rect 6288 5148 6316 5188
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6564 5188 6960 5216
rect 6564 5148 6592 5188
rect 6288 5120 6592 5148
rect 6089 5111 6147 5117
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6788 5120 6837 5148
rect 6788 5108 6794 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6932 5148 6960 5188
rect 9950 5176 9956 5228
rect 10008 5216 10014 5228
rect 10870 5216 10876 5228
rect 10008 5188 10876 5216
rect 10008 5176 10014 5188
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 11146 5176 11152 5228
rect 11204 5216 11210 5228
rect 11425 5219 11483 5225
rect 11425 5216 11437 5219
rect 11204 5188 11437 5216
rect 11204 5176 11210 5188
rect 11425 5185 11437 5188
rect 11471 5185 11483 5219
rect 11425 5179 11483 5185
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5185 11575 5219
rect 11624 5216 11652 5256
rect 11698 5244 11704 5296
rect 11756 5284 11762 5296
rect 12250 5284 12256 5296
rect 11756 5256 12256 5284
rect 11756 5244 11762 5256
rect 12250 5244 12256 5256
rect 12308 5284 12314 5296
rect 13357 5287 13415 5293
rect 12308 5256 13124 5284
rect 12308 5244 12314 5256
rect 12802 5216 12808 5228
rect 11624 5188 12808 5216
rect 11517 5179 11575 5185
rect 8570 5148 8576 5160
rect 6932 5120 8576 5148
rect 6825 5111 6883 5117
rect 8570 5108 8576 5120
rect 8628 5108 8634 5160
rect 8662 5108 8668 5160
rect 8720 5148 8726 5160
rect 8757 5151 8815 5157
rect 8757 5148 8769 5151
rect 8720 5120 8769 5148
rect 8720 5108 8726 5120
rect 8757 5117 8769 5120
rect 8803 5117 8815 5151
rect 8757 5111 8815 5117
rect 9024 5151 9082 5157
rect 9024 5117 9036 5151
rect 9070 5148 9082 5151
rect 9582 5148 9588 5160
rect 9070 5120 9588 5148
rect 9070 5117 9082 5120
rect 9024 5111 9082 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 10321 5151 10379 5157
rect 10321 5117 10333 5151
rect 10367 5148 10379 5151
rect 10413 5151 10471 5157
rect 10413 5148 10425 5151
rect 10367 5120 10425 5148
rect 10367 5117 10379 5120
rect 10321 5111 10379 5117
rect 10413 5117 10425 5120
rect 10459 5117 10471 5151
rect 10413 5111 10471 5117
rect 10686 5108 10692 5160
rect 10744 5148 10750 5160
rect 11532 5148 11560 5179
rect 12802 5176 12808 5188
rect 12860 5176 12866 5228
rect 13096 5225 13124 5256
rect 13357 5253 13369 5287
rect 13403 5284 13415 5287
rect 13449 5287 13507 5293
rect 13449 5284 13461 5287
rect 13403 5256 13461 5284
rect 13403 5253 13415 5256
rect 13357 5247 13415 5253
rect 13449 5253 13461 5256
rect 13495 5284 13507 5287
rect 15286 5284 15292 5296
rect 13495 5256 15292 5284
rect 13495 5253 13507 5256
rect 13449 5247 13507 5253
rect 15286 5244 15292 5256
rect 15344 5244 15350 5296
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 14182 5216 14188 5228
rect 13127 5188 14188 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 14366 5176 14372 5228
rect 14424 5216 14430 5228
rect 15197 5219 15255 5225
rect 15197 5216 15209 5219
rect 14424 5188 15209 5216
rect 14424 5176 14430 5188
rect 15197 5185 15209 5188
rect 15243 5185 15255 5219
rect 15378 5216 15384 5228
rect 15339 5188 15384 5216
rect 15197 5179 15255 5185
rect 15378 5176 15384 5188
rect 15436 5176 15442 5228
rect 15764 5225 15792 5324
rect 15930 5312 15936 5324
rect 15988 5352 15994 5364
rect 16390 5352 16396 5364
rect 15988 5324 16396 5352
rect 15988 5312 15994 5324
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 17129 5355 17187 5361
rect 17129 5321 17141 5355
rect 17175 5352 17187 5355
rect 17494 5352 17500 5364
rect 17175 5324 17500 5352
rect 17175 5321 17187 5324
rect 17129 5315 17187 5321
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 18966 5312 18972 5364
rect 19024 5352 19030 5364
rect 19978 5352 19984 5364
rect 19024 5324 19984 5352
rect 19024 5312 19030 5324
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 20162 5352 20168 5364
rect 20123 5324 20168 5352
rect 20162 5312 20168 5324
rect 20220 5312 20226 5364
rect 16942 5244 16948 5296
rect 17000 5284 17006 5296
rect 17589 5287 17647 5293
rect 17589 5284 17601 5287
rect 17000 5256 17601 5284
rect 17000 5244 17006 5256
rect 17589 5253 17601 5256
rect 17635 5253 17647 5287
rect 17589 5247 17647 5253
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5185 15807 5219
rect 18782 5216 18788 5228
rect 18743 5188 18788 5216
rect 15749 5179 15807 5185
rect 18782 5176 18788 5188
rect 18840 5176 18846 5228
rect 19794 5176 19800 5228
rect 19852 5216 19858 5228
rect 20625 5219 20683 5225
rect 20625 5216 20637 5219
rect 19852 5188 20637 5216
rect 19852 5176 19858 5188
rect 20625 5185 20637 5188
rect 20671 5185 20683 5219
rect 20625 5179 20683 5185
rect 11882 5148 11888 5160
rect 10744 5120 11468 5148
rect 11532 5120 11888 5148
rect 10744 5108 10750 5120
rect 3697 5083 3755 5089
rect 3697 5049 3709 5083
rect 3743 5080 3755 5083
rect 3743 5052 4384 5080
rect 3743 5049 3755 5052
rect 3697 5043 3755 5049
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 2498 5012 2504 5024
rect 2459 4984 2504 5012
rect 2498 4972 2504 4984
rect 2556 4972 2562 5024
rect 2590 4972 2596 5024
rect 2648 5012 2654 5024
rect 3789 5015 3847 5021
rect 2648 4984 2693 5012
rect 2648 4972 2654 4984
rect 3789 4981 3801 5015
rect 3835 5012 3847 5015
rect 4062 5012 4068 5024
rect 3835 4984 4068 5012
rect 3835 4981 3847 4984
rect 3789 4975 3847 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4356 5021 4384 5052
rect 5718 5040 5724 5092
rect 5776 5080 5782 5092
rect 6641 5083 6699 5089
rect 5776 5052 6316 5080
rect 5776 5040 5782 5052
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 4981 4399 5015
rect 4706 5012 4712 5024
rect 4667 4984 4712 5012
rect 4341 4975 4399 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 6178 5012 6184 5024
rect 6139 4984 6184 5012
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 6288 5012 6316 5052
rect 6641 5049 6653 5083
rect 6687 5080 6699 5083
rect 7070 5083 7128 5089
rect 7070 5080 7082 5083
rect 6687 5052 7082 5080
rect 6687 5049 6699 5052
rect 6641 5043 6699 5049
rect 7070 5049 7082 5052
rect 7116 5049 7128 5083
rect 7070 5043 7128 5049
rect 7558 5040 7564 5092
rect 7616 5080 7622 5092
rect 7616 5052 9168 5080
rect 7616 5040 7622 5052
rect 8570 5012 8576 5024
rect 6288 4984 8576 5012
rect 8570 4972 8576 4984
rect 8628 4972 8634 5024
rect 9140 5012 9168 5052
rect 9214 5040 9220 5092
rect 9272 5080 9278 5092
rect 10226 5080 10232 5092
rect 9272 5052 10232 5080
rect 9272 5040 9278 5052
rect 10226 5040 10232 5052
rect 10284 5040 10290 5092
rect 10502 5040 10508 5092
rect 10560 5080 10566 5092
rect 11333 5083 11391 5089
rect 11333 5080 11345 5083
rect 10560 5052 11345 5080
rect 10560 5040 10566 5052
rect 11333 5049 11345 5052
rect 11379 5049 11391 5083
rect 11440 5080 11468 5120
rect 11882 5108 11888 5120
rect 11940 5108 11946 5160
rect 12250 5108 12256 5160
rect 12308 5148 12314 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12308 5120 12909 5148
rect 12308 5108 12314 5120
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5148 14059 5151
rect 15010 5148 15016 5160
rect 14047 5120 15016 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 15010 5108 15016 5120
rect 15068 5108 15074 5160
rect 16022 5157 16028 5160
rect 16016 5148 16028 5157
rect 15983 5120 16028 5148
rect 16016 5111 16028 5120
rect 16022 5108 16028 5111
rect 16080 5108 16086 5160
rect 17218 5148 17224 5160
rect 16123 5120 17224 5148
rect 11974 5080 11980 5092
rect 11440 5052 11980 5080
rect 11333 5043 11391 5049
rect 11974 5040 11980 5052
rect 12032 5040 12038 5092
rect 12986 5040 12992 5092
rect 13044 5080 13050 5092
rect 14093 5083 14151 5089
rect 14093 5080 14105 5083
rect 13044 5052 14105 5080
rect 13044 5040 13050 5052
rect 14093 5049 14105 5052
rect 14139 5049 14151 5083
rect 14093 5043 14151 5049
rect 9858 5012 9864 5024
rect 9140 4984 9864 5012
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 9950 4972 9956 5024
rect 10008 5012 10014 5024
rect 10137 5015 10195 5021
rect 10137 5012 10149 5015
rect 10008 4984 10149 5012
rect 10008 4972 10014 4984
rect 10137 4981 10149 4984
rect 10183 4981 10195 5015
rect 10137 4975 10195 4981
rect 10965 5015 11023 5021
rect 10965 4981 10977 5015
rect 11011 5012 11023 5015
rect 11422 5012 11428 5024
rect 11011 4984 11428 5012
rect 11011 4981 11023 4984
rect 10965 4975 11023 4981
rect 11422 4972 11428 4984
rect 11480 4972 11486 5024
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12805 5015 12863 5021
rect 12492 4984 12537 5012
rect 12492 4972 12498 4984
rect 12805 4981 12817 5015
rect 12851 5012 12863 5015
rect 12894 5012 12900 5024
rect 12851 4984 12900 5012
rect 12851 4981 12863 4984
rect 12805 4975 12863 4981
rect 12894 4972 12900 4984
rect 12952 5012 12958 5024
rect 13449 5015 13507 5021
rect 13449 5012 13461 5015
rect 12952 4984 13461 5012
rect 12952 4972 12958 4984
rect 13449 4981 13461 4984
rect 13495 4981 13507 5015
rect 13449 4975 13507 4981
rect 13633 5015 13691 5021
rect 13633 4981 13645 5015
rect 13679 5012 13691 5015
rect 13814 5012 13820 5024
rect 13679 4984 13820 5012
rect 13679 4981 13691 4984
rect 13633 4975 13691 4981
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 14108 5012 14136 5043
rect 14366 5040 14372 5092
rect 14424 5080 14430 5092
rect 15105 5083 15163 5089
rect 15105 5080 15117 5083
rect 14424 5052 15117 5080
rect 14424 5040 14430 5052
rect 15105 5049 15117 5052
rect 15151 5049 15163 5083
rect 15105 5043 15163 5049
rect 15286 5040 15292 5092
rect 15344 5080 15350 5092
rect 16123 5080 16151 5120
rect 17218 5108 17224 5120
rect 17276 5108 17282 5160
rect 17402 5148 17408 5160
rect 17363 5120 17408 5148
rect 17402 5108 17408 5120
rect 17460 5108 17466 5160
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 20438 5148 20444 5160
rect 20399 5120 20444 5148
rect 18049 5111 18107 5117
rect 15344 5052 16151 5080
rect 15344 5040 15350 5052
rect 16298 5040 16304 5092
rect 16356 5080 16362 5092
rect 18064 5080 18092 5111
rect 20438 5108 20444 5120
rect 20496 5108 20502 5160
rect 16356 5052 18092 5080
rect 18325 5083 18383 5089
rect 16356 5040 16362 5052
rect 18325 5049 18337 5083
rect 18371 5049 18383 5083
rect 18325 5043 18383 5049
rect 19052 5083 19110 5089
rect 19052 5049 19064 5083
rect 19098 5080 19110 5083
rect 19886 5080 19892 5092
rect 19098 5052 19892 5080
rect 19098 5049 19110 5052
rect 19052 5043 19110 5049
rect 15838 5012 15844 5024
rect 14108 4984 15844 5012
rect 15838 4972 15844 4984
rect 15896 4972 15902 5024
rect 18340 5012 18368 5043
rect 19886 5040 19892 5052
rect 19944 5040 19950 5092
rect 19242 5012 19248 5024
rect 18340 4984 19248 5012
rect 19242 4972 19248 4984
rect 19300 4972 19306 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 2406 4768 2412 4820
rect 2464 4808 2470 4820
rect 2682 4808 2688 4820
rect 2464 4780 2688 4808
rect 2464 4768 2470 4780
rect 2682 4768 2688 4780
rect 2740 4808 2746 4820
rect 2869 4811 2927 4817
rect 2869 4808 2881 4811
rect 2740 4780 2881 4808
rect 2740 4768 2746 4780
rect 2869 4777 2881 4780
rect 2915 4777 2927 4811
rect 2869 4771 2927 4777
rect 3418 4768 3424 4820
rect 3476 4808 3482 4820
rect 3605 4811 3663 4817
rect 3605 4808 3617 4811
rect 3476 4780 3617 4808
rect 3476 4768 3482 4780
rect 3605 4777 3617 4780
rect 3651 4777 3663 4811
rect 4062 4808 4068 4820
rect 4023 4780 4068 4808
rect 3605 4771 3663 4777
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 4525 4811 4583 4817
rect 4525 4777 4537 4811
rect 4571 4808 4583 4811
rect 6638 4808 6644 4820
rect 4571 4780 6644 4808
rect 4571 4777 4583 4780
rect 4525 4771 4583 4777
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 7009 4811 7067 4817
rect 7009 4808 7021 4811
rect 6880 4780 7021 4808
rect 6880 4768 6886 4780
rect 7009 4777 7021 4780
rect 7055 4777 7067 4811
rect 7282 4808 7288 4820
rect 7243 4780 7288 4808
rect 7009 4771 7067 4777
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 7650 4808 7656 4820
rect 7611 4780 7656 4808
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 7745 4811 7803 4817
rect 7745 4777 7757 4811
rect 7791 4808 7803 4811
rect 8297 4811 8355 4817
rect 8297 4808 8309 4811
rect 7791 4780 8309 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 8297 4777 8309 4780
rect 8343 4777 8355 4811
rect 8297 4771 8355 4777
rect 8570 4768 8576 4820
rect 8628 4808 8634 4820
rect 8665 4811 8723 4817
rect 8665 4808 8677 4811
rect 8628 4780 8677 4808
rect 8628 4768 8634 4780
rect 8665 4777 8677 4780
rect 8711 4808 8723 4811
rect 10229 4811 10287 4817
rect 10229 4808 10241 4811
rect 8711 4780 10241 4808
rect 8711 4777 8723 4780
rect 8665 4771 8723 4777
rect 10229 4777 10241 4780
rect 10275 4777 10287 4811
rect 10229 4771 10287 4777
rect 10413 4811 10471 4817
rect 10413 4777 10425 4811
rect 10459 4808 10471 4811
rect 10502 4808 10508 4820
rect 10459 4780 10508 4808
rect 10459 4777 10471 4780
rect 10413 4771 10471 4777
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 10686 4768 10692 4820
rect 10744 4808 10750 4820
rect 10873 4811 10931 4817
rect 10873 4808 10885 4811
rect 10744 4780 10885 4808
rect 10744 4768 10750 4780
rect 10873 4777 10885 4780
rect 10919 4777 10931 4811
rect 10873 4771 10931 4777
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 11793 4811 11851 4817
rect 11793 4808 11805 4811
rect 11480 4780 11805 4808
rect 11480 4768 11486 4780
rect 11793 4777 11805 4780
rect 11839 4777 11851 4811
rect 11793 4771 11851 4777
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 12897 4811 12955 4817
rect 12897 4808 12909 4811
rect 12492 4780 12909 4808
rect 12492 4768 12498 4780
rect 12897 4777 12909 4780
rect 12943 4777 12955 4811
rect 13814 4808 13820 4820
rect 13775 4780 13820 4808
rect 12897 4771 12955 4777
rect 13814 4768 13820 4780
rect 13872 4768 13878 4820
rect 15289 4811 15347 4817
rect 15289 4777 15301 4811
rect 15335 4808 15347 4811
rect 15746 4808 15752 4820
rect 15335 4780 15752 4808
rect 15335 4777 15347 4780
rect 15289 4771 15347 4777
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 16117 4811 16175 4817
rect 16117 4777 16129 4811
rect 16163 4808 16175 4811
rect 16574 4808 16580 4820
rect 16163 4780 16580 4808
rect 16163 4777 16175 4780
rect 16117 4771 16175 4777
rect 16574 4768 16580 4780
rect 16632 4768 16638 4820
rect 17954 4808 17960 4820
rect 17328 4780 17960 4808
rect 11606 4740 11612 4752
rect 5092 4712 10548 4740
rect 1756 4675 1814 4681
rect 1756 4641 1768 4675
rect 1802 4672 1814 4675
rect 2958 4672 2964 4684
rect 1802 4644 2964 4672
rect 1802 4641 1814 4644
rect 1756 4635 1814 4641
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 3418 4672 3424 4684
rect 3379 4644 3424 4672
rect 3418 4632 3424 4644
rect 3476 4632 3482 4684
rect 5092 4681 5120 4712
rect 10520 4684 10548 4712
rect 10704 4712 11612 4740
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4641 4491 4675
rect 4433 4635 4491 4641
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4641 5135 4675
rect 5077 4635 5135 4641
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4573 1547 4607
rect 1489 4567 1547 4573
rect 1504 4468 1532 4567
rect 2866 4564 2872 4616
rect 2924 4604 2930 4616
rect 3970 4604 3976 4616
rect 2924 4576 3976 4604
rect 2924 4564 2930 4576
rect 3970 4564 3976 4576
rect 4028 4604 4034 4616
rect 4448 4604 4476 4635
rect 5718 4632 5724 4684
rect 5776 4672 5782 4684
rect 5885 4675 5943 4681
rect 5885 4672 5897 4675
rect 5776 4644 5897 4672
rect 5776 4632 5782 4644
rect 5885 4641 5897 4644
rect 5931 4672 5943 4675
rect 8757 4675 8815 4681
rect 5931 4644 7880 4672
rect 5931 4641 5943 4644
rect 5885 4635 5943 4641
rect 4614 4604 4620 4616
rect 4028 4576 4476 4604
rect 4575 4576 4620 4604
rect 4028 4564 4034 4576
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 7852 4613 7880 4644
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 9674 4672 9680 4684
rect 8803 4644 9680 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 9861 4675 9919 4681
rect 9861 4641 9873 4675
rect 9907 4641 9919 4675
rect 9861 4635 9919 4641
rect 5629 4607 5687 4613
rect 5629 4604 5641 4607
rect 5092 4576 5641 4604
rect 1854 4468 1860 4480
rect 1504 4440 1860 4468
rect 1854 4428 1860 4440
rect 1912 4468 1918 4480
rect 5092 4468 5120 4576
rect 5629 4573 5641 4576
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 8849 4607 8907 4613
rect 8849 4604 8861 4607
rect 8444 4576 8861 4604
rect 8444 4564 8450 4576
rect 8849 4573 8861 4576
rect 8895 4573 8907 4607
rect 9876 4604 9904 4635
rect 10502 4632 10508 4684
rect 10560 4632 10566 4684
rect 10704 4604 10732 4712
rect 11606 4700 11612 4712
rect 11664 4700 11670 4752
rect 12253 4743 12311 4749
rect 12253 4709 12265 4743
rect 12299 4740 12311 4743
rect 17328 4740 17356 4780
rect 17954 4768 17960 4780
rect 18012 4768 18018 4820
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 19794 4808 19800 4820
rect 19392 4780 19800 4808
rect 19392 4768 19398 4780
rect 19794 4768 19800 4780
rect 19852 4768 19858 4820
rect 12299 4712 17356 4740
rect 17396 4743 17454 4749
rect 12299 4709 12311 4712
rect 12253 4703 12311 4709
rect 17396 4709 17408 4743
rect 17442 4740 17454 4743
rect 17678 4740 17684 4752
rect 17442 4712 17684 4740
rect 17442 4709 17454 4712
rect 17396 4703 17454 4709
rect 17678 4700 17684 4712
rect 17736 4700 17742 4752
rect 18506 4700 18512 4752
rect 18564 4740 18570 4752
rect 21174 4740 21180 4752
rect 18564 4712 21180 4740
rect 18564 4700 18570 4712
rect 21174 4700 21180 4712
rect 21232 4700 21238 4752
rect 10781 4675 10839 4681
rect 10781 4641 10793 4675
rect 10827 4672 10839 4675
rect 10870 4672 10876 4684
rect 10827 4644 10876 4672
rect 10827 4641 10839 4644
rect 10781 4635 10839 4641
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 11514 4672 11520 4684
rect 10980 4644 11520 4672
rect 9876 4576 10732 4604
rect 8849 4567 8907 4573
rect 6638 4496 6644 4548
rect 6696 4536 6702 4548
rect 9490 4536 9496 4548
rect 6696 4508 9496 4536
rect 6696 4496 6702 4508
rect 9490 4496 9496 4508
rect 9548 4536 9554 4548
rect 10980 4536 11008 4644
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 12158 4672 12164 4684
rect 11992 4644 12164 4672
rect 11057 4607 11115 4613
rect 11057 4573 11069 4607
rect 11103 4604 11115 4607
rect 11698 4604 11704 4616
rect 11103 4576 11704 4604
rect 11103 4573 11115 4576
rect 11057 4567 11115 4573
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 11992 4613 12020 4644
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 12805 4675 12863 4681
rect 12805 4641 12817 4675
rect 12851 4672 12863 4675
rect 13630 4672 13636 4684
rect 12851 4644 13636 4672
rect 12851 4641 12863 4644
rect 12805 4635 12863 4641
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 13909 4675 13967 4681
rect 13909 4641 13921 4675
rect 13955 4672 13967 4675
rect 14550 4672 14556 4684
rect 13955 4644 14556 4672
rect 13955 4641 13967 4644
rect 13909 4635 13967 4641
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 14642 4632 14648 4684
rect 14700 4672 14706 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 14700 4644 15669 4672
rect 14700 4632 14706 4644
rect 15657 4641 15669 4644
rect 15703 4672 15715 4675
rect 16117 4675 16175 4681
rect 16117 4672 16129 4675
rect 15703 4644 16129 4672
rect 15703 4641 15715 4644
rect 15657 4635 15715 4641
rect 16117 4641 16129 4644
rect 16163 4641 16175 4675
rect 16117 4635 16175 4641
rect 16301 4675 16359 4681
rect 16301 4641 16313 4675
rect 16347 4641 16359 4675
rect 16301 4635 16359 4641
rect 11885 4607 11943 4613
rect 11885 4573 11897 4607
rect 11931 4573 11943 4607
rect 11885 4567 11943 4573
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 11900 4536 11928 4567
rect 12066 4564 12072 4616
rect 12124 4604 12130 4616
rect 12989 4607 13047 4613
rect 12989 4604 13001 4607
rect 12124 4576 13001 4604
rect 12124 4564 12130 4576
rect 12989 4573 13001 4576
rect 13035 4604 13047 4607
rect 14001 4607 14059 4613
rect 14001 4604 14013 4607
rect 13035 4576 14013 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 14001 4573 14013 4576
rect 14047 4604 14059 4607
rect 14366 4604 14372 4616
rect 14047 4576 14372 4604
rect 14047 4573 14059 4576
rect 14001 4567 14059 4573
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 15378 4604 15384 4616
rect 14476 4576 15384 4604
rect 13449 4539 13507 4545
rect 13449 4536 13461 4539
rect 9548 4508 11008 4536
rect 11072 4508 11744 4536
rect 11900 4508 13461 4536
rect 9548 4496 9554 4508
rect 1912 4440 5120 4468
rect 5261 4471 5319 4477
rect 1912 4428 1918 4440
rect 5261 4437 5273 4471
rect 5307 4468 5319 4471
rect 9858 4468 9864 4480
rect 5307 4440 9864 4468
rect 5307 4437 5319 4440
rect 5261 4431 5319 4437
rect 9858 4428 9864 4440
rect 9916 4428 9922 4480
rect 10042 4468 10048 4480
rect 10003 4440 10048 4468
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 10229 4471 10287 4477
rect 10229 4437 10241 4471
rect 10275 4468 10287 4471
rect 11072 4468 11100 4508
rect 10275 4440 11100 4468
rect 11425 4471 11483 4477
rect 10275 4437 10287 4440
rect 10229 4431 10287 4437
rect 11425 4437 11437 4471
rect 11471 4468 11483 4471
rect 11606 4468 11612 4480
rect 11471 4440 11612 4468
rect 11471 4437 11483 4440
rect 11425 4431 11483 4437
rect 11606 4428 11612 4440
rect 11664 4428 11670 4480
rect 11716 4468 11744 4508
rect 13449 4505 13461 4508
rect 13495 4505 13507 4539
rect 13449 4499 13507 4505
rect 12253 4471 12311 4477
rect 12253 4468 12265 4471
rect 11716 4440 12265 4468
rect 12253 4437 12265 4440
rect 12299 4437 12311 4471
rect 12253 4431 12311 4437
rect 12437 4471 12495 4477
rect 12437 4437 12449 4471
rect 12483 4468 12495 4471
rect 12894 4468 12900 4480
rect 12483 4440 12900 4468
rect 12483 4437 12495 4440
rect 12437 4431 12495 4437
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 13262 4428 13268 4480
rect 13320 4468 13326 4480
rect 14476 4468 14504 4576
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 15562 4564 15568 4616
rect 15620 4604 15626 4616
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15620 4576 15761 4604
rect 15620 4564 15626 4576
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4604 15991 4607
rect 16022 4604 16028 4616
rect 15979 4576 16028 4604
rect 15979 4573 15991 4576
rect 15933 4567 15991 4573
rect 16022 4564 16028 4576
rect 16080 4564 16086 4616
rect 15194 4496 15200 4548
rect 15252 4536 15258 4548
rect 16316 4536 16344 4635
rect 16390 4632 16396 4684
rect 16448 4672 16454 4684
rect 17126 4672 17132 4684
rect 16448 4644 17132 4672
rect 16448 4632 16454 4644
rect 17126 4632 17132 4644
rect 17184 4632 17190 4684
rect 19426 4672 19432 4684
rect 19387 4644 19432 4672
rect 19426 4632 19432 4644
rect 19484 4632 19490 4684
rect 19978 4632 19984 4684
rect 20036 4672 20042 4684
rect 20073 4675 20131 4681
rect 20073 4672 20085 4675
rect 20036 4644 20085 4672
rect 20036 4632 20042 4644
rect 20073 4641 20085 4644
rect 20119 4672 20131 4675
rect 20806 4672 20812 4684
rect 20119 4644 20812 4672
rect 20119 4641 20131 4644
rect 20073 4635 20131 4641
rect 20806 4632 20812 4644
rect 20864 4632 20870 4684
rect 16574 4604 16580 4616
rect 16535 4576 16580 4604
rect 16574 4564 16580 4576
rect 16632 4564 16638 4616
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19521 4607 19579 4613
rect 19521 4604 19533 4607
rect 19392 4576 19533 4604
rect 19392 4564 19398 4576
rect 19521 4573 19533 4576
rect 19567 4573 19579 4607
rect 19521 4567 19579 4573
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4604 19763 4607
rect 19886 4604 19892 4616
rect 19751 4576 19892 4604
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 19886 4564 19892 4576
rect 19944 4564 19950 4616
rect 20346 4604 20352 4616
rect 20307 4576 20352 4604
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 20530 4564 20536 4616
rect 20588 4604 20594 4616
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 20588 4576 20913 4604
rect 20588 4564 20594 4576
rect 20901 4573 20913 4576
rect 20947 4573 20959 4607
rect 20901 4567 20959 4573
rect 15252 4508 16344 4536
rect 15252 4496 15258 4508
rect 13320 4440 14504 4468
rect 14829 4471 14887 4477
rect 13320 4428 13326 4440
rect 14829 4437 14841 4471
rect 14875 4468 14887 4471
rect 16206 4468 16212 4480
rect 14875 4440 16212 4468
rect 14875 4437 14887 4440
rect 14829 4431 14887 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 18509 4471 18567 4477
rect 18509 4437 18521 4471
rect 18555 4468 18567 4471
rect 18966 4468 18972 4480
rect 18555 4440 18972 4468
rect 18555 4437 18567 4440
rect 18509 4431 18567 4437
rect 18966 4428 18972 4440
rect 19024 4428 19030 4480
rect 19061 4471 19119 4477
rect 19061 4437 19073 4471
rect 19107 4468 19119 4471
rect 20070 4468 20076 4480
rect 19107 4440 20076 4468
rect 19107 4437 19119 4440
rect 19061 4431 19119 4437
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 3418 4224 3424 4276
rect 3476 4224 3482 4276
rect 3697 4267 3755 4273
rect 3697 4233 3709 4267
rect 3743 4264 3755 4267
rect 4706 4264 4712 4276
rect 3743 4236 4712 4264
rect 3743 4233 3755 4236
rect 3697 4227 3755 4233
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 6089 4267 6147 4273
rect 6089 4233 6101 4267
rect 6135 4264 6147 4267
rect 7098 4264 7104 4276
rect 6135 4236 7104 4264
rect 6135 4233 6147 4236
rect 6089 4227 6147 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 7558 4224 7564 4276
rect 7616 4264 7622 4276
rect 8202 4264 8208 4276
rect 7616 4236 8208 4264
rect 7616 4224 7622 4236
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 10042 4224 10048 4276
rect 10100 4264 10106 4276
rect 13262 4264 13268 4276
rect 10100 4236 13268 4264
rect 10100 4224 10106 4236
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 13354 4224 13360 4276
rect 13412 4264 13418 4276
rect 13412 4236 14044 4264
rect 13412 4224 13418 4236
rect 3436 4196 3464 4224
rect 6822 4196 6828 4208
rect 3436 4168 6828 4196
rect 6822 4156 6828 4168
rect 6880 4156 6886 4208
rect 10962 4196 10968 4208
rect 10336 4168 10968 4196
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 2958 4128 2964 4140
rect 2547 4100 2964 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 3418 4128 3424 4140
rect 3379 4100 3424 4128
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 4430 4128 4436 4140
rect 4264 4100 4436 4128
rect 4264 4069 4292 4100
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4128 4583 4131
rect 5074 4128 5080 4140
rect 4571 4100 5080 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 5074 4088 5080 4100
rect 5132 4128 5138 4140
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 5132 4100 5457 4128
rect 5132 4088 5138 4100
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 5445 4091 5503 4097
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7285 4131 7343 4137
rect 7285 4128 7297 4131
rect 6972 4100 7297 4128
rect 6972 4088 6978 4100
rect 7285 4097 7297 4100
rect 7331 4097 7343 4131
rect 7285 4091 7343 4097
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4128 7527 4131
rect 8110 4128 8116 4140
rect 7515 4100 8116 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8570 4128 8576 4140
rect 8531 4100 8576 4128
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 10336 4128 10364 4168
rect 10962 4156 10968 4168
rect 11020 4156 11026 4208
rect 14016 4196 14044 4236
rect 14366 4224 14372 4276
rect 14424 4264 14430 4276
rect 14461 4267 14519 4273
rect 14461 4264 14473 4267
rect 14424 4236 14473 4264
rect 14424 4224 14430 4236
rect 14461 4233 14473 4236
rect 14507 4233 14519 4267
rect 14461 4227 14519 4233
rect 14550 4224 14556 4276
rect 14608 4264 14614 4276
rect 14737 4267 14795 4273
rect 14737 4264 14749 4267
rect 14608 4236 14749 4264
rect 14608 4224 14614 4236
rect 14737 4233 14749 4236
rect 14783 4233 14795 4267
rect 14737 4227 14795 4233
rect 14918 4224 14924 4276
rect 14976 4264 14982 4276
rect 14976 4236 15424 4264
rect 14976 4224 14982 4236
rect 14182 4196 14188 4208
rect 11440 4168 11744 4196
rect 14016 4168 14188 4196
rect 11440 4128 11468 4168
rect 11606 4128 11612 4140
rect 9640 4100 10364 4128
rect 10428 4100 11468 4128
rect 11567 4100 11612 4128
rect 9640 4088 9646 4100
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 3697 4063 3755 4069
rect 3697 4060 3709 4063
rect 1443 4032 3709 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 3697 4029 3709 4032
rect 3743 4029 3755 4063
rect 3697 4023 3755 4029
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 4706 4020 4712 4072
rect 4764 4060 4770 4072
rect 5258 4060 5264 4072
rect 4764 4032 5120 4060
rect 5219 4032 5264 4060
rect 4764 4020 4770 4032
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3992 2283 3995
rect 3142 3992 3148 4004
rect 2271 3964 3148 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 3142 3952 3148 3964
rect 3200 3952 3206 4004
rect 3237 3995 3295 4001
rect 3237 3961 3249 3995
rect 3283 3992 3295 3995
rect 5092 3992 5120 4032
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 5353 4063 5411 4069
rect 5353 4029 5365 4063
rect 5399 4060 5411 4063
rect 6089 4063 6147 4069
rect 6089 4060 6101 4063
rect 5399 4032 6101 4060
rect 5399 4029 5411 4032
rect 5353 4023 5411 4029
rect 6089 4029 6101 4032
rect 6135 4029 6147 4063
rect 6089 4023 6147 4029
rect 6181 4063 6239 4069
rect 6181 4029 6193 4063
rect 6227 4060 6239 4063
rect 6270 4060 6276 4072
rect 6227 4032 6276 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 7190 4060 7196 4072
rect 7151 4032 7196 4060
rect 7190 4020 7196 4032
rect 7248 4020 7254 4072
rect 8018 4060 8024 4072
rect 7979 4032 8024 4060
rect 8018 4020 8024 4032
rect 8076 4020 8082 4072
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 8588 4032 10241 4060
rect 5166 3992 5172 4004
rect 3283 3964 4936 3992
rect 5092 3964 5172 3992
rect 3283 3961 3295 3964
rect 3237 3955 3295 3961
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 2869 3927 2927 3933
rect 2869 3924 2881 3927
rect 2363 3896 2881 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 2869 3893 2881 3896
rect 2915 3893 2927 3927
rect 3326 3924 3332 3936
rect 3287 3896 3332 3924
rect 2869 3887 2927 3893
rect 3326 3884 3332 3896
rect 3384 3884 3390 3936
rect 3881 3927 3939 3933
rect 3881 3893 3893 3927
rect 3927 3924 3939 3927
rect 4154 3924 4160 3936
rect 3927 3896 4160 3924
rect 3927 3893 3939 3896
rect 3881 3887 3939 3893
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 4246 3884 4252 3936
rect 4304 3924 4310 3936
rect 4908 3933 4936 3964
rect 5166 3952 5172 3964
rect 5224 3952 5230 4004
rect 8588 3992 8616 4032
rect 10229 4029 10241 4032
rect 10275 4029 10287 4063
rect 10229 4023 10287 4029
rect 6840 3964 8616 3992
rect 8840 3995 8898 4001
rect 4341 3927 4399 3933
rect 4341 3924 4353 3927
rect 4304 3896 4353 3924
rect 4304 3884 4310 3896
rect 4341 3893 4353 3896
rect 4387 3893 4399 3927
rect 4341 3887 4399 3893
rect 4893 3927 4951 3933
rect 4893 3893 4905 3927
rect 4939 3893 4951 3927
rect 6362 3924 6368 3936
rect 6323 3896 6368 3924
rect 4893 3887 4951 3893
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 6840 3933 6868 3964
rect 8840 3961 8852 3995
rect 8886 3992 8898 3995
rect 10428 3992 10456 4100
rect 11606 4088 11612 4100
rect 11664 4088 11670 4140
rect 11716 4137 11744 4168
rect 14182 4156 14188 4168
rect 14240 4196 14246 4208
rect 14240 4168 15332 4196
rect 14240 4156 14246 4168
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 12066 4128 12072 4140
rect 11747 4100 12072 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12618 4128 12624 4140
rect 12452 4100 12624 4128
rect 10502 4020 10508 4072
rect 10560 4060 10566 4072
rect 10560 4032 10605 4060
rect 10560 4020 10566 4032
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 12452 4060 12480 4100
rect 12618 4088 12624 4100
rect 12676 4128 12682 4140
rect 13081 4131 13139 4137
rect 13081 4128 13093 4131
rect 12676 4100 13093 4128
rect 12676 4088 12682 4100
rect 13081 4097 13093 4100
rect 13127 4097 13139 4131
rect 13081 4091 13139 4097
rect 15010 4088 15016 4140
rect 15068 4128 15074 4140
rect 15304 4137 15332 4168
rect 15197 4131 15255 4137
rect 15197 4128 15209 4131
rect 15068 4100 15209 4128
rect 15068 4088 15074 4100
rect 15197 4097 15209 4100
rect 15243 4097 15255 4131
rect 15197 4091 15255 4097
rect 15289 4131 15347 4137
rect 15289 4097 15301 4131
rect 15335 4097 15347 4131
rect 15396 4128 15424 4236
rect 15470 4224 15476 4276
rect 15528 4264 15534 4276
rect 16850 4264 16856 4276
rect 15528 4236 16856 4264
rect 15528 4224 15534 4236
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 19610 4264 19616 4276
rect 19168 4236 19616 4264
rect 16761 4199 16819 4205
rect 16761 4165 16773 4199
rect 16807 4196 16819 4199
rect 17034 4196 17040 4208
rect 16807 4168 17040 4196
rect 16807 4165 16819 4168
rect 16761 4159 16819 4165
rect 17034 4156 17040 4168
rect 17092 4156 17098 4208
rect 17126 4156 17132 4208
rect 17184 4196 17190 4208
rect 19168 4196 19196 4236
rect 19610 4224 19616 4236
rect 19668 4224 19674 4276
rect 19705 4267 19763 4273
rect 19705 4233 19717 4267
rect 19751 4264 19763 4267
rect 20438 4264 20444 4276
rect 19751 4236 20444 4264
rect 19751 4233 19763 4236
rect 19705 4227 19763 4233
rect 20438 4224 20444 4236
rect 20496 4224 20502 4276
rect 17184 4168 18092 4196
rect 17184 4156 17190 4168
rect 16390 4128 16396 4140
rect 15396 4100 16252 4128
rect 16351 4100 16396 4128
rect 15289 4091 15347 4097
rect 10836 4032 12480 4060
rect 10836 4020 10842 4032
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 16117 4063 16175 4069
rect 16117 4060 16129 4063
rect 12584 4032 12629 4060
rect 13188 4032 16129 4060
rect 12584 4020 12590 4032
rect 8886 3964 10456 3992
rect 8886 3961 8898 3964
rect 8840 3955 8898 3961
rect 10594 3952 10600 4004
rect 10652 3992 10658 4004
rect 11422 3992 11428 4004
rect 10652 3964 11428 3992
rect 10652 3952 10658 3964
rect 11422 3952 11428 3964
rect 11480 3952 11486 4004
rect 11517 3995 11575 4001
rect 11517 3961 11529 3995
rect 11563 3992 11575 3995
rect 12434 3992 12440 4004
rect 11563 3964 12440 3992
rect 11563 3961 11575 3964
rect 11517 3955 11575 3961
rect 12434 3952 12440 3964
rect 12492 3952 12498 4004
rect 13188 3992 13216 4032
rect 16117 4029 16129 4032
rect 16163 4029 16175 4063
rect 16224 4060 16252 4100
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 17405 4131 17463 4137
rect 17405 4097 17417 4131
rect 17451 4097 17463 4131
rect 17405 4091 17463 4097
rect 16224 4032 17356 4060
rect 16117 4023 16175 4029
rect 13354 4001 13360 4004
rect 13348 3992 13360 4001
rect 12544 3964 13216 3992
rect 13315 3964 13360 3992
rect 12544 3936 12572 3964
rect 13348 3955 13360 3964
rect 13354 3952 13360 3955
rect 13412 3952 13418 4004
rect 13814 3952 13820 4004
rect 13872 3992 13878 4004
rect 14918 3992 14924 4004
rect 13872 3964 14924 3992
rect 13872 3952 13878 3964
rect 14918 3952 14924 3964
rect 14976 3952 14982 4004
rect 15010 3952 15016 4004
rect 15068 3992 15074 4004
rect 17221 3995 17279 4001
rect 17221 3992 17233 3995
rect 15068 3964 17233 3992
rect 15068 3952 15074 3964
rect 17221 3961 17233 3964
rect 17267 3961 17279 3995
rect 17221 3955 17279 3961
rect 6825 3927 6883 3933
rect 6825 3893 6837 3927
rect 6871 3893 6883 3927
rect 6825 3887 6883 3893
rect 8205 3927 8263 3933
rect 8205 3893 8217 3927
rect 8251 3924 8263 3927
rect 9214 3924 9220 3936
rect 8251 3896 9220 3924
rect 8251 3893 8263 3896
rect 8205 3887 8263 3893
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 9953 3927 10011 3933
rect 9953 3893 9965 3927
rect 9999 3924 10011 3927
rect 10226 3924 10232 3936
rect 9999 3896 10232 3924
rect 9999 3893 10011 3896
rect 9953 3887 10011 3893
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 11149 3927 11207 3933
rect 11149 3893 11161 3927
rect 11195 3924 11207 3927
rect 11790 3924 11796 3936
rect 11195 3896 11796 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12526 3884 12532 3936
rect 12584 3884 12590 3936
rect 12713 3927 12771 3933
rect 12713 3893 12725 3927
rect 12759 3924 12771 3927
rect 12986 3924 12992 3936
rect 12759 3896 12992 3924
rect 12759 3893 12771 3896
rect 12713 3887 12771 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 14458 3924 14464 3936
rect 13136 3896 14464 3924
rect 13136 3884 13142 3896
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 15105 3927 15163 3933
rect 15105 3893 15117 3927
rect 15151 3924 15163 3927
rect 15470 3924 15476 3936
rect 15151 3896 15476 3924
rect 15151 3893 15163 3896
rect 15105 3887 15163 3893
rect 15470 3884 15476 3896
rect 15528 3884 15534 3936
rect 15746 3924 15752 3936
rect 15707 3896 15752 3924
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 15838 3884 15844 3936
rect 15896 3924 15902 3936
rect 16209 3927 16267 3933
rect 16209 3924 16221 3927
rect 15896 3896 16221 3924
rect 15896 3884 15902 3896
rect 16209 3893 16221 3896
rect 16255 3893 16267 3927
rect 17126 3924 17132 3936
rect 17087 3896 17132 3924
rect 16209 3887 16267 3893
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 17328 3924 17356 4032
rect 17420 4004 17448 4091
rect 17678 4088 17684 4140
rect 17736 4128 17742 4140
rect 18064 4137 18092 4168
rect 19076 4168 19196 4196
rect 18049 4131 18107 4137
rect 17736 4100 18000 4128
rect 17736 4088 17742 4100
rect 17972 4060 18000 4100
rect 18049 4097 18061 4131
rect 18095 4097 18107 4131
rect 18049 4091 18107 4097
rect 19076 4060 19104 4168
rect 20162 4156 20168 4208
rect 20220 4196 20226 4208
rect 20220 4168 20300 4196
rect 20220 4156 20226 4168
rect 20272 4137 20300 4168
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 17972 4032 19104 4060
rect 19150 4020 19156 4072
rect 19208 4060 19214 4072
rect 19518 4060 19524 4072
rect 19208 4032 19524 4060
rect 19208 4020 19214 4032
rect 19518 4020 19524 4032
rect 19576 4020 19582 4072
rect 20070 4060 20076 4072
rect 20031 4032 20076 4060
rect 20070 4020 20076 4032
rect 20128 4020 20134 4072
rect 20717 4063 20775 4069
rect 20717 4029 20729 4063
rect 20763 4060 20775 4063
rect 20806 4060 20812 4072
rect 20763 4032 20812 4060
rect 20763 4029 20775 4032
rect 20717 4023 20775 4029
rect 20806 4020 20812 4032
rect 20864 4020 20870 4072
rect 17402 3952 17408 4004
rect 17460 3992 17466 4004
rect 18316 3995 18374 4001
rect 18316 3992 18328 3995
rect 17460 3964 17908 3992
rect 17460 3952 17466 3964
rect 17678 3924 17684 3936
rect 17328 3896 17684 3924
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 17880 3924 17908 3964
rect 18064 3964 18328 3992
rect 18064 3924 18092 3964
rect 18316 3961 18328 3964
rect 18362 3992 18374 3995
rect 18690 3992 18696 4004
rect 18362 3964 18696 3992
rect 18362 3961 18374 3964
rect 18316 3955 18374 3961
rect 18690 3952 18696 3964
rect 18748 3952 18754 4004
rect 19702 3952 19708 4004
rect 19760 3992 19766 4004
rect 20165 3995 20223 4001
rect 20165 3992 20177 3995
rect 19760 3964 20177 3992
rect 19760 3952 19766 3964
rect 20165 3961 20177 3964
rect 20211 3961 20223 3995
rect 20165 3955 20223 3961
rect 17880 3896 18092 3924
rect 19429 3927 19487 3933
rect 19429 3893 19441 3927
rect 19475 3924 19487 3927
rect 19886 3924 19892 3936
rect 19475 3896 19892 3924
rect 19475 3893 19487 3896
rect 19429 3887 19487 3893
rect 19886 3884 19892 3896
rect 19944 3884 19950 3936
rect 20438 3884 20444 3936
rect 20496 3924 20502 3936
rect 20901 3927 20959 3933
rect 20901 3924 20913 3927
rect 20496 3896 20913 3924
rect 20496 3884 20502 3896
rect 20901 3893 20913 3896
rect 20947 3893 20959 3927
rect 20901 3887 20959 3893
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 934 3680 940 3732
rect 992 3720 998 3732
rect 2866 3720 2872 3732
rect 992 3692 2872 3720
rect 992 3680 998 3692
rect 2866 3680 2872 3692
rect 2924 3680 2930 3732
rect 3326 3680 3332 3732
rect 3384 3720 3390 3732
rect 4157 3723 4215 3729
rect 4157 3720 4169 3723
rect 3384 3692 4169 3720
rect 3384 3680 3390 3692
rect 4157 3689 4169 3692
rect 4203 3689 4215 3723
rect 4157 3683 4215 3689
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 4304 3692 4349 3720
rect 4304 3680 4310 3692
rect 4706 3680 4712 3732
rect 4764 3720 4770 3732
rect 4801 3723 4859 3729
rect 4801 3720 4813 3723
rect 4764 3692 4813 3720
rect 4764 3680 4770 3692
rect 4801 3689 4813 3692
rect 4847 3689 4859 3723
rect 4801 3683 4859 3689
rect 5813 3723 5871 3729
rect 5813 3689 5825 3723
rect 5859 3720 5871 3723
rect 8294 3720 8300 3732
rect 5859 3692 8300 3720
rect 5859 3689 5871 3692
rect 5813 3683 5871 3689
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 9122 3720 9128 3732
rect 8404 3692 9128 3720
rect 5905 3655 5963 3661
rect 5905 3652 5917 3655
rect 4724 3624 5917 3652
rect 2216 3587 2274 3593
rect 2216 3553 2228 3587
rect 2262 3584 2274 3587
rect 3326 3584 3332 3596
rect 2262 3556 3332 3584
rect 2262 3553 2274 3556
rect 2216 3547 2274 3553
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4724 3584 4752 3624
rect 5905 3621 5917 3624
rect 5951 3621 5963 3655
rect 7742 3652 7748 3664
rect 5905 3615 5963 3621
rect 7116 3624 7748 3652
rect 5353 3587 5411 3593
rect 5353 3584 5365 3587
rect 4212 3556 4752 3584
rect 4908 3556 5365 3584
rect 4212 3544 4218 3556
rect 1486 3516 1492 3528
rect 1447 3488 1492 3516
rect 1486 3476 1492 3488
rect 1544 3476 1550 3528
rect 1946 3516 1952 3528
rect 1907 3488 1952 3516
rect 1946 3476 1952 3488
rect 2004 3476 2010 3528
rect 3142 3476 3148 3528
rect 3200 3516 3206 3528
rect 3200 3488 3464 3516
rect 3200 3476 3206 3488
rect 3329 3451 3387 3457
rect 3329 3448 3341 3451
rect 3068 3420 3341 3448
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 3068 3380 3096 3420
rect 3329 3417 3341 3420
rect 3375 3417 3387 3451
rect 3436 3448 3464 3488
rect 4246 3476 4252 3528
rect 4304 3516 4310 3528
rect 4908 3525 4936 3556
rect 5353 3553 5365 3556
rect 5399 3584 5411 3587
rect 5534 3584 5540 3596
rect 5399 3556 5540 3584
rect 5399 3553 5411 3556
rect 5353 3547 5411 3553
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 7009 3587 7067 3593
rect 7009 3584 7021 3587
rect 6972 3556 7021 3584
rect 6972 3544 6978 3556
rect 7009 3553 7021 3556
rect 7055 3553 7067 3587
rect 7009 3547 7067 3553
rect 7116 3528 7144 3624
rect 7742 3612 7748 3624
rect 7800 3612 7806 3664
rect 8110 3652 8116 3664
rect 8071 3624 8116 3652
rect 8110 3612 8116 3624
rect 8168 3612 8174 3664
rect 7558 3544 7564 3596
rect 7616 3584 7622 3596
rect 8021 3587 8079 3593
rect 8021 3584 8033 3587
rect 7616 3556 8033 3584
rect 7616 3544 7622 3556
rect 8021 3553 8033 3556
rect 8067 3584 8079 3587
rect 8404 3584 8432 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9674 3720 9680 3732
rect 9635 3692 9680 3720
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 10045 3723 10103 3729
rect 10045 3689 10057 3723
rect 10091 3720 10103 3723
rect 10318 3720 10324 3732
rect 10091 3692 10324 3720
rect 10091 3689 10103 3692
rect 10045 3683 10103 3689
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 11330 3720 11336 3732
rect 10928 3692 11336 3720
rect 10928 3680 10934 3692
rect 11330 3680 11336 3692
rect 11388 3680 11394 3732
rect 11514 3680 11520 3732
rect 11572 3720 11578 3732
rect 12253 3723 12311 3729
rect 12253 3720 12265 3723
rect 11572 3692 12265 3720
rect 11572 3680 11578 3692
rect 12253 3689 12265 3692
rect 12299 3689 12311 3723
rect 12434 3720 12440 3732
rect 12395 3692 12440 3720
rect 12253 3683 12311 3689
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 12805 3723 12863 3729
rect 12805 3689 12817 3723
rect 12851 3720 12863 3723
rect 13449 3723 13507 3729
rect 13449 3720 13461 3723
rect 12851 3692 13461 3720
rect 12851 3689 12863 3692
rect 12805 3683 12863 3689
rect 13449 3689 13461 3692
rect 13495 3689 13507 3723
rect 13906 3720 13912 3732
rect 13867 3692 13912 3720
rect 13449 3683 13507 3689
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 15746 3680 15752 3732
rect 15804 3720 15810 3732
rect 15804 3692 17724 3720
rect 15804 3680 15810 3692
rect 9214 3612 9220 3664
rect 9272 3652 9278 3664
rect 12894 3652 12900 3664
rect 9272 3624 12020 3652
rect 12855 3624 12900 3652
rect 9272 3612 9278 3624
rect 8067 3556 8432 3584
rect 8067 3553 8079 3556
rect 8021 3547 8079 3553
rect 8662 3544 8668 3596
rect 8720 3584 8726 3596
rect 8849 3587 8907 3593
rect 8849 3584 8861 3587
rect 8720 3556 8861 3584
rect 8720 3544 8726 3556
rect 8849 3553 8861 3556
rect 8895 3553 8907 3587
rect 8849 3547 8907 3553
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3584 9183 3587
rect 9398 3584 9404 3596
rect 9171 3556 9404 3584
rect 9171 3553 9183 3556
rect 9125 3547 9183 3553
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 11048 3587 11106 3593
rect 11048 3553 11060 3587
rect 11094 3584 11106 3587
rect 11882 3584 11888 3596
rect 11094 3556 11888 3584
rect 11094 3553 11106 3556
rect 11048 3547 11106 3553
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 11992 3584 12020 3624
rect 12894 3612 12900 3624
rect 12952 3612 12958 3664
rect 13538 3612 13544 3664
rect 13596 3652 13602 3664
rect 16574 3652 16580 3664
rect 13596 3624 14596 3652
rect 13596 3612 13602 3624
rect 13630 3584 13636 3596
rect 11992 3556 13636 3584
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 13817 3587 13875 3593
rect 13817 3553 13829 3587
rect 13863 3553 13875 3587
rect 14458 3584 14464 3596
rect 14419 3556 14464 3584
rect 13817 3547 13875 3553
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4304 3488 4905 3516
rect 4304 3476 4310 3488
rect 4893 3485 4905 3488
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3516 5135 3519
rect 5166 3516 5172 3528
rect 5123 3488 5172 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 5316 3488 6009 3516
rect 5316 3476 5322 3488
rect 5997 3485 6009 3488
rect 6043 3485 6055 3519
rect 7098 3516 7104 3528
rect 7059 3488 7104 3516
rect 5997 3479 6055 3485
rect 7098 3476 7104 3488
rect 7156 3476 7162 3528
rect 7190 3476 7196 3528
rect 7248 3516 7254 3528
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 7248 3488 7297 3516
rect 7248 3476 7254 3488
rect 7285 3485 7297 3488
rect 7331 3516 7343 3519
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 7331 3488 8309 3516
rect 7331 3485 7343 3488
rect 7285 3479 7343 3485
rect 8297 3485 8309 3488
rect 8343 3516 8355 3519
rect 8386 3516 8392 3528
rect 8343 3488 8392 3516
rect 8343 3485 8355 3488
rect 8297 3479 8355 3485
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 10134 3516 10140 3528
rect 10095 3488 10140 3516
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 10226 3476 10232 3528
rect 10284 3516 10290 3528
rect 10778 3516 10784 3528
rect 10284 3488 10329 3516
rect 10739 3488 10784 3516
rect 10284 3476 10290 3488
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 12158 3476 12164 3528
rect 12216 3516 12222 3528
rect 12989 3519 13047 3525
rect 12216 3488 12756 3516
rect 12216 3476 12222 3488
rect 5445 3451 5503 3457
rect 5445 3448 5457 3451
rect 3436 3420 5457 3448
rect 3329 3411 3387 3417
rect 5445 3417 5457 3420
rect 5491 3417 5503 3451
rect 5445 3411 5503 3417
rect 6362 3408 6368 3460
rect 6420 3448 6426 3460
rect 12618 3448 12624 3460
rect 6420 3420 10824 3448
rect 6420 3408 6426 3420
rect 3016 3352 3096 3380
rect 4157 3383 4215 3389
rect 3016 3340 3022 3352
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 4433 3383 4491 3389
rect 4433 3380 4445 3383
rect 4203 3352 4445 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 4433 3349 4445 3352
rect 4479 3349 4491 3383
rect 4433 3343 4491 3349
rect 6270 3340 6276 3392
rect 6328 3380 6334 3392
rect 6641 3383 6699 3389
rect 6641 3380 6653 3383
rect 6328 3352 6653 3380
rect 6328 3340 6334 3352
rect 6641 3349 6653 3352
rect 6687 3349 6699 3383
rect 7650 3380 7656 3392
rect 7611 3352 7656 3380
rect 6641 3343 6699 3349
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 8202 3340 8208 3392
rect 8260 3380 8266 3392
rect 8846 3380 8852 3392
rect 8260 3352 8852 3380
rect 8260 3340 8266 3352
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 8938 3340 8944 3392
rect 8996 3380 9002 3392
rect 10410 3380 10416 3392
rect 8996 3352 10416 3380
rect 8996 3340 9002 3352
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 10796 3380 10824 3420
rect 11716 3420 12624 3448
rect 11716 3380 11744 3420
rect 12618 3408 12624 3420
rect 12676 3408 12682 3460
rect 12728 3448 12756 3488
rect 12989 3485 13001 3519
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 13004 3448 13032 3479
rect 12728 3420 13032 3448
rect 13832 3448 13860 3547
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 14568 3584 14596 3624
rect 15304 3624 16580 3652
rect 15304 3593 15332 3624
rect 16574 3612 16580 3624
rect 16632 3612 16638 3664
rect 17696 3652 17724 3692
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 18417 3723 18475 3729
rect 18417 3720 18429 3723
rect 18012 3692 18429 3720
rect 18012 3680 18018 3692
rect 18417 3689 18429 3692
rect 18463 3689 18475 3723
rect 18417 3683 18475 3689
rect 18509 3723 18567 3729
rect 18509 3689 18521 3723
rect 18555 3720 18567 3723
rect 18598 3720 18604 3732
rect 18555 3692 18604 3720
rect 18555 3689 18567 3692
rect 18509 3683 18567 3689
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 19153 3723 19211 3729
rect 19153 3689 19165 3723
rect 19199 3720 19211 3723
rect 19334 3720 19340 3732
rect 19199 3692 19340 3720
rect 19199 3689 19211 3692
rect 19153 3683 19211 3689
rect 19334 3680 19340 3692
rect 19392 3680 19398 3732
rect 19518 3720 19524 3732
rect 19479 3692 19524 3720
rect 19518 3680 19524 3692
rect 19576 3680 19582 3732
rect 19794 3680 19800 3732
rect 19852 3720 19858 3732
rect 20162 3720 20168 3732
rect 19852 3692 20168 3720
rect 19852 3680 19858 3692
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 19613 3655 19671 3661
rect 19613 3652 19625 3655
rect 17696 3624 19625 3652
rect 19613 3621 19625 3624
rect 19659 3621 19671 3655
rect 19613 3615 19671 3621
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14568 3556 14749 3584
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 15841 3587 15899 3593
rect 15841 3553 15853 3587
rect 15887 3584 15899 3587
rect 15930 3584 15936 3596
rect 15887 3556 15936 3584
rect 15887 3553 15899 3556
rect 15841 3547 15899 3553
rect 15930 3544 15936 3556
rect 15988 3544 15994 3596
rect 16108 3587 16166 3593
rect 16108 3553 16120 3587
rect 16154 3584 16166 3587
rect 16390 3584 16396 3596
rect 16154 3556 16396 3584
rect 16154 3553 16166 3556
rect 16108 3547 16166 3553
rect 16390 3544 16396 3556
rect 16448 3544 16454 3596
rect 17310 3544 17316 3596
rect 17368 3584 17374 3596
rect 17497 3587 17555 3593
rect 17497 3584 17509 3587
rect 17368 3556 17509 3584
rect 17368 3544 17374 3556
rect 17497 3553 17509 3556
rect 17543 3553 17555 3587
rect 20165 3587 20223 3593
rect 20165 3584 20177 3587
rect 17497 3547 17555 3553
rect 17604 3556 20177 3584
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3516 14151 3519
rect 14366 3516 14372 3528
rect 14139 3488 14372 3516
rect 14139 3485 14151 3488
rect 14093 3479 14151 3485
rect 14366 3476 14372 3488
rect 14424 3476 14430 3528
rect 16850 3476 16856 3528
rect 16908 3516 16914 3528
rect 17604 3516 17632 3556
rect 20165 3553 20177 3556
rect 20211 3553 20223 3587
rect 20165 3547 20223 3553
rect 18690 3516 18696 3528
rect 16908 3488 17632 3516
rect 18603 3488 18696 3516
rect 16908 3476 16914 3488
rect 18690 3476 18696 3488
rect 18748 3516 18754 3528
rect 19794 3516 19800 3528
rect 18748 3488 19800 3516
rect 18748 3476 18754 3488
rect 19794 3476 19800 3488
rect 19852 3476 19858 3528
rect 20901 3519 20959 3525
rect 20901 3485 20913 3519
rect 20947 3485 20959 3519
rect 20901 3479 20959 3485
rect 20916 3448 20944 3479
rect 13832 3420 15884 3448
rect 12158 3380 12164 3392
rect 10796 3352 11744 3380
rect 12119 3352 12164 3380
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 12253 3383 12311 3389
rect 12253 3349 12265 3383
rect 12299 3380 12311 3383
rect 12894 3380 12900 3392
rect 12299 3352 12900 3380
rect 12299 3349 12311 3352
rect 12253 3343 12311 3349
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13262 3340 13268 3392
rect 13320 3380 13326 3392
rect 14550 3380 14556 3392
rect 13320 3352 14556 3380
rect 13320 3340 13326 3352
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 15470 3380 15476 3392
rect 15431 3352 15476 3380
rect 15470 3340 15476 3352
rect 15528 3340 15534 3392
rect 15856 3380 15884 3420
rect 16776 3420 20944 3448
rect 16776 3380 16804 3420
rect 15856 3352 16804 3380
rect 17221 3383 17279 3389
rect 17221 3349 17233 3383
rect 17267 3380 17279 3383
rect 17402 3380 17408 3392
rect 17267 3352 17408 3380
rect 17267 3349 17279 3352
rect 17221 3343 17279 3349
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 17681 3383 17739 3389
rect 17681 3349 17693 3383
rect 17727 3380 17739 3383
rect 17862 3380 17868 3392
rect 17727 3352 17868 3380
rect 17727 3349 17739 3352
rect 17681 3343 17739 3349
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 18049 3383 18107 3389
rect 18049 3349 18061 3383
rect 18095 3380 18107 3383
rect 19702 3380 19708 3392
rect 18095 3352 19708 3380
rect 18095 3349 18107 3352
rect 18049 3343 18107 3349
rect 19702 3340 19708 3352
rect 19760 3340 19766 3392
rect 20070 3340 20076 3392
rect 20128 3380 20134 3392
rect 20349 3383 20407 3389
rect 20349 3380 20361 3383
rect 20128 3352 20361 3380
rect 20128 3340 20134 3352
rect 20349 3349 20361 3352
rect 20395 3349 20407 3383
rect 20349 3343 20407 3349
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 1673 3179 1731 3185
rect 1673 3145 1685 3179
rect 1719 3176 1731 3179
rect 2498 3176 2504 3188
rect 1719 3148 2504 3176
rect 1719 3145 1731 3148
rect 1673 3139 1731 3145
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 2590 3136 2596 3188
rect 2648 3176 2654 3188
rect 2685 3179 2743 3185
rect 2685 3176 2697 3179
rect 2648 3148 2697 3176
rect 2648 3136 2654 3148
rect 2685 3145 2697 3148
rect 2731 3145 2743 3179
rect 2685 3139 2743 3145
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 5258 3176 5264 3188
rect 3384 3148 5264 3176
rect 3384 3136 3390 3148
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 5721 3179 5779 3185
rect 5721 3145 5733 3179
rect 5767 3176 5779 3179
rect 6178 3176 6184 3188
rect 5767 3148 6184 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 6380 3148 8217 3176
rect 6380 3052 6408 3148
rect 8205 3145 8217 3148
rect 8251 3145 8263 3179
rect 8205 3139 8263 3145
rect 8386 3136 8392 3188
rect 8444 3176 8450 3188
rect 8846 3176 8852 3188
rect 8444 3148 8852 3176
rect 8444 3136 8450 3148
rect 8846 3136 8852 3148
rect 8904 3176 8910 3188
rect 9861 3179 9919 3185
rect 9861 3176 9873 3179
rect 8904 3148 9873 3176
rect 8904 3136 8910 3148
rect 9861 3145 9873 3148
rect 9907 3145 9919 3179
rect 9861 3139 9919 3145
rect 10962 3136 10968 3188
rect 11020 3176 11026 3188
rect 12342 3176 12348 3188
rect 11020 3148 12348 3176
rect 11020 3136 11026 3148
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12618 3136 12624 3188
rect 12676 3176 12682 3188
rect 13262 3176 13268 3188
rect 12676 3148 13268 3176
rect 12676 3136 12682 3148
rect 13262 3136 13268 3148
rect 13320 3136 13326 3188
rect 13722 3176 13728 3188
rect 13683 3148 13728 3176
rect 13722 3136 13728 3148
rect 13780 3176 13786 3188
rect 13998 3176 14004 3188
rect 13780 3148 14004 3176
rect 13780 3136 13786 3148
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 14366 3136 14372 3188
rect 14424 3176 14430 3188
rect 14645 3179 14703 3185
rect 14645 3176 14657 3179
rect 14424 3148 14657 3176
rect 14424 3136 14430 3148
rect 14645 3145 14657 3148
rect 14691 3176 14703 3179
rect 14734 3176 14740 3188
rect 14691 3148 14740 3176
rect 14691 3145 14703 3148
rect 14645 3139 14703 3145
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 14829 3179 14887 3185
rect 14829 3145 14841 3179
rect 14875 3176 14887 3179
rect 15010 3176 15016 3188
rect 14875 3148 15016 3176
rect 14875 3145 14887 3148
rect 14829 3139 14887 3145
rect 15010 3136 15016 3148
rect 15068 3136 15074 3188
rect 16114 3176 16120 3188
rect 15120 3148 16120 3176
rect 12066 3108 12072 3120
rect 12027 3080 12072 3108
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 12529 3111 12587 3117
rect 12529 3077 12541 3111
rect 12575 3108 12587 3111
rect 13817 3111 13875 3117
rect 12575 3080 13768 3108
rect 12575 3077 12587 3080
rect 12529 3071 12587 3077
rect 13740 3052 13768 3080
rect 13817 3077 13829 3111
rect 13863 3108 13875 3111
rect 15120 3108 15148 3148
rect 16114 3136 16120 3148
rect 16172 3136 16178 3188
rect 16393 3179 16451 3185
rect 16393 3145 16405 3179
rect 16439 3176 16451 3179
rect 17126 3176 17132 3188
rect 16439 3148 17132 3176
rect 16439 3145 16451 3148
rect 16393 3139 16451 3145
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 18233 3179 18291 3185
rect 17276 3148 17908 3176
rect 17276 3136 17282 3148
rect 15657 3111 15715 3117
rect 15657 3108 15669 3111
rect 13863 3080 15148 3108
rect 15304 3080 15669 3108
rect 13863 3077 13875 3080
rect 13817 3071 13875 3077
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3040 2375 3043
rect 3326 3040 3332 3052
rect 2363 3012 3332 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 6273 3043 6331 3049
rect 6273 3040 6285 3043
rect 5776 3012 6285 3040
rect 5776 3000 5782 3012
rect 6273 3009 6285 3012
rect 6319 3040 6331 3043
rect 6362 3040 6368 3052
rect 6319 3012 6368 3040
rect 6319 3009 6331 3012
rect 6273 3003 6331 3009
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 10226 3040 10232 3052
rect 10060 3012 10232 3040
rect 1486 2932 1492 2984
rect 1544 2972 1550 2984
rect 2041 2975 2099 2981
rect 2041 2972 2053 2975
rect 1544 2944 2053 2972
rect 1544 2932 1550 2944
rect 2041 2941 2053 2944
rect 2087 2941 2099 2975
rect 2041 2935 2099 2941
rect 3786 2932 3792 2984
rect 3844 2972 3850 2984
rect 3881 2975 3939 2981
rect 3881 2972 3893 2975
rect 3844 2944 3893 2972
rect 3844 2932 3850 2944
rect 3881 2941 3893 2944
rect 3927 2941 3939 2975
rect 5810 2972 5816 2984
rect 3881 2935 3939 2941
rect 4080 2944 5816 2972
rect 1670 2864 1676 2916
rect 1728 2904 1734 2916
rect 4080 2904 4108 2944
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 6730 2932 6736 2984
rect 6788 2972 6794 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6788 2944 6837 2972
rect 6788 2932 6794 2944
rect 6825 2941 6837 2944
rect 6871 2972 6883 2975
rect 8481 2975 8539 2981
rect 8481 2972 8493 2975
rect 6871 2944 8493 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 8481 2941 8493 2944
rect 8527 2972 8539 2975
rect 8570 2972 8576 2984
rect 8527 2944 8576 2972
rect 8527 2941 8539 2944
rect 8481 2935 8539 2941
rect 8570 2932 8576 2944
rect 8628 2932 8634 2984
rect 8748 2975 8806 2981
rect 8748 2941 8760 2975
rect 8794 2972 8806 2975
rect 10060 2972 10088 3012
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 11974 3000 11980 3052
rect 12032 3040 12038 3052
rect 13078 3040 13084 3052
rect 12032 3012 12296 3040
rect 13039 3012 13084 3040
rect 12032 3000 12038 3012
rect 8794 2944 10088 2972
rect 8794 2941 8806 2944
rect 8748 2935 8806 2941
rect 10134 2932 10140 2984
rect 10192 2972 10198 2984
rect 10689 2975 10747 2981
rect 10192 2944 10237 2972
rect 10192 2932 10198 2944
rect 10689 2941 10701 2975
rect 10735 2972 10747 2975
rect 10778 2972 10784 2984
rect 10735 2944 10784 2972
rect 10735 2941 10747 2944
rect 10689 2935 10747 2941
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 10956 2975 11014 2981
rect 10956 2941 10968 2975
rect 11002 2972 11014 2975
rect 12158 2972 12164 2984
rect 11002 2944 12164 2972
rect 11002 2941 11014 2944
rect 10956 2935 11014 2941
rect 12158 2932 12164 2944
rect 12216 2932 12222 2984
rect 12268 2972 12296 3012
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3040 13323 3043
rect 13354 3040 13360 3052
rect 13311 3012 13360 3040
rect 13311 3009 13323 3012
rect 13265 3003 13323 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 13722 3000 13728 3052
rect 13780 3000 13786 3052
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 14277 3043 14335 3049
rect 14277 3040 14289 3043
rect 14056 3012 14289 3040
rect 14056 3000 14062 3012
rect 14277 3009 14289 3012
rect 14323 3009 14335 3043
rect 14458 3040 14464 3052
rect 14419 3012 14464 3040
rect 14277 3003 14335 3009
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 14734 3000 14740 3052
rect 14792 3040 14798 3052
rect 15304 3049 15332 3080
rect 15657 3077 15669 3080
rect 15703 3077 15715 3111
rect 15657 3071 15715 3077
rect 16025 3111 16083 3117
rect 16025 3077 16037 3111
rect 16071 3108 16083 3111
rect 17770 3108 17776 3120
rect 16071 3080 17776 3108
rect 16071 3077 16083 3080
rect 16025 3071 16083 3077
rect 17770 3068 17776 3080
rect 17828 3068 17834 3120
rect 17880 3108 17908 3148
rect 18233 3145 18245 3179
rect 18279 3176 18291 3179
rect 18506 3176 18512 3188
rect 18279 3148 18512 3176
rect 18279 3145 18291 3148
rect 18233 3139 18291 3145
rect 18506 3136 18512 3148
rect 18564 3136 18570 3188
rect 19426 3176 19432 3188
rect 19387 3148 19432 3176
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 19610 3136 19616 3188
rect 19668 3176 19674 3188
rect 20438 3176 20444 3188
rect 19668 3148 20444 3176
rect 19668 3136 19674 3148
rect 20438 3136 20444 3148
rect 20496 3136 20502 3188
rect 20714 3136 20720 3188
rect 20772 3136 20778 3188
rect 20070 3108 20076 3120
rect 17880 3080 20076 3108
rect 20070 3068 20076 3080
rect 20128 3068 20134 3120
rect 20732 3108 20760 3136
rect 20180 3080 20760 3108
rect 15289 3043 15347 3049
rect 15289 3040 15301 3043
rect 14792 3012 15301 3040
rect 14792 3000 14798 3012
rect 15289 3009 15301 3012
rect 15335 3009 15347 3043
rect 15289 3003 15347 3009
rect 15473 3043 15531 3049
rect 15473 3009 15485 3043
rect 15519 3040 15531 3043
rect 16390 3040 16396 3052
rect 15519 3012 16396 3040
rect 15519 3009 15531 3012
rect 15473 3003 15531 3009
rect 16390 3000 16396 3012
rect 16448 3040 16454 3052
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 16448 3012 17049 3040
rect 16448 3000 16454 3012
rect 17037 3009 17049 3012
rect 17083 3040 17095 3043
rect 17126 3040 17132 3052
rect 17083 3012 17132 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 17494 3000 17500 3052
rect 17552 3040 17558 3052
rect 18877 3043 18935 3049
rect 17552 3012 18828 3040
rect 17552 3000 17558 3012
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 12268 2944 13001 2972
rect 12989 2941 13001 2944
rect 13035 2941 13047 2975
rect 12989 2935 13047 2941
rect 13538 2932 13544 2984
rect 13596 2972 13602 2984
rect 14185 2975 14243 2981
rect 14185 2972 14197 2975
rect 13596 2944 14197 2972
rect 13596 2932 13602 2944
rect 14185 2941 14197 2944
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 15102 2932 15108 2984
rect 15160 2972 15166 2984
rect 15197 2975 15255 2981
rect 15197 2972 15209 2975
rect 15160 2944 15209 2972
rect 15160 2932 15166 2944
rect 15197 2941 15209 2944
rect 15243 2941 15255 2975
rect 15197 2935 15255 2941
rect 15378 2932 15384 2984
rect 15436 2972 15442 2984
rect 15841 2975 15899 2981
rect 15841 2972 15853 2975
rect 15436 2944 15853 2972
rect 15436 2932 15442 2944
rect 15841 2941 15853 2944
rect 15887 2941 15899 2975
rect 16758 2972 16764 2984
rect 16719 2944 16764 2972
rect 15841 2935 15899 2941
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 16850 2932 16856 2984
rect 16908 2972 16914 2984
rect 17402 2972 17408 2984
rect 16908 2944 16953 2972
rect 17363 2944 17408 2972
rect 16908 2932 16914 2944
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 4154 2913 4160 2916
rect 1728 2876 4108 2904
rect 1728 2864 1734 2876
rect 4148 2867 4160 2913
rect 4212 2904 4218 2916
rect 6086 2904 6092 2916
rect 4212 2876 4248 2904
rect 6047 2876 6092 2904
rect 4154 2864 4160 2867
rect 4212 2864 4218 2876
rect 6086 2864 6092 2876
rect 6144 2864 6150 2916
rect 7092 2907 7150 2913
rect 7092 2873 7104 2907
rect 7138 2904 7150 2907
rect 7190 2904 7196 2916
rect 7138 2876 7196 2904
rect 7138 2873 7150 2876
rect 7092 2867 7150 2873
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 9582 2904 9588 2916
rect 8680 2876 9588 2904
rect 2038 2796 2044 2848
rect 2096 2836 2102 2848
rect 2133 2839 2191 2845
rect 2133 2836 2145 2839
rect 2096 2808 2145 2836
rect 2096 2796 2102 2808
rect 2133 2805 2145 2808
rect 2179 2805 2191 2839
rect 2133 2799 2191 2805
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3053 2839 3111 2845
rect 3053 2836 3065 2839
rect 2832 2808 3065 2836
rect 2832 2796 2838 2808
rect 3053 2805 3065 2808
rect 3099 2805 3111 2839
rect 3053 2799 3111 2805
rect 3142 2796 3148 2848
rect 3200 2836 3206 2848
rect 3200 2808 3245 2836
rect 3200 2796 3206 2808
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 5350 2836 5356 2848
rect 4304 2808 5356 2836
rect 4304 2796 4310 2808
rect 5350 2796 5356 2808
rect 5408 2796 5414 2848
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 6914 2836 6920 2848
rect 6227 2808 6920 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 8680 2836 8708 2876
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 9858 2864 9864 2916
rect 9916 2904 9922 2916
rect 11238 2904 11244 2916
rect 9916 2876 11244 2904
rect 9916 2864 9922 2876
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 18322 2904 18328 2916
rect 11348 2876 18328 2904
rect 8444 2808 8708 2836
rect 8444 2796 8450 2808
rect 8754 2796 8760 2848
rect 8812 2836 8818 2848
rect 9306 2836 9312 2848
rect 8812 2808 9312 2836
rect 8812 2796 8818 2808
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 10042 2796 10048 2848
rect 10100 2836 10106 2848
rect 10226 2836 10232 2848
rect 10100 2808 10232 2836
rect 10100 2796 10106 2808
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 10321 2839 10379 2845
rect 10321 2805 10333 2839
rect 10367 2836 10379 2839
rect 11348 2836 11376 2876
rect 18322 2864 18328 2876
rect 18380 2864 18386 2916
rect 18598 2904 18604 2916
rect 18559 2876 18604 2904
rect 18598 2864 18604 2876
rect 18656 2864 18662 2916
rect 10367 2808 11376 2836
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 11422 2796 11428 2848
rect 11480 2836 11486 2848
rect 11974 2836 11980 2848
rect 11480 2808 11980 2836
rect 11480 2796 11486 2808
rect 11974 2796 11980 2808
rect 12032 2796 12038 2848
rect 12529 2839 12587 2845
rect 12529 2805 12541 2839
rect 12575 2836 12587 2839
rect 12621 2839 12679 2845
rect 12621 2836 12633 2839
rect 12575 2808 12633 2836
rect 12575 2805 12587 2808
rect 12529 2799 12587 2805
rect 12621 2805 12633 2808
rect 12667 2805 12679 2839
rect 12621 2799 12679 2805
rect 17589 2839 17647 2845
rect 17589 2805 17601 2839
rect 17635 2836 17647 2839
rect 18414 2836 18420 2848
rect 17635 2808 18420 2836
rect 17635 2805 17647 2808
rect 17589 2799 17647 2805
rect 18414 2796 18420 2808
rect 18472 2796 18478 2848
rect 18690 2836 18696 2848
rect 18651 2808 18696 2836
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 18800 2836 18828 3012
rect 18877 3009 18889 3043
rect 18923 3040 18935 3043
rect 18966 3040 18972 3052
rect 18923 3012 18972 3040
rect 18923 3009 18935 3012
rect 18877 3003 18935 3009
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 19794 3000 19800 3052
rect 19852 3040 19858 3052
rect 19981 3043 20039 3049
rect 19981 3040 19993 3043
rect 19852 3012 19993 3040
rect 19852 3000 19858 3012
rect 19981 3009 19993 3012
rect 20027 3009 20039 3043
rect 20180 3040 20208 3080
rect 19981 3003 20039 3009
rect 20088 3012 20208 3040
rect 19242 2932 19248 2984
rect 19300 2972 19306 2984
rect 19334 2972 19340 2984
rect 19300 2944 19340 2972
rect 19300 2932 19306 2944
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 19889 2975 19947 2981
rect 19889 2941 19901 2975
rect 19935 2972 19947 2975
rect 20088 2972 20116 3012
rect 20438 2972 20444 2984
rect 19935 2944 20116 2972
rect 20399 2944 20444 2972
rect 19935 2941 19947 2944
rect 19889 2935 19947 2941
rect 20438 2932 20444 2944
rect 20496 2932 20502 2984
rect 22554 2972 22560 2984
rect 20640 2944 22560 2972
rect 20640 2916 20668 2944
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 19797 2907 19855 2913
rect 19797 2873 19809 2907
rect 19843 2904 19855 2907
rect 20530 2904 20536 2916
rect 19843 2876 20536 2904
rect 19843 2873 19855 2876
rect 19797 2867 19855 2873
rect 20530 2864 20536 2876
rect 20588 2864 20594 2916
rect 20622 2864 20628 2916
rect 20680 2864 20686 2916
rect 20717 2907 20775 2913
rect 20717 2873 20729 2907
rect 20763 2904 20775 2907
rect 22186 2904 22192 2916
rect 20763 2876 22192 2904
rect 20763 2873 20775 2876
rect 20717 2867 20775 2873
rect 22186 2864 22192 2876
rect 22244 2864 22250 2916
rect 19242 2836 19248 2848
rect 18800 2808 19248 2836
rect 19242 2796 19248 2808
rect 19300 2796 19306 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1394 2592 1400 2644
rect 1452 2632 1458 2644
rect 1949 2635 2007 2641
rect 1949 2632 1961 2635
rect 1452 2604 1961 2632
rect 1452 2592 1458 2604
rect 1949 2601 1961 2604
rect 1995 2601 2007 2635
rect 1949 2595 2007 2601
rect 2130 2592 2136 2644
rect 2188 2632 2194 2644
rect 2317 2635 2375 2641
rect 2317 2632 2329 2635
rect 2188 2604 2329 2632
rect 2188 2592 2194 2604
rect 2317 2601 2329 2604
rect 2363 2601 2375 2635
rect 2317 2595 2375 2601
rect 2961 2635 3019 2641
rect 2961 2601 2973 2635
rect 3007 2632 3019 2635
rect 3142 2632 3148 2644
rect 3007 2604 3148 2632
rect 3007 2601 3019 2604
rect 2961 2595 3019 2601
rect 3142 2592 3148 2604
rect 3200 2592 3206 2644
rect 3326 2632 3332 2644
rect 3287 2604 3332 2632
rect 3326 2592 3332 2604
rect 3384 2632 3390 2644
rect 4706 2632 4712 2644
rect 3384 2604 4712 2632
rect 3384 2592 3390 2604
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 5445 2635 5503 2641
rect 5445 2601 5457 2635
rect 5491 2632 5503 2635
rect 5626 2632 5632 2644
rect 5491 2604 5632 2632
rect 5491 2601 5503 2604
rect 5445 2595 5503 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2632 5871 2635
rect 6546 2632 6552 2644
rect 5859 2604 6552 2632
rect 5859 2601 5871 2604
rect 5813 2595 5871 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 6914 2632 6920 2644
rect 6875 2604 6920 2632
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7285 2635 7343 2641
rect 7285 2632 7297 2635
rect 7248 2604 7297 2632
rect 7248 2592 7254 2604
rect 7285 2601 7297 2604
rect 7331 2601 7343 2635
rect 7285 2595 7343 2601
rect 10137 2635 10195 2641
rect 10137 2601 10149 2635
rect 10183 2632 10195 2635
rect 10183 2604 10548 2632
rect 10183 2601 10195 2604
rect 10137 2595 10195 2601
rect 1854 2524 1860 2576
rect 1912 2564 1918 2576
rect 2409 2567 2467 2573
rect 2409 2564 2421 2567
rect 1912 2536 2421 2564
rect 1912 2524 1918 2536
rect 2409 2533 2421 2536
rect 2455 2533 2467 2567
rect 2409 2527 2467 2533
rect 2700 2536 3188 2564
rect 1946 2456 1952 2508
rect 2004 2496 2010 2508
rect 2700 2496 2728 2536
rect 2004 2468 2728 2496
rect 3160 2496 3188 2536
rect 3234 2524 3240 2576
rect 3292 2564 3298 2576
rect 4310 2567 4368 2573
rect 4310 2564 4322 2567
rect 3292 2536 4322 2564
rect 3292 2524 3298 2536
rect 4310 2533 4322 2536
rect 4356 2533 4368 2567
rect 4310 2527 4368 2533
rect 6181 2567 6239 2573
rect 6181 2533 6193 2567
rect 6227 2564 6239 2567
rect 7650 2564 7656 2576
rect 6227 2536 7656 2564
rect 6227 2533 6239 2536
rect 6181 2527 6239 2533
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 8110 2524 8116 2576
rect 8168 2564 8174 2576
rect 8297 2567 8355 2573
rect 8297 2564 8309 2567
rect 8168 2536 8309 2564
rect 8168 2524 8174 2536
rect 8297 2533 8309 2536
rect 8343 2564 8355 2567
rect 8478 2564 8484 2576
rect 8343 2536 8484 2564
rect 8343 2533 8355 2536
rect 8297 2527 8355 2533
rect 8478 2524 8484 2536
rect 8536 2524 8542 2576
rect 9306 2524 9312 2576
rect 9364 2564 9370 2576
rect 9364 2536 10456 2564
rect 9364 2524 9370 2536
rect 3786 2496 3792 2508
rect 3160 2468 3792 2496
rect 2004 2456 2010 2468
rect 3786 2456 3792 2468
rect 3844 2496 3850 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3844 2468 4077 2496
rect 3844 2456 3850 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4154 2456 4160 2508
rect 4212 2496 4218 2508
rect 5074 2496 5080 2508
rect 4212 2468 5080 2496
rect 4212 2456 4218 2468
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 7377 2499 7435 2505
rect 7377 2496 7389 2499
rect 5868 2468 7389 2496
rect 5868 2456 5874 2468
rect 7377 2465 7389 2468
rect 7423 2496 7435 2499
rect 8202 2496 8208 2508
rect 7423 2468 8208 2496
rect 7423 2465 7435 2468
rect 7377 2459 7435 2465
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 8386 2496 8392 2508
rect 8347 2468 8392 2496
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 8846 2496 8852 2508
rect 8588 2468 8852 2496
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2682 2428 2688 2440
rect 2639 2400 2688 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2682 2388 2688 2400
rect 2740 2388 2746 2440
rect 3418 2428 3424 2440
rect 3379 2400 3424 2428
rect 3418 2388 3424 2400
rect 3476 2388 3482 2440
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 4172 2428 4200 2456
rect 3651 2400 4200 2428
rect 6273 2431 6331 2437
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 6273 2397 6285 2431
rect 6319 2397 6331 2431
rect 6273 2391 6331 2397
rect 6288 2360 6316 2391
rect 6362 2388 6368 2440
rect 6420 2428 6426 2440
rect 8588 2437 8616 2468
rect 8846 2456 8852 2468
rect 8904 2456 8910 2508
rect 9122 2496 9128 2508
rect 9083 2468 9128 2496
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 9950 2456 9956 2508
rect 10008 2496 10014 2508
rect 10008 2468 10364 2496
rect 10008 2456 10014 2468
rect 7561 2431 7619 2437
rect 6420 2400 6465 2428
rect 6420 2388 6426 2400
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 7607 2400 8585 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 8662 2388 8668 2440
rect 8720 2428 8726 2440
rect 10336 2437 10364 2468
rect 10229 2431 10287 2437
rect 10229 2428 10241 2431
rect 8720 2400 10241 2428
rect 8720 2388 8726 2400
rect 10229 2397 10241 2400
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 7929 2363 7987 2369
rect 7929 2360 7941 2363
rect 6288 2332 7941 2360
rect 7929 2329 7941 2332
rect 7975 2329 7987 2363
rect 7929 2323 7987 2329
rect 8294 2320 8300 2372
rect 8352 2360 8358 2372
rect 9769 2363 9827 2369
rect 9769 2360 9781 2363
rect 8352 2332 9781 2360
rect 8352 2320 8358 2332
rect 9769 2329 9781 2332
rect 9815 2329 9827 2363
rect 10428 2360 10456 2536
rect 10520 2496 10548 2604
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11241 2635 11299 2641
rect 11241 2632 11253 2635
rect 11112 2604 11253 2632
rect 11112 2592 11118 2604
rect 11241 2601 11253 2604
rect 11287 2601 11299 2635
rect 14274 2632 14280 2644
rect 11241 2595 11299 2601
rect 11808 2604 14280 2632
rect 11149 2567 11207 2573
rect 11149 2533 11161 2567
rect 11195 2564 11207 2567
rect 11808 2564 11836 2604
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 14369 2635 14427 2641
rect 14369 2601 14381 2635
rect 14415 2632 14427 2635
rect 16209 2635 16267 2641
rect 14415 2604 15884 2632
rect 14415 2601 14427 2604
rect 14369 2595 14427 2601
rect 11195 2536 11836 2564
rect 12069 2567 12127 2573
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 12250 2564 12256 2576
rect 12115 2536 12256 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 12250 2524 12256 2536
rect 12308 2524 12314 2576
rect 12897 2567 12955 2573
rect 12897 2533 12909 2567
rect 12943 2564 12955 2567
rect 13170 2564 13176 2576
rect 12943 2536 13176 2564
rect 12943 2533 12955 2536
rect 12897 2527 12955 2533
rect 13170 2524 13176 2536
rect 13228 2524 13234 2576
rect 13354 2524 13360 2576
rect 13412 2564 13418 2576
rect 13412 2536 14044 2564
rect 13412 2524 13418 2536
rect 10962 2496 10968 2508
rect 10520 2468 10968 2496
rect 10962 2456 10968 2468
rect 11020 2496 11026 2508
rect 11330 2496 11336 2508
rect 11020 2468 11336 2496
rect 11020 2456 11026 2468
rect 11330 2456 11336 2468
rect 11388 2456 11394 2508
rect 11790 2496 11796 2508
rect 11751 2468 11796 2496
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 13446 2496 13452 2508
rect 12667 2468 13452 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 13446 2456 13452 2468
rect 13504 2456 13510 2508
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2496 13783 2499
rect 13906 2496 13912 2508
rect 13771 2468 13912 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 13906 2456 13912 2468
rect 13964 2456 13970 2508
rect 11425 2431 11483 2437
rect 11425 2397 11437 2431
rect 11471 2428 11483 2431
rect 11698 2428 11704 2440
rect 11471 2400 11704 2428
rect 11471 2397 11483 2400
rect 11425 2391 11483 2397
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 14016 2437 14044 2536
rect 14090 2524 14096 2576
rect 14148 2564 14154 2576
rect 15749 2567 15807 2573
rect 15749 2564 15761 2567
rect 14148 2536 15761 2564
rect 14148 2524 14154 2536
rect 15749 2533 15761 2536
rect 15795 2533 15807 2567
rect 15856 2564 15884 2604
rect 16209 2601 16221 2635
rect 16255 2632 16267 2635
rect 16298 2632 16304 2644
rect 16255 2604 16304 2632
rect 16255 2601 16267 2604
rect 16209 2595 16267 2601
rect 16298 2592 16304 2604
rect 16356 2592 16362 2644
rect 16666 2632 16672 2644
rect 16627 2604 16672 2632
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 17126 2592 17132 2644
rect 17184 2632 17190 2644
rect 17494 2632 17500 2644
rect 17184 2604 17500 2632
rect 17184 2592 17190 2604
rect 17494 2592 17500 2604
rect 17552 2592 17558 2644
rect 17678 2592 17684 2644
rect 17736 2632 17742 2644
rect 17862 2632 17868 2644
rect 17736 2604 17868 2632
rect 17736 2592 17742 2604
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 18230 2592 18236 2644
rect 18288 2632 18294 2644
rect 18325 2635 18383 2641
rect 18325 2632 18337 2635
rect 18288 2604 18337 2632
rect 18288 2592 18294 2604
rect 18325 2601 18337 2604
rect 18371 2601 18383 2635
rect 18325 2595 18383 2601
rect 18785 2635 18843 2641
rect 18785 2601 18797 2635
rect 18831 2632 18843 2635
rect 19150 2632 19156 2644
rect 18831 2604 19156 2632
rect 18831 2601 18843 2604
rect 18785 2595 18843 2601
rect 19150 2592 19156 2604
rect 19208 2592 19214 2644
rect 19337 2635 19395 2641
rect 19337 2601 19349 2635
rect 19383 2632 19395 2635
rect 19518 2632 19524 2644
rect 19383 2604 19524 2632
rect 19383 2601 19395 2604
rect 19337 2595 19395 2601
rect 19518 2592 19524 2604
rect 19576 2592 19582 2644
rect 19702 2632 19708 2644
rect 19663 2604 19708 2632
rect 19702 2592 19708 2604
rect 19760 2592 19766 2644
rect 17589 2567 17647 2573
rect 17589 2564 17601 2567
rect 15856 2536 17601 2564
rect 15749 2527 15807 2533
rect 17589 2533 17601 2536
rect 17635 2533 17647 2567
rect 19058 2564 19064 2576
rect 17589 2527 17647 2533
rect 17788 2536 19064 2564
rect 14734 2496 14740 2508
rect 14695 2468 14740 2496
rect 14734 2456 14740 2468
rect 14792 2456 14798 2508
rect 14826 2456 14832 2508
rect 14884 2496 14890 2508
rect 15286 2496 15292 2508
rect 14884 2468 14929 2496
rect 15028 2468 15292 2496
rect 14884 2456 14890 2468
rect 15028 2437 15056 2468
rect 15286 2456 15292 2468
rect 15344 2456 15350 2508
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 16577 2499 16635 2505
rect 16577 2465 16589 2499
rect 16623 2496 16635 2499
rect 17788 2496 17816 2536
rect 19058 2524 19064 2536
rect 19116 2524 19122 2576
rect 19242 2524 19248 2576
rect 19300 2564 19306 2576
rect 19797 2567 19855 2573
rect 19797 2564 19809 2567
rect 19300 2536 19809 2564
rect 19300 2524 19306 2536
rect 19797 2533 19809 2536
rect 19843 2533 19855 2567
rect 20622 2564 20628 2576
rect 20583 2536 20628 2564
rect 19797 2527 19855 2533
rect 20622 2524 20628 2536
rect 20680 2524 20686 2576
rect 18693 2499 18751 2505
rect 18693 2496 18705 2499
rect 16623 2468 17816 2496
rect 17972 2468 18705 2496
rect 16623 2465 16635 2468
rect 16577 2459 16635 2465
rect 13817 2431 13875 2437
rect 13817 2428 13829 2431
rect 13096 2400 13829 2428
rect 13096 2360 13124 2400
rect 13817 2397 13829 2400
rect 13863 2397 13875 2431
rect 13817 2391 13875 2397
rect 14001 2431 14059 2437
rect 14001 2397 14013 2431
rect 14047 2428 14059 2431
rect 15013 2431 15071 2437
rect 15013 2428 15025 2431
rect 14047 2400 15025 2428
rect 14047 2397 14059 2400
rect 14001 2391 14059 2397
rect 15013 2397 15025 2400
rect 15059 2397 15071 2431
rect 15013 2391 15071 2397
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2428 15255 2431
rect 15488 2428 15516 2459
rect 15243 2400 15516 2428
rect 15243 2397 15255 2400
rect 15197 2391 15255 2397
rect 16482 2388 16488 2440
rect 16540 2428 16546 2440
rect 16761 2431 16819 2437
rect 16761 2428 16773 2431
rect 16540 2400 16773 2428
rect 16540 2388 16546 2400
rect 16761 2397 16773 2400
rect 16807 2397 16819 2431
rect 16761 2391 16819 2397
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 17862 2428 17868 2440
rect 17823 2400 17868 2428
rect 17681 2391 17739 2397
rect 10428 2332 13124 2360
rect 13357 2363 13415 2369
rect 9769 2323 9827 2329
rect 13357 2329 13369 2363
rect 13403 2360 13415 2363
rect 17696 2360 17724 2391
rect 17862 2388 17868 2400
rect 17920 2388 17926 2440
rect 13403 2332 17724 2360
rect 13403 2329 13415 2332
rect 13357 2323 13415 2329
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 4798 2292 4804 2304
rect 3476 2264 4804 2292
rect 3476 2252 3482 2264
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 5902 2252 5908 2304
rect 5960 2292 5966 2304
rect 9122 2292 9128 2304
rect 5960 2264 9128 2292
rect 5960 2252 5966 2264
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 9309 2295 9367 2301
rect 9309 2261 9321 2295
rect 9355 2292 9367 2295
rect 9674 2292 9680 2304
rect 9355 2264 9680 2292
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 10778 2292 10784 2304
rect 10739 2264 10784 2292
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 12710 2252 12716 2304
rect 12768 2292 12774 2304
rect 15197 2295 15255 2301
rect 15197 2292 15209 2295
rect 12768 2264 15209 2292
rect 12768 2252 12774 2264
rect 15197 2261 15209 2264
rect 15243 2261 15255 2295
rect 17218 2292 17224 2304
rect 17179 2264 17224 2292
rect 15197 2255 15255 2261
rect 17218 2252 17224 2264
rect 17276 2252 17282 2304
rect 17310 2252 17316 2304
rect 17368 2292 17374 2304
rect 17972 2292 18000 2468
rect 18693 2465 18705 2468
rect 18739 2465 18751 2499
rect 18693 2459 18751 2465
rect 20070 2456 20076 2508
rect 20128 2496 20134 2508
rect 20349 2499 20407 2505
rect 20349 2496 20361 2499
rect 20128 2468 20361 2496
rect 20128 2456 20134 2468
rect 20349 2465 20361 2468
rect 20395 2465 20407 2499
rect 20349 2459 20407 2465
rect 18966 2428 18972 2440
rect 18927 2400 18972 2428
rect 18966 2388 18972 2400
rect 19024 2388 19030 2440
rect 19886 2428 19892 2440
rect 19847 2400 19892 2428
rect 19886 2388 19892 2400
rect 19944 2388 19950 2440
rect 18322 2320 18328 2372
rect 18380 2360 18386 2372
rect 21450 2360 21456 2372
rect 18380 2332 21456 2360
rect 18380 2320 18386 2332
rect 21450 2320 21456 2332
rect 21508 2320 21514 2372
rect 17368 2264 18000 2292
rect 17368 2252 17374 2264
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 5074 2048 5080 2100
rect 5132 2088 5138 2100
rect 9950 2088 9956 2100
rect 5132 2060 9956 2088
rect 5132 2048 5138 2060
rect 9950 2048 9956 2060
rect 10008 2048 10014 2100
rect 10778 2048 10784 2100
rect 10836 2088 10842 2100
rect 10836 2060 14228 2088
rect 10836 2048 10842 2060
rect 198 1980 204 2032
rect 256 2020 262 2032
rect 8386 2020 8392 2032
rect 256 1992 8392 2020
rect 256 1980 262 1992
rect 8386 1980 8392 1992
rect 8444 1980 8450 2032
rect 2038 1912 2044 1964
rect 2096 1952 2102 1964
rect 7190 1952 7196 1964
rect 2096 1924 7196 1952
rect 2096 1912 2102 1924
rect 7190 1912 7196 1924
rect 7248 1912 7254 1964
rect 14200 1952 14228 2060
rect 14734 2048 14740 2100
rect 14792 2088 14798 2100
rect 20898 2088 20904 2100
rect 14792 2060 20904 2088
rect 14792 2048 14798 2060
rect 20898 2048 20904 2060
rect 20956 2048 20962 2100
rect 14274 1980 14280 2032
rect 14332 2020 14338 2032
rect 18966 2020 18972 2032
rect 14332 1992 18972 2020
rect 14332 1980 14338 1992
rect 18966 1980 18972 1992
rect 19024 1980 19030 2032
rect 20254 1952 20260 1964
rect 14200 1924 20260 1952
rect 20254 1912 20260 1924
rect 20312 1912 20318 1964
rect 1302 1844 1308 1896
rect 1360 1884 1366 1896
rect 7558 1884 7564 1896
rect 1360 1856 7564 1884
rect 1360 1844 1366 1856
rect 7558 1844 7564 1856
rect 7616 1844 7622 1896
rect 7742 1844 7748 1896
rect 7800 1884 7806 1896
rect 14826 1884 14832 1896
rect 7800 1856 14832 1884
rect 7800 1844 7806 1856
rect 14826 1844 14832 1856
rect 14884 1844 14890 1896
rect 15470 1844 15476 1896
rect 15528 1884 15534 1896
rect 17402 1884 17408 1896
rect 15528 1856 17408 1884
rect 15528 1844 15534 1856
rect 17402 1844 17408 1856
rect 17460 1844 17466 1896
rect 5350 1776 5356 1828
rect 5408 1816 5414 1828
rect 7374 1816 7380 1828
rect 5408 1788 7380 1816
rect 5408 1776 5414 1788
rect 7374 1776 7380 1788
rect 7432 1816 7438 1828
rect 17310 1816 17316 1828
rect 7432 1788 17316 1816
rect 7432 1776 7438 1788
rect 17310 1776 17316 1788
rect 17368 1776 17374 1828
rect 566 1708 572 1760
rect 624 1748 630 1760
rect 8110 1748 8116 1760
rect 624 1720 8116 1748
rect 624 1708 630 1720
rect 8110 1708 8116 1720
rect 8168 1708 8174 1760
rect 12986 1708 12992 1760
rect 13044 1748 13050 1760
rect 15470 1748 15476 1760
rect 13044 1720 15476 1748
rect 13044 1708 13050 1720
rect 15470 1708 15476 1720
rect 15528 1708 15534 1760
rect 2406 1640 2412 1692
rect 2464 1680 2470 1692
rect 7098 1680 7104 1692
rect 2464 1652 7104 1680
rect 2464 1640 2470 1652
rect 7098 1640 7104 1652
rect 7156 1640 7162 1692
rect 2774 1572 2780 1624
rect 2832 1612 2838 1624
rect 6822 1612 6828 1624
rect 2832 1584 6828 1612
rect 2832 1572 2838 1584
rect 6822 1572 6828 1584
rect 6880 1572 6886 1624
rect 9674 1368 9680 1420
rect 9732 1408 9738 1420
rect 15102 1408 15108 1420
rect 9732 1380 15108 1408
rect 9732 1368 9738 1380
rect 15102 1368 15108 1380
rect 15160 1368 15166 1420
rect 16758 1300 16764 1352
rect 16816 1340 16822 1352
rect 17954 1340 17960 1352
rect 16816 1312 17960 1340
rect 16816 1300 16822 1312
rect 17954 1300 17960 1312
rect 18012 1300 18018 1352
rect 12802 1232 12808 1284
rect 12860 1272 12866 1284
rect 14366 1272 14372 1284
rect 12860 1244 14372 1272
rect 12860 1232 12866 1244
rect 14366 1232 14372 1244
rect 14424 1232 14430 1284
rect 16574 1096 16580 1148
rect 16632 1136 16638 1148
rect 17126 1136 17132 1148
rect 16632 1108 17132 1136
rect 16632 1096 16638 1108
rect 17126 1096 17132 1108
rect 17184 1096 17190 1148
<< via1 >>
rect 3884 21224 3936 21276
rect 8300 21224 8352 21276
rect 4068 20952 4120 21004
rect 6000 20952 6052 21004
rect 3792 20612 3844 20664
rect 11612 20612 11664 20664
rect 15292 20612 15344 20664
rect 19524 20612 19576 20664
rect 8760 20544 8812 20596
rect 19340 20544 19392 20596
rect 4988 20408 5040 20460
rect 12256 20408 12308 20460
rect 572 20272 624 20324
rect 5356 20272 5408 20324
rect 7564 20272 7616 20324
rect 15108 20272 15160 20324
rect 8484 20204 8536 20256
rect 8668 20204 8720 20256
rect 9312 20204 9364 20256
rect 14004 20204 14056 20256
rect 15016 20204 15068 20256
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 1952 19975 2004 19984
rect 1952 19941 1961 19975
rect 1961 19941 1995 19975
rect 1995 19941 2004 19975
rect 1952 19932 2004 19941
rect 2320 19864 2372 19916
rect 7564 20000 7616 20052
rect 7656 20000 7708 20052
rect 12716 20000 12768 20052
rect 13820 20000 13872 20052
rect 19064 20000 19116 20052
rect 3516 19864 3568 19916
rect 2780 19796 2832 19848
rect 4896 19864 4948 19916
rect 5356 19864 5408 19916
rect 6092 19907 6144 19916
rect 6092 19873 6101 19907
rect 6101 19873 6135 19907
rect 6135 19873 6144 19907
rect 6092 19864 6144 19873
rect 1676 19728 1728 19780
rect 3792 19728 3844 19780
rect 5264 19796 5316 19848
rect 5172 19728 5224 19780
rect 5356 19728 5408 19780
rect 4068 19703 4120 19712
rect 4068 19669 4077 19703
rect 4077 19669 4111 19703
rect 4111 19669 4120 19703
rect 4068 19660 4120 19669
rect 6184 19660 6236 19712
rect 6644 19796 6696 19848
rect 8024 19932 8076 19984
rect 8392 19864 8444 19916
rect 9036 19839 9088 19848
rect 9036 19805 9045 19839
rect 9045 19805 9079 19839
rect 9079 19805 9088 19839
rect 9036 19796 9088 19805
rect 9864 19932 9916 19984
rect 9496 19864 9548 19916
rect 12164 19932 12216 19984
rect 12256 19932 12308 19984
rect 15476 19932 15528 19984
rect 16580 19932 16632 19984
rect 12440 19864 12492 19916
rect 12624 19907 12676 19916
rect 12624 19873 12633 19907
rect 12633 19873 12667 19907
rect 12667 19873 12676 19907
rect 12624 19864 12676 19873
rect 13912 19907 13964 19916
rect 13912 19873 13921 19907
rect 13921 19873 13955 19907
rect 13955 19873 13964 19907
rect 13912 19864 13964 19873
rect 14464 19907 14516 19916
rect 14464 19873 14473 19907
rect 14473 19873 14507 19907
rect 14507 19873 14516 19907
rect 14464 19864 14516 19873
rect 15108 19864 15160 19916
rect 15660 19907 15712 19916
rect 15660 19873 15669 19907
rect 15669 19873 15703 19907
rect 15703 19873 15712 19907
rect 15660 19864 15712 19873
rect 19156 19975 19208 19984
rect 10232 19839 10284 19848
rect 10232 19805 10241 19839
rect 10241 19805 10275 19839
rect 10275 19805 10284 19839
rect 10232 19796 10284 19805
rect 10324 19839 10376 19848
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 10324 19796 10376 19805
rect 12072 19839 12124 19848
rect 12072 19805 12081 19839
rect 12081 19805 12115 19839
rect 12115 19805 12124 19839
rect 15844 19839 15896 19848
rect 12072 19796 12124 19805
rect 15844 19805 15853 19839
rect 15853 19805 15887 19839
rect 15887 19805 15896 19839
rect 15844 19796 15896 19805
rect 17224 19864 17276 19916
rect 8944 19728 8996 19780
rect 13452 19728 13504 19780
rect 15292 19728 15344 19780
rect 9680 19660 9732 19712
rect 12808 19660 12860 19712
rect 13820 19660 13872 19712
rect 17500 19728 17552 19780
rect 18788 19864 18840 19916
rect 19156 19941 19165 19975
rect 19165 19941 19199 19975
rect 19199 19941 19208 19975
rect 19156 19932 19208 19941
rect 21824 20000 21876 20052
rect 20628 19975 20680 19984
rect 20628 19941 20637 19975
rect 20637 19941 20671 19975
rect 20671 19941 20680 19975
rect 20628 19932 20680 19941
rect 19708 19864 19760 19916
rect 20352 19907 20404 19916
rect 20352 19873 20361 19907
rect 20361 19873 20395 19907
rect 20395 19873 20404 19907
rect 20352 19864 20404 19873
rect 22192 19796 22244 19848
rect 21456 19728 21508 19780
rect 18880 19660 18932 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 4068 19456 4120 19508
rect 6828 19456 6880 19508
rect 8392 19499 8444 19508
rect 8392 19465 8401 19499
rect 8401 19465 8435 19499
rect 8435 19465 8444 19499
rect 8392 19456 8444 19465
rect 8760 19456 8812 19508
rect 10324 19456 10376 19508
rect 12440 19499 12492 19508
rect 12440 19465 12449 19499
rect 12449 19465 12483 19499
rect 12483 19465 12492 19499
rect 12440 19456 12492 19465
rect 15660 19456 15712 19508
rect 16580 19456 16632 19508
rect 19156 19456 19208 19508
rect 3516 19320 3568 19372
rect 4252 19320 4304 19372
rect 16212 19388 16264 19440
rect 1676 19295 1728 19304
rect 1676 19261 1685 19295
rect 1685 19261 1719 19295
rect 1719 19261 1728 19295
rect 1676 19252 1728 19261
rect 1860 19252 1912 19304
rect 2044 19252 2096 19304
rect 4068 19252 4120 19304
rect 4160 19252 4212 19304
rect 1308 19184 1360 19236
rect 4344 19184 4396 19236
rect 6644 19320 6696 19372
rect 8024 19320 8076 19372
rect 5356 19252 5408 19304
rect 10140 19320 10192 19372
rect 10324 19320 10376 19372
rect 12072 19320 12124 19372
rect 13636 19320 13688 19372
rect 15108 19320 15160 19372
rect 15936 19320 15988 19372
rect 2780 19116 2832 19168
rect 2964 19116 3016 19168
rect 3516 19116 3568 19168
rect 3792 19159 3844 19168
rect 3792 19125 3801 19159
rect 3801 19125 3835 19159
rect 3835 19125 3844 19159
rect 3792 19116 3844 19125
rect 4896 19116 4948 19168
rect 5172 19116 5224 19168
rect 5356 19116 5408 19168
rect 7748 19184 7800 19236
rect 8116 19184 8168 19236
rect 9404 19252 9456 19304
rect 9680 19252 9732 19304
rect 12532 19252 12584 19304
rect 14924 19252 14976 19304
rect 9220 19184 9272 19236
rect 9956 19184 10008 19236
rect 6276 19116 6328 19168
rect 6460 19116 6512 19168
rect 10048 19116 10100 19168
rect 11796 19116 11848 19168
rect 14280 19184 14332 19236
rect 16120 19184 16172 19236
rect 16580 19252 16632 19304
rect 17224 19295 17276 19304
rect 17224 19261 17233 19295
rect 17233 19261 17267 19295
rect 17267 19261 17276 19295
rect 17224 19252 17276 19261
rect 18604 19320 18656 19372
rect 18972 19363 19024 19372
rect 18972 19329 18981 19363
rect 18981 19329 19015 19363
rect 19015 19329 19024 19363
rect 18972 19320 19024 19329
rect 19340 19320 19392 19372
rect 16672 19184 16724 19236
rect 17960 19252 18012 19304
rect 18144 19252 18196 19304
rect 18512 19184 18564 19236
rect 19800 19252 19852 19304
rect 19524 19184 19576 19236
rect 12716 19116 12768 19168
rect 13452 19116 13504 19168
rect 13544 19116 13596 19168
rect 14096 19159 14148 19168
rect 14096 19125 14105 19159
rect 14105 19125 14139 19159
rect 14139 19125 14148 19159
rect 14096 19116 14148 19125
rect 15016 19116 15068 19168
rect 15936 19159 15988 19168
rect 15936 19125 15945 19159
rect 15945 19125 15979 19159
rect 15979 19125 15988 19159
rect 15936 19116 15988 19125
rect 16396 19116 16448 19168
rect 17776 19116 17828 19168
rect 18972 19116 19024 19168
rect 19432 19116 19484 19168
rect 20812 19252 20864 19304
rect 20168 19116 20220 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 4712 18912 4764 18964
rect 4804 18912 4856 18964
rect 5816 18912 5868 18964
rect 6184 18955 6236 18964
rect 6184 18921 6193 18955
rect 6193 18921 6227 18955
rect 6227 18921 6236 18955
rect 6184 18912 6236 18921
rect 1952 18887 2004 18896
rect 1952 18853 1961 18887
rect 1961 18853 1995 18887
rect 1995 18853 2004 18887
rect 1952 18844 2004 18853
rect 5080 18844 5132 18896
rect 5724 18844 5776 18896
rect 8852 18844 8904 18896
rect 2320 18776 2372 18828
rect 2228 18708 2280 18760
rect 4160 18776 4212 18828
rect 4804 18776 4856 18828
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 7380 18776 7432 18828
rect 8760 18776 8812 18828
rect 10232 18912 10284 18964
rect 9404 18844 9456 18896
rect 10048 18887 10100 18896
rect 9680 18776 9732 18828
rect 10048 18853 10057 18887
rect 10057 18853 10091 18887
rect 10091 18853 10100 18887
rect 10048 18844 10100 18853
rect 14280 18912 14332 18964
rect 15292 18912 15344 18964
rect 15476 18912 15528 18964
rect 16212 18912 16264 18964
rect 19984 18912 20036 18964
rect 12992 18844 13044 18896
rect 14096 18844 14148 18896
rect 17132 18844 17184 18896
rect 18144 18887 18196 18896
rect 18144 18853 18153 18887
rect 18153 18853 18187 18887
rect 18187 18853 18196 18887
rect 18144 18844 18196 18853
rect 10600 18776 10652 18828
rect 11520 18776 11572 18828
rect 12072 18776 12124 18828
rect 12256 18776 12308 18828
rect 17224 18776 17276 18828
rect 17776 18776 17828 18828
rect 18696 18776 18748 18828
rect 3424 18751 3476 18760
rect 3424 18717 3433 18751
rect 3433 18717 3467 18751
rect 3467 18717 3476 18751
rect 3424 18708 3476 18717
rect 3516 18640 3568 18692
rect 2780 18572 2832 18624
rect 5172 18708 5224 18760
rect 6276 18751 6328 18760
rect 6276 18717 6285 18751
rect 6285 18717 6319 18751
rect 6319 18717 6328 18751
rect 6276 18708 6328 18717
rect 6644 18708 6696 18760
rect 9128 18751 9180 18760
rect 9128 18717 9137 18751
rect 9137 18717 9171 18751
rect 9171 18717 9180 18751
rect 9128 18708 9180 18717
rect 8484 18640 8536 18692
rect 10048 18708 10100 18760
rect 11152 18708 11204 18760
rect 5356 18572 5408 18624
rect 5724 18615 5776 18624
rect 5724 18581 5733 18615
rect 5733 18581 5767 18615
rect 5767 18581 5776 18615
rect 5724 18572 5776 18581
rect 5908 18572 5960 18624
rect 7288 18572 7340 18624
rect 7748 18572 7800 18624
rect 9220 18572 9272 18624
rect 10600 18640 10652 18692
rect 12900 18708 12952 18760
rect 9588 18572 9640 18624
rect 13820 18572 13872 18624
rect 14096 18572 14148 18624
rect 16212 18615 16264 18624
rect 16212 18581 16221 18615
rect 16221 18581 16255 18615
rect 16255 18581 16264 18615
rect 16212 18572 16264 18581
rect 17960 18572 18012 18624
rect 18972 18572 19024 18624
rect 19248 18844 19300 18896
rect 19340 18819 19392 18828
rect 19340 18785 19349 18819
rect 19349 18785 19383 18819
rect 19383 18785 19392 18819
rect 19340 18776 19392 18785
rect 19708 18776 19760 18828
rect 19248 18751 19300 18760
rect 19248 18717 19257 18751
rect 19257 18717 19291 18751
rect 19291 18717 19300 18751
rect 19248 18708 19300 18717
rect 22560 18708 22612 18760
rect 20352 18640 20404 18692
rect 20904 18572 20956 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 2228 18232 2280 18284
rect 4436 18300 4488 18352
rect 3516 18232 3568 18284
rect 5724 18368 5776 18420
rect 6000 18368 6052 18420
rect 7656 18368 7708 18420
rect 9036 18368 9088 18420
rect 9496 18411 9548 18420
rect 9496 18377 9505 18411
rect 9505 18377 9539 18411
rect 9539 18377 9548 18411
rect 9496 18368 9548 18377
rect 9588 18368 9640 18420
rect 9680 18368 9732 18420
rect 10048 18368 10100 18420
rect 12072 18411 12124 18420
rect 12072 18377 12081 18411
rect 12081 18377 12115 18411
rect 12115 18377 12124 18411
rect 12072 18368 12124 18377
rect 12624 18368 12676 18420
rect 12716 18368 12768 18420
rect 15936 18368 15988 18420
rect 16120 18411 16172 18420
rect 16120 18377 16129 18411
rect 16129 18377 16163 18411
rect 16163 18377 16172 18411
rect 16120 18368 16172 18377
rect 3792 18164 3844 18216
rect 4344 18164 4396 18216
rect 4712 18275 4764 18284
rect 4712 18241 4721 18275
rect 4721 18241 4755 18275
rect 4755 18241 4764 18275
rect 4712 18232 4764 18241
rect 2964 18096 3016 18148
rect 4528 18096 4580 18148
rect 4804 18096 4856 18148
rect 5356 18207 5408 18216
rect 5356 18173 5390 18207
rect 5390 18173 5408 18207
rect 5356 18164 5408 18173
rect 7748 18232 7800 18284
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 9220 18232 9272 18284
rect 9588 18164 9640 18216
rect 9772 18164 9824 18216
rect 10324 18164 10376 18216
rect 10600 18164 10652 18216
rect 13912 18300 13964 18352
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 13636 18232 13688 18284
rect 15476 18232 15528 18284
rect 15936 18232 15988 18284
rect 16764 18275 16816 18284
rect 16764 18241 16773 18275
rect 16773 18241 16807 18275
rect 16807 18241 16816 18275
rect 16764 18232 16816 18241
rect 12716 18164 12768 18216
rect 13820 18207 13872 18216
rect 13820 18173 13829 18207
rect 13829 18173 13863 18207
rect 13863 18173 13872 18207
rect 13820 18164 13872 18173
rect 18696 18368 18748 18420
rect 18512 18300 18564 18352
rect 20904 18232 20956 18284
rect 18420 18164 18472 18216
rect 18604 18164 18656 18216
rect 19340 18207 19392 18216
rect 19340 18173 19349 18207
rect 19349 18173 19383 18207
rect 19383 18173 19392 18207
rect 19340 18164 19392 18173
rect 19616 18164 19668 18216
rect 8576 18096 8628 18148
rect 9680 18096 9732 18148
rect 10140 18096 10192 18148
rect 11244 18096 11296 18148
rect 11796 18096 11848 18148
rect 13176 18096 13228 18148
rect 4344 18028 4396 18080
rect 4436 18071 4488 18080
rect 4436 18037 4445 18071
rect 4445 18037 4479 18071
rect 4479 18037 4488 18071
rect 4436 18028 4488 18037
rect 5356 18028 5408 18080
rect 6460 18071 6512 18080
rect 6460 18037 6469 18071
rect 6469 18037 6503 18071
rect 6503 18037 6512 18071
rect 6460 18028 6512 18037
rect 9772 18028 9824 18080
rect 10048 18028 10100 18080
rect 12532 18028 12584 18080
rect 14372 18028 14424 18080
rect 16304 18096 16356 18148
rect 19708 18096 19760 18148
rect 19800 18096 19852 18148
rect 16948 18028 17000 18080
rect 18420 18071 18472 18080
rect 18420 18037 18429 18071
rect 18429 18037 18463 18071
rect 18463 18037 18472 18071
rect 18420 18028 18472 18037
rect 20076 18071 20128 18080
rect 20076 18037 20085 18071
rect 20085 18037 20119 18071
rect 20119 18037 20128 18071
rect 20076 18028 20128 18037
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 204 17824 256 17876
rect 1860 17867 1912 17876
rect 1860 17833 1869 17867
rect 1869 17833 1903 17867
rect 1903 17833 1912 17867
rect 1860 17824 1912 17833
rect 2872 17867 2924 17876
rect 2872 17833 2881 17867
rect 2881 17833 2915 17867
rect 2915 17833 2924 17867
rect 2872 17824 2924 17833
rect 3056 17824 3108 17876
rect 3240 17824 3292 17876
rect 3424 17824 3476 17876
rect 4344 17824 4396 17876
rect 5080 17867 5132 17876
rect 5080 17833 5089 17867
rect 5089 17833 5123 17867
rect 5123 17833 5132 17867
rect 5080 17824 5132 17833
rect 6828 17867 6880 17876
rect 6828 17833 6837 17867
rect 6837 17833 6871 17867
rect 6871 17833 6880 17867
rect 6828 17824 6880 17833
rect 6920 17824 6972 17876
rect 7104 17824 7156 17876
rect 7380 17824 7432 17876
rect 8576 17867 8628 17876
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 8576 17824 8628 17833
rect 9128 17824 9180 17876
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 10048 17824 10100 17876
rect 13084 17867 13136 17876
rect 940 17688 992 17740
rect 1768 17731 1820 17740
rect 1768 17697 1777 17731
rect 1777 17697 1811 17731
rect 1811 17697 1820 17731
rect 1768 17688 1820 17697
rect 2596 17688 2648 17740
rect 3424 17731 3476 17740
rect 3424 17697 3433 17731
rect 3433 17697 3467 17731
rect 3467 17697 3476 17731
rect 3424 17688 3476 17697
rect 2504 17620 2556 17672
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 4528 17620 4580 17672
rect 5448 17731 5500 17740
rect 5448 17697 5457 17731
rect 5457 17697 5491 17731
rect 5491 17697 5500 17731
rect 5448 17688 5500 17697
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 6828 17688 6880 17740
rect 7196 17688 7248 17740
rect 7104 17663 7156 17672
rect 7104 17629 7113 17663
rect 7113 17629 7147 17663
rect 7147 17629 7156 17663
rect 7104 17620 7156 17629
rect 6092 17552 6144 17604
rect 11888 17756 11940 17808
rect 13084 17833 13093 17867
rect 13093 17833 13127 17867
rect 13127 17833 13136 17867
rect 13084 17824 13136 17833
rect 15936 17824 15988 17876
rect 16672 17824 16724 17876
rect 17500 17824 17552 17876
rect 8392 17688 8444 17740
rect 8668 17688 8720 17740
rect 8760 17688 8812 17740
rect 8300 17620 8352 17672
rect 9036 17663 9088 17672
rect 9036 17629 9045 17663
rect 9045 17629 9079 17663
rect 9079 17629 9088 17663
rect 9036 17620 9088 17629
rect 9404 17688 9456 17740
rect 10140 17663 10192 17672
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 10968 17688 11020 17740
rect 11244 17688 11296 17740
rect 12072 17688 12124 17740
rect 11888 17620 11940 17672
rect 12256 17663 12308 17672
rect 12256 17629 12265 17663
rect 12265 17629 12299 17663
rect 12299 17629 12308 17663
rect 12256 17620 12308 17629
rect 12532 17688 12584 17740
rect 13084 17688 13136 17740
rect 14648 17688 14700 17740
rect 15200 17688 15252 17740
rect 21456 17824 21508 17876
rect 20260 17756 20312 17808
rect 16580 17688 16632 17740
rect 19156 17731 19208 17740
rect 19156 17697 19165 17731
rect 19165 17697 19199 17731
rect 19199 17697 19208 17731
rect 19156 17688 19208 17697
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 15476 17620 15528 17672
rect 3148 17484 3200 17536
rect 7104 17484 7156 17536
rect 7840 17484 7892 17536
rect 11612 17484 11664 17536
rect 13176 17484 13228 17536
rect 15660 17484 15712 17536
rect 16764 17552 16816 17604
rect 17408 17552 17460 17604
rect 19248 17620 19300 17672
rect 19892 17620 19944 17672
rect 20444 17663 20496 17672
rect 20444 17629 20453 17663
rect 20453 17629 20487 17663
rect 20487 17629 20496 17663
rect 20444 17620 20496 17629
rect 20904 17620 20956 17672
rect 18604 17552 18656 17604
rect 21732 17552 21784 17604
rect 15936 17484 15988 17536
rect 16488 17484 16540 17536
rect 18880 17484 18932 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 2044 17280 2096 17332
rect 2780 17280 2832 17332
rect 3056 17280 3108 17332
rect 5540 17280 5592 17332
rect 7840 17280 7892 17332
rect 8300 17323 8352 17332
rect 8300 17289 8309 17323
rect 8309 17289 8343 17323
rect 8343 17289 8352 17323
rect 8300 17280 8352 17289
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 9772 17280 9824 17332
rect 12348 17280 12400 17332
rect 12440 17323 12492 17332
rect 12440 17289 12449 17323
rect 12449 17289 12483 17323
rect 12483 17289 12492 17323
rect 12440 17280 12492 17289
rect 13728 17280 13780 17332
rect 10784 17212 10836 17264
rect 4252 17144 4304 17196
rect 4712 17144 4764 17196
rect 5264 17144 5316 17196
rect 6460 17144 6512 17196
rect 6644 17144 6696 17196
rect 1676 17051 1728 17060
rect 1676 17017 1685 17051
rect 1685 17017 1719 17051
rect 1719 17017 1728 17051
rect 1676 17008 1728 17017
rect 2872 17076 2924 17128
rect 3884 17076 3936 17128
rect 2228 17008 2280 17060
rect 2412 17051 2464 17060
rect 2412 17017 2446 17051
rect 2446 17017 2464 17051
rect 2412 17008 2464 17017
rect 1768 16940 1820 16992
rect 4896 17076 4948 17128
rect 8024 17144 8076 17196
rect 7656 17076 7708 17128
rect 8852 17119 8904 17128
rect 8852 17085 8861 17119
rect 8861 17085 8895 17119
rect 8895 17085 8904 17119
rect 8852 17076 8904 17085
rect 9588 17144 9640 17196
rect 10968 17187 11020 17196
rect 10968 17153 10977 17187
rect 10977 17153 11011 17187
rect 11011 17153 11020 17187
rect 10968 17144 11020 17153
rect 12256 17212 12308 17264
rect 13452 17212 13504 17264
rect 16580 17280 16632 17332
rect 19064 17323 19116 17332
rect 19064 17289 19073 17323
rect 19073 17289 19107 17323
rect 19107 17289 19116 17323
rect 19064 17280 19116 17289
rect 19156 17280 19208 17332
rect 11612 17144 11664 17196
rect 12992 17144 13044 17196
rect 13636 17144 13688 17196
rect 16672 17212 16724 17264
rect 19340 17212 19392 17264
rect 19524 17212 19576 17264
rect 19708 17212 19760 17264
rect 11152 17076 11204 17128
rect 11796 17076 11848 17128
rect 12532 17076 12584 17128
rect 14096 17119 14148 17128
rect 14096 17085 14130 17119
rect 14130 17085 14148 17119
rect 14096 17076 14148 17085
rect 15292 17076 15344 17128
rect 4436 16940 4488 16992
rect 4712 16983 4764 16992
rect 4712 16949 4721 16983
rect 4721 16949 4755 16983
rect 4755 16949 4764 16983
rect 4712 16940 4764 16949
rect 5632 16940 5684 16992
rect 7472 17008 7524 17060
rect 8576 17008 8628 17060
rect 12716 17008 12768 17060
rect 12900 17008 12952 17060
rect 13728 17008 13780 17060
rect 14188 17008 14240 17060
rect 18880 17144 18932 17196
rect 20444 17144 20496 17196
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 16028 17008 16080 17060
rect 9680 16940 9732 16992
rect 10048 16940 10100 16992
rect 10508 16940 10560 16992
rect 12808 16983 12860 16992
rect 12808 16949 12817 16983
rect 12817 16949 12851 16983
rect 12851 16949 12860 16983
rect 12808 16940 12860 16949
rect 15936 16940 15988 16992
rect 16580 17076 16632 17128
rect 19064 17076 19116 17128
rect 19340 17076 19392 17128
rect 20536 17076 20588 17128
rect 19156 17008 19208 17060
rect 21640 17008 21692 17060
rect 17960 16940 18012 16992
rect 18420 16983 18472 16992
rect 18420 16949 18429 16983
rect 18429 16949 18463 16983
rect 18463 16949 18472 16983
rect 18420 16940 18472 16949
rect 19432 16983 19484 16992
rect 19432 16949 19441 16983
rect 19441 16949 19475 16983
rect 19475 16949 19484 16983
rect 19432 16940 19484 16949
rect 20628 16940 20680 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1768 16736 1820 16788
rect 2044 16779 2096 16788
rect 2044 16745 2053 16779
rect 2053 16745 2087 16779
rect 2087 16745 2096 16779
rect 2044 16736 2096 16745
rect 2596 16779 2648 16788
rect 2596 16745 2605 16779
rect 2605 16745 2639 16779
rect 2639 16745 2648 16779
rect 2596 16736 2648 16745
rect 4436 16779 4488 16788
rect 2780 16668 2832 16720
rect 3240 16668 3292 16720
rect 3976 16668 4028 16720
rect 4436 16745 4445 16779
rect 4445 16745 4479 16779
rect 4479 16745 4488 16779
rect 4436 16736 4488 16745
rect 4528 16736 4580 16788
rect 4344 16668 4396 16720
rect 6000 16668 6052 16720
rect 6828 16736 6880 16788
rect 7104 16736 7156 16788
rect 9588 16736 9640 16788
rect 11060 16736 11112 16788
rect 11980 16736 12032 16788
rect 15568 16736 15620 16788
rect 15660 16736 15712 16788
rect 16304 16779 16356 16788
rect 16304 16745 16313 16779
rect 16313 16745 16347 16779
rect 16347 16745 16356 16779
rect 16304 16736 16356 16745
rect 16396 16736 16448 16788
rect 18328 16779 18380 16788
rect 18328 16745 18337 16779
rect 18337 16745 18371 16779
rect 18371 16745 18380 16779
rect 18328 16736 18380 16745
rect 19616 16736 19668 16788
rect 20076 16736 20128 16788
rect 1860 16600 1912 16652
rect 3424 16600 3476 16652
rect 2412 16464 2464 16516
rect 3332 16532 3384 16584
rect 5172 16532 5224 16584
rect 5356 16600 5408 16652
rect 5540 16643 5592 16652
rect 5540 16609 5574 16643
rect 5574 16609 5592 16643
rect 5540 16600 5592 16609
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 8300 16668 8352 16720
rect 10968 16668 11020 16720
rect 12072 16668 12124 16720
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 10600 16600 10652 16652
rect 11888 16600 11940 16652
rect 11980 16600 12032 16652
rect 14372 16600 14424 16652
rect 14556 16600 14608 16652
rect 15476 16668 15528 16720
rect 18052 16668 18104 16720
rect 18972 16668 19024 16720
rect 19156 16668 19208 16720
rect 15660 16643 15712 16652
rect 7472 16575 7524 16584
rect 3884 16464 3936 16516
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 7472 16532 7524 16541
rect 7656 16532 7708 16584
rect 12900 16532 12952 16584
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 16488 16600 16540 16652
rect 16580 16600 16632 16652
rect 17776 16643 17828 16652
rect 17776 16609 17785 16643
rect 17785 16609 17819 16643
rect 17819 16609 17828 16643
rect 17776 16600 17828 16609
rect 16028 16532 16080 16584
rect 16764 16575 16816 16584
rect 16764 16541 16773 16575
rect 16773 16541 16807 16575
rect 16807 16541 16816 16575
rect 16764 16532 16816 16541
rect 6276 16464 6328 16516
rect 6920 16396 6972 16448
rect 8576 16396 8628 16448
rect 8852 16396 8904 16448
rect 11796 16396 11848 16448
rect 12992 16396 13044 16448
rect 14096 16396 14148 16448
rect 18604 16396 18656 16448
rect 20076 16600 20128 16652
rect 18788 16464 18840 16516
rect 19248 16532 19300 16584
rect 18972 16396 19024 16448
rect 20628 16396 20680 16448
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1492 16192 1544 16244
rect 4712 16192 4764 16244
rect 5356 16192 5408 16244
rect 6000 16235 6052 16244
rect 5448 16124 5500 16176
rect 6000 16201 6009 16235
rect 6009 16201 6043 16235
rect 6043 16201 6052 16235
rect 6000 16192 6052 16201
rect 7472 16192 7524 16244
rect 10140 16192 10192 16244
rect 10324 16192 10376 16244
rect 10508 16124 10560 16176
rect 3332 16099 3384 16108
rect 3332 16065 3341 16099
rect 3341 16065 3375 16099
rect 3375 16065 3384 16099
rect 3332 16056 3384 16065
rect 4252 16056 4304 16108
rect 5172 16056 5224 16108
rect 5632 16056 5684 16108
rect 1492 16031 1544 16040
rect 1492 15997 1501 16031
rect 1501 15997 1535 16031
rect 1535 15997 1544 16031
rect 1492 15988 1544 15997
rect 2136 15988 2188 16040
rect 2320 16031 2372 16040
rect 2320 15997 2329 16031
rect 2329 15997 2363 16031
rect 2363 15997 2372 16031
rect 2320 15988 2372 15997
rect 4160 16031 4212 16040
rect 4160 15997 4169 16031
rect 4169 15997 4203 16031
rect 4203 15997 4212 16031
rect 4160 15988 4212 15997
rect 6276 15988 6328 16040
rect 6460 15988 6512 16040
rect 6644 15988 6696 16040
rect 9588 16056 9640 16108
rect 12164 16192 12216 16244
rect 11796 16124 11848 16176
rect 13820 16192 13872 16244
rect 14372 16192 14424 16244
rect 15016 16192 15068 16244
rect 15660 16192 15712 16244
rect 16764 16192 16816 16244
rect 17592 16192 17644 16244
rect 13544 16124 13596 16176
rect 12992 16099 13044 16108
rect 8760 15988 8812 16040
rect 10600 15988 10652 16040
rect 11244 15988 11296 16040
rect 11336 15988 11388 16040
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 13268 16056 13320 16108
rect 14096 16099 14148 16108
rect 14096 16065 14105 16099
rect 14105 16065 14139 16099
rect 14139 16065 14148 16099
rect 14096 16056 14148 16065
rect 15200 16099 15252 16108
rect 15200 16065 15209 16099
rect 15209 16065 15243 16099
rect 15243 16065 15252 16099
rect 15200 16056 15252 16065
rect 15292 16056 15344 16108
rect 18788 16056 18840 16108
rect 19248 16124 19300 16176
rect 19340 16056 19392 16108
rect 20352 16056 20404 16108
rect 1400 15920 1452 15972
rect 4712 15920 4764 15972
rect 6920 15920 6972 15972
rect 8208 15920 8260 15972
rect 8392 15920 8444 15972
rect 11796 15920 11848 15972
rect 16396 15988 16448 16040
rect 16672 15988 16724 16040
rect 19248 15988 19300 16040
rect 19984 15988 20036 16040
rect 3240 15895 3292 15904
rect 3240 15861 3249 15895
rect 3249 15861 3283 15895
rect 3283 15861 3292 15895
rect 3240 15852 3292 15861
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 6736 15852 6788 15904
rect 6828 15852 6880 15904
rect 7656 15852 7708 15904
rect 8852 15895 8904 15904
rect 8852 15861 8861 15895
rect 8861 15861 8895 15895
rect 8895 15861 8904 15895
rect 8852 15852 8904 15861
rect 9680 15852 9732 15904
rect 10876 15852 10928 15904
rect 11888 15895 11940 15904
rect 11888 15861 11897 15895
rect 11897 15861 11931 15895
rect 11931 15861 11940 15895
rect 11888 15852 11940 15861
rect 12716 15852 12768 15904
rect 17960 15920 18012 15972
rect 15292 15852 15344 15904
rect 15752 15852 15804 15904
rect 16212 15852 16264 15904
rect 16856 15852 16908 15904
rect 17132 15852 17184 15904
rect 18144 15852 18196 15904
rect 18512 15852 18564 15904
rect 19340 15852 19392 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 2412 15648 2464 15700
rect 3516 15648 3568 15700
rect 4068 15648 4120 15700
rect 5724 15648 5776 15700
rect 6184 15648 6236 15700
rect 7196 15648 7248 15700
rect 7288 15648 7340 15700
rect 7656 15648 7708 15700
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 3240 15512 3292 15564
rect 6092 15580 6144 15632
rect 8852 15648 8904 15700
rect 12992 15648 13044 15700
rect 15292 15691 15344 15700
rect 8760 15580 8812 15632
rect 9220 15580 9272 15632
rect 1768 15444 1820 15496
rect 2596 15487 2648 15496
rect 2596 15453 2605 15487
rect 2605 15453 2639 15487
rect 2639 15453 2648 15487
rect 2596 15444 2648 15453
rect 3608 15487 3660 15496
rect 3608 15453 3617 15487
rect 3617 15453 3651 15487
rect 3651 15453 3660 15487
rect 3608 15444 3660 15453
rect 5540 15512 5592 15564
rect 5724 15555 5776 15564
rect 5724 15521 5733 15555
rect 5733 15521 5767 15555
rect 5767 15521 5776 15555
rect 5724 15512 5776 15521
rect 7564 15512 7616 15564
rect 4804 15487 4856 15496
rect 4160 15376 4212 15428
rect 4804 15453 4813 15487
rect 4813 15453 4847 15487
rect 4847 15453 4856 15487
rect 4804 15444 4856 15453
rect 5908 15487 5960 15496
rect 5908 15453 5917 15487
rect 5917 15453 5951 15487
rect 5951 15453 5960 15487
rect 5908 15444 5960 15453
rect 7104 15444 7156 15496
rect 7472 15444 7524 15496
rect 8576 15512 8628 15564
rect 8852 15512 8904 15564
rect 8208 15487 8260 15496
rect 8208 15453 8217 15487
rect 8217 15453 8251 15487
rect 8251 15453 8260 15487
rect 8208 15444 8260 15453
rect 9312 15444 9364 15496
rect 8484 15376 8536 15428
rect 11336 15580 11388 15632
rect 14096 15580 14148 15632
rect 15292 15657 15301 15691
rect 15301 15657 15335 15691
rect 15335 15657 15344 15691
rect 15292 15648 15344 15657
rect 18236 15648 18288 15700
rect 18328 15691 18380 15700
rect 18328 15657 18337 15691
rect 18337 15657 18371 15691
rect 18371 15657 18380 15691
rect 18328 15648 18380 15657
rect 18788 15648 18840 15700
rect 19340 15691 19392 15700
rect 17960 15580 18012 15632
rect 18052 15580 18104 15632
rect 10416 15555 10468 15564
rect 10416 15521 10425 15555
rect 10425 15521 10459 15555
rect 10459 15521 10468 15555
rect 10416 15512 10468 15521
rect 11244 15555 11296 15564
rect 11244 15521 11253 15555
rect 11253 15521 11287 15555
rect 11287 15521 11296 15555
rect 11244 15512 11296 15521
rect 11980 15512 12032 15564
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 10692 15487 10744 15496
rect 10692 15453 10701 15487
rect 10701 15453 10735 15487
rect 10735 15453 10744 15487
rect 10692 15444 10744 15453
rect 13544 15512 13596 15564
rect 14556 15512 14608 15564
rect 15016 15512 15068 15564
rect 15660 15555 15712 15564
rect 12900 15487 12952 15496
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 12900 15444 12952 15453
rect 13912 15444 13964 15496
rect 15660 15521 15669 15555
rect 15669 15521 15703 15555
rect 15703 15521 15712 15555
rect 15660 15512 15712 15521
rect 16672 15555 16724 15564
rect 16672 15521 16681 15555
rect 16681 15521 16715 15555
rect 16715 15521 16724 15555
rect 16672 15512 16724 15521
rect 17684 15555 17736 15564
rect 17684 15521 17693 15555
rect 17693 15521 17727 15555
rect 17727 15521 17736 15555
rect 17684 15512 17736 15521
rect 18328 15512 18380 15564
rect 18696 15623 18748 15632
rect 18696 15589 18705 15623
rect 18705 15589 18739 15623
rect 18739 15589 18748 15623
rect 18696 15580 18748 15589
rect 19340 15657 19349 15691
rect 19349 15657 19383 15691
rect 19383 15657 19392 15691
rect 19340 15648 19392 15657
rect 19800 15580 19852 15632
rect 15476 15444 15528 15496
rect 16028 15444 16080 15496
rect 16764 15487 16816 15496
rect 16764 15453 16773 15487
rect 16773 15453 16807 15487
rect 16807 15453 16816 15487
rect 16764 15444 16816 15453
rect 17868 15487 17920 15496
rect 17868 15453 17877 15487
rect 17877 15453 17911 15487
rect 17911 15453 17920 15487
rect 17868 15444 17920 15453
rect 4252 15351 4304 15360
rect 4252 15317 4261 15351
rect 4261 15317 4295 15351
rect 4295 15317 4304 15351
rect 4252 15308 4304 15317
rect 5172 15308 5224 15360
rect 6920 15308 6972 15360
rect 12164 15308 12216 15360
rect 14556 15308 14608 15360
rect 14648 15308 14700 15360
rect 17960 15308 18012 15360
rect 19248 15444 19300 15496
rect 20628 15444 20680 15496
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 3792 15104 3844 15156
rect 5724 15104 5776 15156
rect 6920 15104 6972 15156
rect 11796 15147 11848 15156
rect 6092 15036 6144 15088
rect 11796 15113 11805 15147
rect 11805 15113 11839 15147
rect 11839 15113 11848 15147
rect 11796 15104 11848 15113
rect 12808 15104 12860 15156
rect 17500 15104 17552 15156
rect 17868 15104 17920 15156
rect 7196 14968 7248 15020
rect 8116 14968 8168 15020
rect 13176 15036 13228 15088
rect 2044 14875 2096 14884
rect 2044 14841 2078 14875
rect 2078 14841 2096 14875
rect 2044 14832 2096 14841
rect 2228 14832 2280 14884
rect 4804 14900 4856 14952
rect 5080 14943 5132 14952
rect 5080 14909 5089 14943
rect 5089 14909 5123 14943
rect 5123 14909 5132 14943
rect 5080 14900 5132 14909
rect 5632 14900 5684 14952
rect 11888 14968 11940 15020
rect 5356 14875 5408 14884
rect 5356 14841 5390 14875
rect 5390 14841 5408 14875
rect 5356 14832 5408 14841
rect 9128 14832 9180 14884
rect 9588 14832 9640 14884
rect 10692 14875 10744 14884
rect 10692 14841 10726 14875
rect 10726 14841 10744 14875
rect 10692 14832 10744 14841
rect 13268 14900 13320 14952
rect 13912 14900 13964 14952
rect 12440 14832 12492 14884
rect 16028 14900 16080 14952
rect 18328 15036 18380 15088
rect 18420 14968 18472 15020
rect 19708 15011 19760 15020
rect 3516 14764 3568 14816
rect 5448 14764 5500 14816
rect 5908 14764 5960 14816
rect 6920 14764 6972 14816
rect 7472 14764 7524 14816
rect 7656 14764 7708 14816
rect 14556 14832 14608 14884
rect 15292 14832 15344 14884
rect 17960 14900 18012 14952
rect 17224 14832 17276 14884
rect 18512 14943 18564 14952
rect 18512 14909 18521 14943
rect 18521 14909 18555 14943
rect 18555 14909 18564 14943
rect 18512 14900 18564 14909
rect 11888 14764 11940 14816
rect 11980 14764 12032 14816
rect 12532 14764 12584 14816
rect 12808 14807 12860 14816
rect 12808 14773 12817 14807
rect 12817 14773 12851 14807
rect 12851 14773 12860 14807
rect 12808 14764 12860 14773
rect 13084 14764 13136 14816
rect 13636 14764 13688 14816
rect 15568 14807 15620 14816
rect 15568 14773 15577 14807
rect 15577 14773 15611 14807
rect 15611 14773 15620 14807
rect 15568 14764 15620 14773
rect 16212 14764 16264 14816
rect 17960 14764 18012 14816
rect 19432 14943 19484 14952
rect 19432 14909 19441 14943
rect 19441 14909 19475 14943
rect 19475 14909 19484 14943
rect 19432 14900 19484 14909
rect 19708 14977 19717 15011
rect 19717 14977 19751 15011
rect 19751 14977 19760 15011
rect 19708 14968 19760 14977
rect 20352 14968 20404 15020
rect 20812 14900 20864 14952
rect 19524 14807 19576 14816
rect 19524 14773 19533 14807
rect 19533 14773 19567 14807
rect 19567 14773 19576 14807
rect 19524 14764 19576 14773
rect 19984 14764 20036 14816
rect 20536 14807 20588 14816
rect 20536 14773 20545 14807
rect 20545 14773 20579 14807
rect 20579 14773 20588 14807
rect 20536 14764 20588 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 2872 14603 2924 14612
rect 2872 14569 2881 14603
rect 2881 14569 2915 14603
rect 2915 14569 2924 14603
rect 2872 14560 2924 14569
rect 4160 14560 4212 14612
rect 4252 14492 4304 14544
rect 5908 14560 5960 14612
rect 6368 14560 6420 14612
rect 8760 14560 8812 14612
rect 2044 14356 2096 14408
rect 3608 14424 3660 14476
rect 5632 14492 5684 14544
rect 6092 14492 6144 14544
rect 6552 14492 6604 14544
rect 8024 14492 8076 14544
rect 3516 14399 3568 14408
rect 3516 14365 3525 14399
rect 3525 14365 3559 14399
rect 3559 14365 3568 14399
rect 3516 14356 3568 14365
rect 7564 14424 7616 14476
rect 9588 14560 9640 14612
rect 10508 14560 10560 14612
rect 10968 14560 11020 14612
rect 13360 14560 13412 14612
rect 18420 14603 18472 14612
rect 9772 14492 9824 14544
rect 10692 14492 10744 14544
rect 14648 14492 14700 14544
rect 15108 14492 15160 14544
rect 16212 14492 16264 14544
rect 17868 14492 17920 14544
rect 18420 14569 18429 14603
rect 18429 14569 18463 14603
rect 18463 14569 18472 14603
rect 18420 14560 18472 14569
rect 18604 14560 18656 14612
rect 20536 14560 20588 14612
rect 18788 14492 18840 14544
rect 19248 14492 19300 14544
rect 19616 14492 19668 14544
rect 4804 14356 4856 14408
rect 5080 14288 5132 14340
rect 7380 14356 7432 14408
rect 9588 14424 9640 14476
rect 10048 14424 10100 14476
rect 11152 14424 11204 14476
rect 11336 14467 11388 14476
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 3608 14220 3660 14272
rect 4068 14220 4120 14272
rect 5448 14220 5500 14272
rect 7104 14288 7156 14340
rect 9312 14356 9364 14408
rect 9772 14356 9824 14408
rect 10048 14288 10100 14340
rect 10784 14356 10836 14408
rect 11060 14356 11112 14408
rect 11336 14433 11345 14467
rect 11345 14433 11379 14467
rect 11379 14433 11388 14467
rect 11336 14424 11388 14433
rect 13360 14467 13412 14476
rect 13360 14433 13369 14467
rect 13369 14433 13403 14467
rect 13403 14433 13412 14467
rect 13360 14424 13412 14433
rect 14372 14467 14424 14476
rect 14372 14433 14381 14467
rect 14381 14433 14415 14467
rect 14415 14433 14424 14467
rect 14372 14424 14424 14433
rect 15292 14467 15344 14476
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 11520 14399 11572 14408
rect 11520 14365 11529 14399
rect 11529 14365 11563 14399
rect 11563 14365 11572 14399
rect 11520 14356 11572 14365
rect 11888 14356 11940 14408
rect 12716 14356 12768 14408
rect 13544 14399 13596 14408
rect 13544 14365 13553 14399
rect 13553 14365 13587 14399
rect 13587 14365 13596 14399
rect 13544 14356 13596 14365
rect 14096 14356 14148 14408
rect 15292 14433 15301 14467
rect 15301 14433 15335 14467
rect 15335 14433 15344 14467
rect 15292 14424 15344 14433
rect 16028 14424 16080 14476
rect 17592 14424 17644 14476
rect 18696 14424 18748 14476
rect 16212 14356 16264 14408
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 6644 14220 6696 14272
rect 7380 14220 7432 14272
rect 7472 14220 7524 14272
rect 9128 14220 9180 14272
rect 13176 14288 13228 14340
rect 15936 14288 15988 14340
rect 16672 14288 16724 14340
rect 10600 14220 10652 14272
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 11980 14220 12032 14229
rect 13912 14220 13964 14272
rect 18052 14356 18104 14408
rect 18144 14288 18196 14340
rect 18788 14288 18840 14340
rect 17224 14220 17276 14272
rect 17408 14220 17460 14272
rect 19708 14356 19760 14408
rect 20720 14356 20772 14408
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 2872 13948 2924 14000
rect 3332 13948 3384 14000
rect 4160 14016 4212 14068
rect 5356 14059 5408 14068
rect 5356 14025 5365 14059
rect 5365 14025 5399 14059
rect 5399 14025 5408 14059
rect 5356 14016 5408 14025
rect 5540 14016 5592 14068
rect 6276 14016 6328 14068
rect 6644 14016 6696 14068
rect 7196 14016 7248 14068
rect 8116 14016 8168 14068
rect 9128 14016 9180 14068
rect 9864 14016 9916 14068
rect 10416 14016 10468 14068
rect 11152 14059 11204 14068
rect 11152 14025 11161 14059
rect 11161 14025 11195 14059
rect 11195 14025 11204 14059
rect 11152 14016 11204 14025
rect 14188 14016 14240 14068
rect 16764 14059 16816 14068
rect 1676 13812 1728 13864
rect 3700 13880 3752 13932
rect 1584 13744 1636 13796
rect 3884 13812 3936 13864
rect 5908 13880 5960 13932
rect 6736 13880 6788 13932
rect 8944 13948 8996 14000
rect 11888 13948 11940 14000
rect 16764 14025 16773 14059
rect 16773 14025 16807 14059
rect 16807 14025 16816 14059
rect 16764 14016 16816 14025
rect 18696 14016 18748 14068
rect 19616 14016 19668 14068
rect 20168 14016 20220 14068
rect 20904 14059 20956 14068
rect 20904 14025 20913 14059
rect 20913 14025 20947 14059
rect 20947 14025 20956 14059
rect 20904 14016 20956 14025
rect 7472 13880 7524 13932
rect 7656 13880 7708 13932
rect 10600 13923 10652 13932
rect 8116 13855 8168 13864
rect 8116 13821 8150 13855
rect 8150 13821 8168 13855
rect 8116 13812 8168 13821
rect 10600 13889 10609 13923
rect 10609 13889 10643 13923
rect 10643 13889 10652 13923
rect 10600 13880 10652 13889
rect 10784 13923 10836 13932
rect 10784 13889 10793 13923
rect 10793 13889 10827 13923
rect 10827 13889 10836 13923
rect 10784 13880 10836 13889
rect 11520 13880 11572 13932
rect 17408 13923 17460 13932
rect 11612 13855 11664 13864
rect 5448 13744 5500 13796
rect 5908 13744 5960 13796
rect 6368 13744 6420 13796
rect 7472 13744 7524 13796
rect 8300 13744 8352 13796
rect 9128 13744 9180 13796
rect 11612 13821 11621 13855
rect 11621 13821 11655 13855
rect 11655 13821 11664 13855
rect 11612 13812 11664 13821
rect 13544 13812 13596 13864
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 20076 13880 20128 13932
rect 10140 13744 10192 13796
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 2044 13676 2096 13728
rect 2964 13719 3016 13728
rect 2964 13685 2973 13719
rect 2973 13685 3007 13719
rect 3007 13685 3016 13719
rect 2964 13676 3016 13685
rect 7104 13676 7156 13728
rect 11060 13676 11112 13728
rect 11520 13719 11572 13728
rect 11520 13685 11529 13719
rect 11529 13685 11563 13719
rect 11563 13685 11572 13719
rect 11520 13676 11572 13685
rect 14096 13744 14148 13796
rect 14648 13744 14700 13796
rect 13820 13676 13872 13728
rect 15384 13855 15436 13864
rect 15384 13821 15418 13855
rect 15418 13821 15436 13855
rect 15384 13812 15436 13821
rect 17592 13812 17644 13864
rect 17960 13812 18012 13864
rect 18328 13855 18380 13864
rect 18328 13821 18362 13855
rect 18362 13821 18380 13855
rect 18328 13812 18380 13821
rect 15292 13744 15344 13796
rect 15936 13744 15988 13796
rect 18788 13744 18840 13796
rect 16212 13676 16264 13728
rect 16580 13676 16632 13728
rect 17224 13719 17276 13728
rect 17224 13685 17233 13719
rect 17233 13685 17267 13719
rect 17267 13685 17276 13719
rect 17224 13676 17276 13685
rect 17592 13676 17644 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 2044 13472 2096 13524
rect 3424 13472 3476 13524
rect 3700 13515 3752 13524
rect 3700 13481 3709 13515
rect 3709 13481 3743 13515
rect 3743 13481 3752 13515
rect 3700 13472 3752 13481
rect 4160 13515 4212 13524
rect 4160 13481 4169 13515
rect 4169 13481 4203 13515
rect 4203 13481 4212 13515
rect 4160 13472 4212 13481
rect 5632 13472 5684 13524
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 8208 13515 8260 13524
rect 8208 13481 8217 13515
rect 8217 13481 8251 13515
rect 8251 13481 8260 13515
rect 8208 13472 8260 13481
rect 9956 13472 10008 13524
rect 10508 13472 10560 13524
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 11152 13515 11204 13524
rect 11152 13481 11161 13515
rect 11161 13481 11195 13515
rect 11195 13481 11204 13515
rect 11152 13472 11204 13481
rect 11704 13515 11756 13524
rect 11704 13481 11713 13515
rect 11713 13481 11747 13515
rect 11747 13481 11756 13515
rect 11704 13472 11756 13481
rect 11980 13472 12032 13524
rect 12164 13515 12216 13524
rect 12164 13481 12173 13515
rect 12173 13481 12207 13515
rect 12207 13481 12216 13515
rect 12164 13472 12216 13481
rect 13452 13472 13504 13524
rect 15016 13472 15068 13524
rect 15752 13515 15804 13524
rect 2964 13404 3016 13456
rect 6736 13404 6788 13456
rect 7380 13404 7432 13456
rect 7840 13404 7892 13456
rect 2412 13336 2464 13388
rect 5448 13336 5500 13388
rect 2320 13311 2372 13320
rect 2320 13277 2329 13311
rect 2329 13277 2363 13311
rect 2363 13277 2372 13311
rect 2320 13268 2372 13277
rect 4068 13268 4120 13320
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 5724 13311 5776 13320
rect 5724 13277 5733 13311
rect 5733 13277 5767 13311
rect 5767 13277 5776 13311
rect 5724 13268 5776 13277
rect 7104 13336 7156 13388
rect 9588 13404 9640 13456
rect 10784 13404 10836 13456
rect 6552 13268 6604 13320
rect 6828 13268 6880 13320
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 8300 13311 8352 13320
rect 8300 13277 8309 13311
rect 8309 13277 8343 13311
rect 8343 13277 8352 13311
rect 8300 13268 8352 13277
rect 8668 13268 8720 13320
rect 9128 13336 9180 13388
rect 10232 13336 10284 13388
rect 10508 13268 10560 13320
rect 10692 13336 10744 13388
rect 12624 13404 12676 13456
rect 13728 13404 13780 13456
rect 15752 13481 15761 13515
rect 15761 13481 15795 13515
rect 15795 13481 15804 13515
rect 15752 13472 15804 13481
rect 16580 13472 16632 13524
rect 17224 13404 17276 13456
rect 17684 13472 17736 13524
rect 20720 13472 20772 13524
rect 18052 13404 18104 13456
rect 18144 13404 18196 13456
rect 11796 13336 11848 13388
rect 9956 13200 10008 13252
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 13544 13379 13596 13388
rect 12992 13336 13044 13345
rect 13544 13345 13553 13379
rect 13553 13345 13587 13379
rect 13587 13345 13596 13379
rect 13544 13336 13596 13345
rect 14188 13336 14240 13388
rect 14924 13336 14976 13388
rect 15200 13268 15252 13320
rect 16580 13336 16632 13388
rect 17040 13336 17092 13388
rect 18604 13447 18656 13456
rect 18604 13413 18613 13447
rect 18613 13413 18647 13447
rect 18647 13413 18656 13447
rect 18604 13404 18656 13413
rect 18788 13404 18840 13456
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 16764 13268 16816 13320
rect 17408 13268 17460 13320
rect 11796 13200 11848 13252
rect 13268 13200 13320 13252
rect 13544 13200 13596 13252
rect 5080 13132 5132 13184
rect 5908 13132 5960 13184
rect 6736 13175 6788 13184
rect 6736 13141 6745 13175
rect 6745 13141 6779 13175
rect 6779 13141 6788 13175
rect 6736 13132 6788 13141
rect 7012 13132 7064 13184
rect 7748 13132 7800 13184
rect 8208 13132 8260 13184
rect 8576 13132 8628 13184
rect 9312 13132 9364 13184
rect 12348 13132 12400 13184
rect 18420 13200 18472 13252
rect 18972 13268 19024 13320
rect 20168 13268 20220 13320
rect 15384 13132 15436 13184
rect 15936 13132 15988 13184
rect 17224 13132 17276 13184
rect 17500 13132 17552 13184
rect 18696 13132 18748 13184
rect 19708 13132 19760 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 5448 12971 5500 12980
rect 5448 12937 5457 12971
rect 5457 12937 5491 12971
rect 5491 12937 5500 12971
rect 5448 12928 5500 12937
rect 6460 12971 6512 12980
rect 6460 12937 6469 12971
rect 6469 12937 6503 12971
rect 6503 12937 6512 12971
rect 6460 12928 6512 12937
rect 4068 12860 4120 12912
rect 2412 12792 2464 12844
rect 2320 12724 2372 12776
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 3884 12724 3936 12776
rect 4436 12724 4488 12776
rect 3516 12656 3568 12708
rect 5724 12792 5776 12844
rect 6644 12860 6696 12912
rect 8300 12928 8352 12980
rect 8668 12903 8720 12912
rect 8668 12869 8677 12903
rect 8677 12869 8711 12903
rect 8711 12869 8720 12903
rect 8668 12860 8720 12869
rect 4896 12724 4948 12776
rect 6368 12724 6420 12776
rect 5448 12656 5500 12708
rect 6276 12656 6328 12708
rect 2964 12588 3016 12640
rect 5908 12631 5960 12640
rect 5908 12597 5917 12631
rect 5917 12597 5951 12631
rect 5951 12597 5960 12631
rect 6828 12656 6880 12708
rect 7840 12724 7892 12776
rect 9312 12767 9364 12776
rect 9312 12733 9321 12767
rect 9321 12733 9355 12767
rect 9355 12733 9364 12767
rect 9312 12724 9364 12733
rect 11428 12860 11480 12912
rect 14096 12903 14148 12912
rect 14096 12869 14105 12903
rect 14105 12869 14139 12903
rect 14139 12869 14148 12903
rect 14096 12860 14148 12869
rect 14464 12928 14516 12980
rect 16488 12928 16540 12980
rect 16672 12928 16724 12980
rect 18788 12928 18840 12980
rect 20444 12928 20496 12980
rect 17684 12860 17736 12912
rect 10232 12792 10284 12844
rect 10508 12835 10560 12844
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 10784 12792 10836 12844
rect 14556 12792 14608 12844
rect 10968 12724 11020 12776
rect 11152 12724 11204 12776
rect 12072 12724 12124 12776
rect 12440 12724 12492 12776
rect 13912 12724 13964 12776
rect 16396 12792 16448 12844
rect 16764 12835 16816 12844
rect 5908 12588 5960 12597
rect 7380 12588 7432 12640
rect 8944 12631 8996 12640
rect 8944 12597 8953 12631
rect 8953 12597 8987 12631
rect 8987 12597 8996 12631
rect 8944 12588 8996 12597
rect 9864 12588 9916 12640
rect 10232 12588 10284 12640
rect 10416 12588 10468 12640
rect 13176 12656 13228 12708
rect 15660 12767 15712 12776
rect 15660 12733 15669 12767
rect 15669 12733 15703 12767
rect 15703 12733 15712 12767
rect 15660 12724 15712 12733
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 19156 12860 19208 12912
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 17224 12767 17276 12776
rect 17224 12733 17233 12767
rect 17233 12733 17267 12767
rect 17267 12733 17276 12767
rect 17224 12724 17276 12733
rect 18512 12724 18564 12776
rect 18880 12724 18932 12776
rect 11336 12631 11388 12640
rect 11336 12597 11345 12631
rect 11345 12597 11379 12631
rect 11379 12597 11388 12631
rect 11336 12588 11388 12597
rect 13268 12588 13320 12640
rect 15200 12588 15252 12640
rect 17040 12656 17092 12708
rect 17500 12699 17552 12708
rect 17500 12665 17509 12699
rect 17509 12665 17543 12699
rect 17543 12665 17552 12699
rect 17500 12656 17552 12665
rect 17684 12656 17736 12708
rect 20168 12860 20220 12912
rect 20720 12860 20772 12912
rect 19432 12792 19484 12844
rect 19708 12767 19760 12776
rect 19708 12733 19717 12767
rect 19717 12733 19751 12767
rect 19751 12733 19760 12767
rect 19708 12724 19760 12733
rect 19800 12767 19852 12776
rect 19800 12733 19809 12767
rect 19809 12733 19843 12767
rect 19843 12733 19852 12767
rect 19800 12724 19852 12733
rect 16304 12588 16356 12640
rect 18144 12588 18196 12640
rect 18420 12588 18472 12640
rect 19156 12588 19208 12640
rect 20168 12588 20220 12640
rect 20812 12631 20864 12640
rect 20812 12597 20821 12631
rect 20821 12597 20855 12631
rect 20855 12597 20864 12631
rect 20812 12588 20864 12597
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2780 12384 2832 12436
rect 2964 12427 3016 12436
rect 2964 12393 2973 12427
rect 2973 12393 3007 12427
rect 3007 12393 3016 12427
rect 2964 12384 3016 12393
rect 3976 12384 4028 12436
rect 5724 12384 5776 12436
rect 6368 12384 6420 12436
rect 6644 12384 6696 12436
rect 7564 12384 7616 12436
rect 1492 12316 1544 12368
rect 7932 12316 7984 12368
rect 10232 12384 10284 12436
rect 11888 12427 11940 12436
rect 11888 12393 11897 12427
rect 11897 12393 11931 12427
rect 11931 12393 11940 12427
rect 11888 12384 11940 12393
rect 12164 12384 12216 12436
rect 12716 12427 12768 12436
rect 12716 12393 12725 12427
rect 12725 12393 12759 12427
rect 12759 12393 12768 12427
rect 12716 12384 12768 12393
rect 13268 12384 13320 12436
rect 13360 12384 13412 12436
rect 15476 12384 15528 12436
rect 15660 12384 15712 12436
rect 1768 12248 1820 12300
rect 2964 12248 3016 12300
rect 3332 12291 3384 12300
rect 3332 12257 3341 12291
rect 3341 12257 3375 12291
rect 3375 12257 3384 12291
rect 3332 12248 3384 12257
rect 4436 12248 4488 12300
rect 4988 12291 5040 12300
rect 4988 12257 5022 12291
rect 5022 12257 5040 12291
rect 4988 12248 5040 12257
rect 7656 12248 7708 12300
rect 8576 12248 8628 12300
rect 9864 12291 9916 12300
rect 9864 12257 9873 12291
rect 9873 12257 9907 12291
rect 9907 12257 9916 12291
rect 9864 12248 9916 12257
rect 9956 12248 10008 12300
rect 10876 12248 10928 12300
rect 1952 12180 2004 12232
rect 2136 12180 2188 12232
rect 2780 12180 2832 12232
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 3516 12223 3568 12232
rect 3516 12189 3525 12223
rect 3525 12189 3559 12223
rect 3559 12189 3568 12223
rect 3516 12180 3568 12189
rect 6184 12180 6236 12232
rect 6828 12223 6880 12232
rect 6828 12189 6837 12223
rect 6837 12189 6871 12223
rect 6871 12189 6880 12223
rect 6828 12180 6880 12189
rect 3240 12112 3292 12164
rect 5908 12112 5960 12164
rect 6552 12112 6604 12164
rect 7840 12223 7892 12232
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 11336 12223 11388 12232
rect 2136 12044 2188 12096
rect 6460 12044 6512 12096
rect 7104 12044 7156 12096
rect 8116 12112 8168 12164
rect 8668 12112 8720 12164
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 11336 12180 11388 12189
rect 11428 12180 11480 12232
rect 12532 12180 12584 12232
rect 9680 12112 9732 12164
rect 9864 12112 9916 12164
rect 10876 12112 10928 12164
rect 14004 12248 14056 12300
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 13728 12180 13780 12232
rect 14464 12180 14516 12232
rect 16580 12384 16632 12436
rect 17592 12384 17644 12436
rect 17224 12316 17276 12368
rect 19340 12384 19392 12436
rect 19616 12384 19668 12436
rect 19892 12384 19944 12436
rect 20076 12384 20128 12436
rect 21456 12384 21508 12436
rect 18512 12316 18564 12368
rect 18788 12316 18840 12368
rect 19064 12316 19116 12368
rect 19248 12316 19300 12368
rect 15844 12112 15896 12164
rect 18052 12248 18104 12300
rect 20444 12248 20496 12300
rect 9220 12044 9272 12096
rect 9588 12044 9640 12096
rect 10232 12044 10284 12096
rect 13176 12044 13228 12096
rect 14740 12044 14792 12096
rect 15200 12044 15252 12096
rect 16396 12044 16448 12096
rect 19800 12180 19852 12232
rect 18880 12044 18932 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 5632 11840 5684 11892
rect 6276 11840 6328 11892
rect 7840 11883 7892 11892
rect 7840 11849 7849 11883
rect 7849 11849 7883 11883
rect 7883 11849 7892 11883
rect 7840 11840 7892 11849
rect 7932 11840 7984 11892
rect 4620 11772 4672 11824
rect 4896 11772 4948 11824
rect 3240 11704 3292 11756
rect 6552 11772 6604 11824
rect 7748 11772 7800 11824
rect 8668 11772 8720 11824
rect 1400 11568 1452 11620
rect 2596 11636 2648 11688
rect 4252 11568 4304 11620
rect 4620 11568 4672 11620
rect 2320 11500 2372 11552
rect 4068 11500 4120 11552
rect 4988 11636 5040 11688
rect 5908 11679 5960 11688
rect 5908 11645 5917 11679
rect 5917 11645 5951 11679
rect 5951 11645 5960 11679
rect 5908 11636 5960 11645
rect 6736 11636 6788 11688
rect 8760 11704 8812 11756
rect 9220 11772 9272 11824
rect 8208 11679 8260 11688
rect 8208 11645 8217 11679
rect 8217 11645 8251 11679
rect 8251 11645 8260 11679
rect 8208 11636 8260 11645
rect 8944 11636 8996 11688
rect 9588 11840 9640 11892
rect 9680 11840 9732 11892
rect 12164 11840 12216 11892
rect 13544 11840 13596 11892
rect 14740 11840 14792 11892
rect 16028 11840 16080 11892
rect 16212 11840 16264 11892
rect 9588 11704 9640 11756
rect 9956 11704 10008 11756
rect 11888 11772 11940 11824
rect 14372 11772 14424 11824
rect 17776 11772 17828 11824
rect 11796 11704 11848 11756
rect 9496 11636 9548 11688
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12440 11636 12492 11645
rect 15568 11704 15620 11756
rect 16212 11704 16264 11756
rect 17316 11704 17368 11756
rect 18604 11840 18656 11892
rect 20996 11883 21048 11892
rect 20996 11849 21005 11883
rect 21005 11849 21039 11883
rect 21039 11849 21048 11883
rect 20996 11840 21048 11849
rect 19248 11772 19300 11824
rect 21088 11772 21140 11824
rect 14188 11636 14240 11688
rect 6092 11568 6144 11620
rect 6368 11568 6420 11620
rect 7012 11568 7064 11620
rect 8668 11568 8720 11620
rect 10692 11568 10744 11620
rect 10876 11611 10928 11620
rect 10876 11577 10910 11611
rect 10910 11577 10928 11611
rect 10876 11568 10928 11577
rect 11888 11568 11940 11620
rect 9404 11500 9456 11552
rect 9588 11500 9640 11552
rect 9956 11500 10008 11552
rect 11980 11500 12032 11552
rect 12072 11500 12124 11552
rect 15200 11636 15252 11688
rect 16396 11636 16448 11688
rect 16580 11679 16632 11688
rect 16580 11645 16614 11679
rect 16614 11645 16632 11679
rect 16580 11636 16632 11645
rect 16948 11636 17000 11688
rect 17776 11636 17828 11688
rect 17960 11636 18012 11688
rect 18972 11704 19024 11756
rect 19432 11704 19484 11756
rect 20168 11679 20220 11688
rect 20168 11645 20177 11679
rect 20177 11645 20211 11679
rect 20211 11645 20220 11679
rect 20168 11636 20220 11645
rect 20996 11636 21048 11688
rect 15568 11568 15620 11620
rect 15384 11500 15436 11552
rect 19616 11568 19668 11620
rect 17132 11500 17184 11552
rect 18972 11500 19024 11552
rect 19156 11543 19208 11552
rect 19156 11509 19165 11543
rect 19165 11509 19199 11543
rect 19199 11509 19208 11543
rect 19156 11500 19208 11509
rect 19432 11500 19484 11552
rect 20720 11500 20772 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 1492 11296 1544 11348
rect 3240 11339 3292 11348
rect 3240 11305 3249 11339
rect 3249 11305 3283 11339
rect 3283 11305 3292 11339
rect 3240 11296 3292 11305
rect 3332 11296 3384 11348
rect 4068 11339 4120 11348
rect 4068 11305 4077 11339
rect 4077 11305 4111 11339
rect 4111 11305 4120 11339
rect 4068 11296 4120 11305
rect 2596 11228 2648 11280
rect 3884 11228 3936 11280
rect 5816 11296 5868 11348
rect 6276 11296 6328 11348
rect 7104 11296 7156 11348
rect 6736 11228 6788 11280
rect 6828 11228 6880 11280
rect 2688 11160 2740 11212
rect 4160 11160 4212 11212
rect 5080 11203 5132 11212
rect 5080 11169 5089 11203
rect 5089 11169 5123 11203
rect 5123 11169 5132 11203
rect 5080 11160 5132 11169
rect 6920 11160 6972 11212
rect 7748 11203 7800 11212
rect 7748 11169 7782 11203
rect 7782 11169 7800 11203
rect 8116 11228 8168 11280
rect 8392 11228 8444 11280
rect 8760 11296 8812 11348
rect 9036 11296 9088 11348
rect 9680 11296 9732 11348
rect 10232 11296 10284 11348
rect 10692 11296 10744 11348
rect 11704 11296 11756 11348
rect 12072 11296 12124 11348
rect 7748 11160 7800 11169
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 10416 11228 10468 11280
rect 11520 11228 11572 11280
rect 9956 11160 10008 11169
rect 12164 11160 12216 11212
rect 15384 11228 15436 11280
rect 4252 11092 4304 11144
rect 3240 11024 3292 11076
rect 5632 11092 5684 11144
rect 7012 11092 7064 11144
rect 4712 11024 4764 11076
rect 5724 11024 5776 11076
rect 11980 11092 12032 11144
rect 13728 11160 13780 11212
rect 14004 11160 14056 11212
rect 14556 11203 14608 11212
rect 14556 11169 14565 11203
rect 14565 11169 14599 11203
rect 14599 11169 14608 11203
rect 15844 11296 15896 11348
rect 18420 11296 18472 11348
rect 16856 11228 16908 11280
rect 14556 11160 14608 11169
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 12440 11092 12492 11101
rect 4068 10956 4120 11008
rect 11520 11024 11572 11076
rect 11796 11024 11848 11076
rect 12072 11024 12124 11076
rect 16396 11092 16448 11144
rect 12624 10956 12676 11008
rect 12808 10956 12860 11008
rect 13912 11024 13964 11076
rect 17776 11228 17828 11280
rect 17224 11160 17276 11212
rect 19156 11296 19208 11348
rect 19248 11228 19300 11280
rect 20352 11228 20404 11280
rect 17132 11135 17184 11144
rect 17132 11101 17141 11135
rect 17141 11101 17175 11135
rect 17175 11101 17184 11135
rect 17132 11092 17184 11101
rect 18788 11092 18840 11144
rect 17316 11024 17368 11076
rect 17960 11024 18012 11076
rect 14096 10999 14148 11008
rect 14096 10965 14105 10999
rect 14105 10965 14139 10999
rect 14139 10965 14148 10999
rect 14096 10956 14148 10965
rect 14188 10956 14240 11008
rect 16672 10956 16724 11008
rect 18696 11024 18748 11076
rect 20628 11160 20680 11212
rect 19800 10956 19852 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 1768 10752 1820 10804
rect 3240 10795 3292 10804
rect 3240 10761 3249 10795
rect 3249 10761 3283 10795
rect 3283 10761 3292 10795
rect 3240 10752 3292 10761
rect 3792 10752 3844 10804
rect 4252 10752 4304 10804
rect 4344 10684 4396 10736
rect 6736 10752 6788 10804
rect 7380 10752 7432 10804
rect 8576 10752 8628 10804
rect 8944 10752 8996 10804
rect 11796 10752 11848 10804
rect 11980 10752 12032 10804
rect 12992 10752 13044 10804
rect 5264 10684 5316 10736
rect 3240 10548 3292 10600
rect 5448 10616 5500 10668
rect 5908 10659 5960 10668
rect 5908 10625 5917 10659
rect 5917 10625 5951 10659
rect 5951 10625 5960 10659
rect 5908 10616 5960 10625
rect 8116 10684 8168 10736
rect 9312 10727 9364 10736
rect 9312 10693 9321 10727
rect 9321 10693 9355 10727
rect 9355 10693 9364 10727
rect 9312 10684 9364 10693
rect 10784 10684 10836 10736
rect 11336 10684 11388 10736
rect 12532 10684 12584 10736
rect 13176 10684 13228 10736
rect 13452 10727 13504 10736
rect 13452 10693 13461 10727
rect 13461 10693 13495 10727
rect 13495 10693 13504 10727
rect 13452 10684 13504 10693
rect 14372 10752 14424 10804
rect 16028 10752 16080 10804
rect 17224 10752 17276 10804
rect 6368 10616 6420 10668
rect 6828 10548 6880 10600
rect 7564 10616 7616 10668
rect 8208 10548 8260 10600
rect 11244 10616 11296 10668
rect 13728 10616 13780 10668
rect 13912 10659 13964 10668
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 19156 10752 19208 10804
rect 21180 10752 21232 10804
rect 15384 10659 15436 10668
rect 8944 10548 8996 10600
rect 9496 10548 9548 10600
rect 9588 10548 9640 10600
rect 2596 10480 2648 10532
rect 2780 10480 2832 10532
rect 3976 10480 4028 10532
rect 3332 10412 3384 10464
rect 5724 10480 5776 10532
rect 6736 10480 6788 10532
rect 7288 10523 7340 10532
rect 7288 10489 7297 10523
rect 7297 10489 7331 10523
rect 7331 10489 7340 10523
rect 7288 10480 7340 10489
rect 7564 10480 7616 10532
rect 8392 10480 8444 10532
rect 8760 10480 8812 10532
rect 10876 10548 10928 10600
rect 11060 10548 11112 10600
rect 11612 10591 11664 10600
rect 11612 10557 11621 10591
rect 11621 10557 11655 10591
rect 11655 10557 11664 10591
rect 11980 10591 12032 10600
rect 11612 10548 11664 10557
rect 11980 10557 11989 10591
rect 11989 10557 12023 10591
rect 12023 10557 12032 10591
rect 11980 10548 12032 10557
rect 12348 10548 12400 10600
rect 11244 10480 11296 10532
rect 11704 10480 11756 10532
rect 6092 10412 6144 10464
rect 6920 10412 6972 10464
rect 7748 10412 7800 10464
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 10324 10412 10376 10464
rect 11060 10412 11112 10464
rect 12716 10412 12768 10464
rect 13176 10412 13228 10464
rect 14096 10548 14148 10600
rect 14188 10548 14240 10600
rect 15384 10625 15393 10659
rect 15393 10625 15427 10659
rect 15427 10625 15436 10659
rect 15384 10616 15436 10625
rect 15568 10616 15620 10668
rect 16488 10616 16540 10668
rect 16856 10616 16908 10668
rect 17132 10616 17184 10668
rect 20168 10616 20220 10668
rect 20628 10616 20680 10668
rect 16948 10548 17000 10600
rect 13912 10480 13964 10532
rect 14556 10412 14608 10464
rect 14924 10480 14976 10532
rect 18052 10480 18104 10532
rect 18880 10548 18932 10600
rect 18972 10548 19024 10600
rect 20536 10548 20588 10600
rect 20904 10548 20956 10600
rect 18236 10480 18288 10532
rect 18696 10480 18748 10532
rect 18788 10480 18840 10532
rect 17224 10412 17276 10464
rect 17316 10412 17368 10464
rect 17592 10412 17644 10464
rect 19800 10455 19852 10464
rect 19800 10421 19809 10455
rect 19809 10421 19843 10455
rect 19843 10421 19852 10455
rect 19800 10412 19852 10421
rect 20076 10412 20128 10464
rect 21916 10412 21968 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 1676 10251 1728 10260
rect 1676 10217 1685 10251
rect 1685 10217 1719 10251
rect 1719 10217 1728 10251
rect 1676 10208 1728 10217
rect 2872 10208 2924 10260
rect 2780 10140 2832 10192
rect 6368 10208 6420 10260
rect 7748 10208 7800 10260
rect 8668 10208 8720 10260
rect 8852 10208 8904 10260
rect 9220 10251 9272 10260
rect 9220 10217 9229 10251
rect 9229 10217 9263 10251
rect 9263 10217 9272 10251
rect 9220 10208 9272 10217
rect 9496 10208 9548 10260
rect 11336 10208 11388 10260
rect 11704 10208 11756 10260
rect 12440 10208 12492 10260
rect 1860 10072 1912 10124
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 4252 10140 4304 10192
rect 12624 10140 12676 10192
rect 3240 10072 3292 10124
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 5632 10072 5684 10124
rect 5908 10072 5960 10124
rect 7380 10072 7432 10124
rect 8116 10115 8168 10124
rect 8116 10081 8125 10115
rect 8125 10081 8159 10115
rect 8159 10081 8168 10115
rect 8116 10072 8168 10081
rect 8576 10072 8628 10124
rect 9036 10115 9088 10124
rect 9036 10081 9045 10115
rect 9045 10081 9079 10115
rect 9079 10081 9088 10115
rect 9036 10072 9088 10081
rect 9404 10072 9456 10124
rect 9588 10072 9640 10124
rect 9772 10072 9824 10124
rect 10784 10072 10836 10124
rect 11704 10072 11756 10124
rect 12256 10072 12308 10124
rect 12348 10072 12400 10124
rect 13544 10208 13596 10260
rect 15568 10208 15620 10260
rect 15752 10208 15804 10260
rect 17684 10208 17736 10260
rect 18144 10208 18196 10260
rect 20076 10208 20128 10260
rect 20352 10208 20404 10260
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 6184 10047 6236 10056
rect 6184 10013 6193 10047
rect 6193 10013 6227 10047
rect 6227 10013 6236 10047
rect 6184 10004 6236 10013
rect 5264 9936 5316 9988
rect 2320 9868 2372 9920
rect 5448 9911 5500 9920
rect 5448 9877 5457 9911
rect 5457 9877 5491 9911
rect 5491 9877 5500 9911
rect 5448 9868 5500 9877
rect 5540 9868 5592 9920
rect 5908 9868 5960 9920
rect 6552 10004 6604 10056
rect 6920 10004 6972 10056
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 7288 9936 7340 9988
rect 10876 10004 10928 10056
rect 9680 9936 9732 9988
rect 6552 9911 6604 9920
rect 6552 9877 6561 9911
rect 6561 9877 6595 9911
rect 6595 9877 6604 9911
rect 6552 9868 6604 9877
rect 7380 9868 7432 9920
rect 7748 9911 7800 9920
rect 7748 9877 7757 9911
rect 7757 9877 7791 9911
rect 7791 9877 7800 9911
rect 7748 9868 7800 9877
rect 8576 9868 8628 9920
rect 9312 9868 9364 9920
rect 11520 9936 11572 9988
rect 11152 9868 11204 9920
rect 12072 9868 12124 9920
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12992 9936 13044 9988
rect 14280 10072 14332 10124
rect 14556 10072 14608 10124
rect 15384 10072 15436 10124
rect 17408 10072 17460 10124
rect 17592 10072 17644 10124
rect 15108 10004 15160 10056
rect 15200 10004 15252 10056
rect 16488 10004 16540 10056
rect 16856 10004 16908 10056
rect 16948 10004 17000 10056
rect 18144 10072 18196 10124
rect 18696 10140 18748 10192
rect 18788 10140 18840 10192
rect 20260 10140 20312 10192
rect 20720 10140 20772 10192
rect 19156 10072 19208 10124
rect 19340 10115 19392 10124
rect 19340 10081 19374 10115
rect 19374 10081 19392 10115
rect 19340 10072 19392 10081
rect 18788 10004 18840 10056
rect 20904 10047 20956 10056
rect 20904 10013 20913 10047
rect 20913 10013 20947 10047
rect 20947 10013 20956 10047
rect 20904 10004 20956 10013
rect 12440 9868 12492 9877
rect 13728 9868 13780 9920
rect 14096 9868 14148 9920
rect 14372 9868 14424 9920
rect 16488 9868 16540 9920
rect 17132 9868 17184 9920
rect 17776 9936 17828 9988
rect 18972 9868 19024 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 2504 9664 2556 9716
rect 5724 9664 5776 9716
rect 8760 9664 8812 9716
rect 9404 9664 9456 9716
rect 9772 9664 9824 9716
rect 10416 9664 10468 9716
rect 12348 9664 12400 9716
rect 13084 9664 13136 9716
rect 17592 9707 17644 9716
rect 3056 9596 3108 9648
rect 3516 9596 3568 9648
rect 3792 9596 3844 9648
rect 4160 9639 4212 9648
rect 4160 9605 4169 9639
rect 4169 9605 4203 9639
rect 4203 9605 4212 9639
rect 4160 9596 4212 9605
rect 5264 9596 5316 9648
rect 6368 9639 6420 9648
rect 2412 9528 2464 9580
rect 1860 9460 1912 9512
rect 3240 9528 3292 9580
rect 4252 9528 4304 9580
rect 5448 9528 5500 9580
rect 6368 9605 6377 9639
rect 6377 9605 6411 9639
rect 6411 9605 6420 9639
rect 6368 9596 6420 9605
rect 6828 9639 6880 9648
rect 6828 9605 6837 9639
rect 6837 9605 6871 9639
rect 6871 9605 6880 9639
rect 6828 9596 6880 9605
rect 7196 9596 7248 9648
rect 7656 9596 7708 9648
rect 9680 9596 9732 9648
rect 10876 9596 10928 9648
rect 7564 9528 7616 9580
rect 5540 9460 5592 9512
rect 8944 9528 8996 9580
rect 10232 9528 10284 9580
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 13820 9596 13872 9648
rect 2596 9435 2648 9444
rect 2596 9401 2605 9435
rect 2605 9401 2639 9435
rect 2639 9401 2648 9435
rect 2596 9392 2648 9401
rect 2412 9324 2464 9376
rect 2504 9367 2556 9376
rect 2504 9333 2513 9367
rect 2513 9333 2547 9367
rect 2547 9333 2556 9367
rect 2504 9324 2556 9333
rect 2964 9324 3016 9376
rect 3884 9392 3936 9444
rect 3700 9324 3752 9376
rect 5724 9392 5776 9444
rect 9496 9460 9548 9512
rect 7932 9392 7984 9444
rect 8760 9392 8812 9444
rect 8852 9392 8904 9444
rect 5264 9324 5316 9376
rect 5632 9367 5684 9376
rect 5632 9333 5641 9367
rect 5641 9333 5675 9367
rect 5675 9333 5684 9367
rect 5632 9324 5684 9333
rect 5908 9324 5960 9376
rect 9312 9324 9364 9376
rect 9496 9367 9548 9376
rect 9496 9333 9505 9367
rect 9505 9333 9539 9367
rect 9539 9333 9548 9367
rect 9496 9324 9548 9333
rect 9956 9367 10008 9376
rect 9956 9333 9965 9367
rect 9965 9333 9999 9367
rect 9999 9333 10008 9367
rect 9956 9324 10008 9333
rect 10968 9435 11020 9444
rect 10968 9401 10977 9435
rect 10977 9401 11011 9435
rect 11011 9401 11020 9435
rect 10968 9392 11020 9401
rect 11520 9392 11572 9444
rect 11704 9435 11756 9444
rect 11704 9401 11713 9435
rect 11713 9401 11747 9435
rect 11747 9401 11756 9435
rect 11704 9392 11756 9401
rect 11796 9435 11848 9444
rect 11796 9401 11805 9435
rect 11805 9401 11839 9435
rect 11839 9401 11848 9435
rect 12348 9460 12400 9512
rect 12532 9460 12584 9512
rect 14096 9460 14148 9512
rect 14464 9596 14516 9648
rect 14924 9571 14976 9580
rect 14372 9460 14424 9512
rect 14924 9537 14933 9571
rect 14933 9537 14967 9571
rect 14967 9537 14976 9571
rect 14924 9528 14976 9537
rect 15200 9596 15252 9648
rect 15752 9596 15804 9648
rect 17592 9673 17601 9707
rect 17601 9673 17635 9707
rect 17635 9673 17644 9707
rect 17592 9664 17644 9673
rect 17960 9664 18012 9716
rect 17132 9639 17184 9648
rect 17132 9605 17141 9639
rect 17141 9605 17175 9639
rect 17175 9605 17184 9639
rect 17132 9596 17184 9605
rect 20720 9664 20772 9716
rect 19064 9639 19116 9648
rect 19064 9605 19073 9639
rect 19073 9605 19107 9639
rect 19107 9605 19116 9639
rect 19064 9596 19116 9605
rect 19248 9596 19300 9648
rect 11796 9392 11848 9401
rect 12808 9392 12860 9444
rect 15568 9460 15620 9512
rect 15752 9503 15804 9512
rect 15752 9469 15761 9503
rect 15761 9469 15795 9503
rect 15795 9469 15804 9503
rect 15752 9460 15804 9469
rect 17776 9528 17828 9580
rect 17868 9528 17920 9580
rect 17500 9460 17552 9512
rect 19616 9528 19668 9580
rect 19708 9571 19760 9580
rect 19708 9537 19717 9571
rect 19717 9537 19751 9571
rect 19751 9537 19760 9571
rect 19708 9528 19760 9537
rect 19156 9460 19208 9512
rect 10692 9324 10744 9376
rect 11980 9324 12032 9376
rect 15292 9392 15344 9444
rect 16488 9392 16540 9444
rect 16672 9392 16724 9444
rect 17592 9392 17644 9444
rect 12992 9324 13044 9376
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 16304 9324 16356 9376
rect 19248 9392 19300 9444
rect 19616 9392 19668 9444
rect 19800 9460 19852 9512
rect 20904 9392 20956 9444
rect 19432 9324 19484 9376
rect 19708 9324 19760 9376
rect 19800 9324 19852 9376
rect 20536 9367 20588 9376
rect 20536 9333 20545 9367
rect 20545 9333 20579 9367
rect 20579 9333 20588 9367
rect 20536 9324 20588 9333
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2228 9120 2280 9172
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 2596 9120 2648 9172
rect 4712 9120 4764 9172
rect 2320 9095 2372 9104
rect 2320 9061 2329 9095
rect 2329 9061 2363 9095
rect 2363 9061 2372 9095
rect 2320 9052 2372 9061
rect 3332 9095 3384 9104
rect 3332 9061 3341 9095
rect 3341 9061 3375 9095
rect 3375 9061 3384 9095
rect 3332 9052 3384 9061
rect 4160 9052 4212 9104
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 2412 8984 2464 9036
rect 2964 8984 3016 9036
rect 3056 8984 3108 9036
rect 2688 8916 2740 8968
rect 3148 8848 3200 8900
rect 4896 8984 4948 9036
rect 5540 9052 5592 9104
rect 5356 9027 5408 9036
rect 5356 8993 5390 9027
rect 5390 8993 5408 9027
rect 5356 8984 5408 8993
rect 3332 8848 3384 8900
rect 2780 8780 2832 8832
rect 3240 8780 3292 8832
rect 8208 9120 8260 9172
rect 8760 9163 8812 9172
rect 8760 9129 8769 9163
rect 8769 9129 8803 9163
rect 8803 9129 8812 9163
rect 8760 9120 8812 9129
rect 9220 9163 9272 9172
rect 9220 9129 9229 9163
rect 9229 9129 9263 9163
rect 9263 9129 9272 9163
rect 9220 9120 9272 9129
rect 9496 9120 9548 9172
rect 10140 9120 10192 9172
rect 10324 9120 10376 9172
rect 10508 9120 10560 9172
rect 10692 9120 10744 9172
rect 10784 9120 10836 9172
rect 12348 9120 12400 9172
rect 12900 9120 12952 9172
rect 13452 9120 13504 9172
rect 13912 9120 13964 9172
rect 14188 9120 14240 9172
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 15292 9120 15344 9129
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 7564 9052 7616 9104
rect 8116 9052 8168 9104
rect 7656 9027 7708 9036
rect 7656 8993 7690 9027
rect 7690 8993 7708 9027
rect 6828 8848 6880 8900
rect 7656 8984 7708 8993
rect 8944 8984 8996 9036
rect 8760 8916 8812 8968
rect 9312 8984 9364 9036
rect 9956 8984 10008 9036
rect 8392 8848 8444 8900
rect 9772 8916 9824 8968
rect 12072 9052 12124 9104
rect 12440 9052 12492 9104
rect 13176 9052 13228 9104
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 12992 8984 13044 9036
rect 10784 8916 10836 8968
rect 12532 8916 12584 8968
rect 13084 8916 13136 8968
rect 13636 8916 13688 8968
rect 13820 8916 13872 8968
rect 10784 8823 10836 8832
rect 10784 8789 10793 8823
rect 10793 8789 10827 8823
rect 10827 8789 10836 8823
rect 10784 8780 10836 8789
rect 10968 8780 11020 8832
rect 12348 8823 12400 8832
rect 12348 8789 12357 8823
rect 12357 8789 12391 8823
rect 12391 8789 12400 8823
rect 12348 8780 12400 8789
rect 12716 8780 12768 8832
rect 13544 8823 13596 8832
rect 13544 8789 13553 8823
rect 13553 8789 13587 8823
rect 13587 8789 13596 8823
rect 13544 8780 13596 8789
rect 13820 8780 13872 8832
rect 15200 9052 15252 9104
rect 14648 9027 14700 9036
rect 14648 8993 14657 9027
rect 14657 8993 14691 9027
rect 14691 8993 14700 9027
rect 14648 8984 14700 8993
rect 15292 8984 15344 9036
rect 15660 9120 15712 9172
rect 16304 9163 16356 9172
rect 16304 9129 16313 9163
rect 16313 9129 16347 9163
rect 16347 9129 16356 9163
rect 16304 9120 16356 9129
rect 16396 9120 16448 9172
rect 17408 9120 17460 9172
rect 19248 9120 19300 9172
rect 19340 9120 19392 9172
rect 20720 9120 20772 9172
rect 15568 9052 15620 9104
rect 15660 9027 15712 9036
rect 15660 8993 15669 9027
rect 15669 8993 15703 9027
rect 15703 8993 15712 9027
rect 15660 8984 15712 8993
rect 15936 8984 15988 9036
rect 16396 8984 16448 9036
rect 16580 8984 16632 9036
rect 16948 8984 17000 9036
rect 17592 8984 17644 9036
rect 17776 9027 17828 9036
rect 17776 8993 17785 9027
rect 17785 8993 17819 9027
rect 17819 8993 17828 9027
rect 17776 8984 17828 8993
rect 18052 8984 18104 9036
rect 18604 9027 18656 9036
rect 18604 8993 18638 9027
rect 18638 8993 18656 9027
rect 18604 8984 18656 8993
rect 19984 9027 20036 9036
rect 19984 8993 19993 9027
rect 19993 8993 20027 9027
rect 20027 8993 20036 9027
rect 19984 8984 20036 8993
rect 14740 8916 14792 8968
rect 14832 8916 14884 8968
rect 15108 8916 15160 8968
rect 17040 8916 17092 8968
rect 17960 8959 18012 8968
rect 17960 8925 17969 8959
rect 17969 8925 18003 8959
rect 18003 8925 18012 8959
rect 17960 8916 18012 8925
rect 19340 8916 19392 8968
rect 19892 8916 19944 8968
rect 14096 8780 14148 8832
rect 14280 8780 14332 8832
rect 14648 8780 14700 8832
rect 16396 8848 16448 8900
rect 15568 8780 15620 8832
rect 16672 8780 16724 8832
rect 19432 8848 19484 8900
rect 19616 8848 19668 8900
rect 19800 8780 19852 8832
rect 19984 8780 20036 8832
rect 21272 8780 21324 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2504 8576 2556 8628
rect 3608 8619 3660 8628
rect 3608 8585 3617 8619
rect 3617 8585 3651 8619
rect 3651 8585 3660 8619
rect 3608 8576 3660 8585
rect 5356 8619 5408 8628
rect 5356 8585 5365 8619
rect 5365 8585 5399 8619
rect 5399 8585 5408 8619
rect 5356 8576 5408 8585
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 3240 8508 3292 8560
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2872 8483 2924 8492
rect 2044 8440 2096 8449
rect 1768 8347 1820 8356
rect 1768 8313 1777 8347
rect 1777 8313 1811 8347
rect 1811 8313 1820 8347
rect 1768 8304 1820 8313
rect 1400 8279 1452 8288
rect 1400 8245 1409 8279
rect 1409 8245 1443 8279
rect 1443 8245 1452 8279
rect 1400 8236 1452 8245
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3332 8440 3384 8492
rect 3976 8483 4028 8492
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 5632 8440 5684 8492
rect 3424 8415 3476 8424
rect 3424 8381 3433 8415
rect 3433 8381 3467 8415
rect 3467 8381 3476 8415
rect 3424 8372 3476 8381
rect 9312 8619 9364 8628
rect 9312 8585 9321 8619
rect 9321 8585 9355 8619
rect 9355 8585 9364 8619
rect 9312 8576 9364 8585
rect 10968 8576 11020 8628
rect 12992 8576 13044 8628
rect 18512 8576 18564 8628
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 3516 8304 3568 8356
rect 4160 8304 4212 8356
rect 4344 8304 4396 8356
rect 4712 8304 4764 8356
rect 7104 8347 7156 8356
rect 7104 8313 7138 8347
rect 7138 8313 7156 8347
rect 7104 8304 7156 8313
rect 7380 8372 7432 8424
rect 8024 8372 8076 8424
rect 11428 8508 11480 8560
rect 12808 8508 12860 8560
rect 13084 8508 13136 8560
rect 13912 8508 13964 8560
rect 14740 8508 14792 8560
rect 9312 8440 9364 8492
rect 10232 8440 10284 8492
rect 10416 8440 10468 8492
rect 11336 8440 11388 8492
rect 12348 8440 12400 8492
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 14372 8440 14424 8492
rect 15936 8508 15988 8560
rect 17224 8508 17276 8560
rect 18328 8508 18380 8560
rect 18972 8576 19024 8628
rect 19248 8576 19300 8628
rect 19984 8576 20036 8628
rect 20536 8576 20588 8628
rect 17868 8440 17920 8492
rect 19340 8440 19392 8492
rect 8300 8372 8352 8424
rect 12440 8372 12492 8424
rect 12808 8372 12860 8424
rect 13636 8372 13688 8424
rect 13820 8415 13872 8424
rect 13820 8381 13829 8415
rect 13829 8381 13863 8415
rect 13863 8381 13872 8415
rect 13820 8372 13872 8381
rect 14556 8372 14608 8424
rect 8668 8304 8720 8356
rect 10048 8304 10100 8356
rect 10232 8304 10284 8356
rect 10416 8304 10468 8356
rect 12532 8304 12584 8356
rect 13084 8304 13136 8356
rect 15016 8372 15068 8424
rect 15752 8372 15804 8424
rect 15936 8372 15988 8424
rect 17132 8372 17184 8424
rect 18972 8372 19024 8424
rect 20168 8508 20220 8560
rect 16304 8304 16356 8356
rect 17040 8304 17092 8356
rect 5172 8236 5224 8288
rect 7380 8236 7432 8288
rect 7564 8236 7616 8288
rect 8484 8279 8536 8288
rect 8484 8245 8493 8279
rect 8493 8245 8527 8279
rect 8527 8245 8536 8279
rect 8484 8236 8536 8245
rect 10600 8236 10652 8288
rect 12164 8236 12216 8288
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 12440 8236 12492 8245
rect 13268 8236 13320 8288
rect 13452 8279 13504 8288
rect 13452 8245 13461 8279
rect 13461 8245 13495 8279
rect 13495 8245 13504 8279
rect 13452 8236 13504 8245
rect 19984 8440 20036 8492
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 20444 8372 20496 8424
rect 19800 8304 19852 8356
rect 19432 8279 19484 8288
rect 19432 8245 19441 8279
rect 19441 8245 19475 8279
rect 19475 8245 19484 8279
rect 19432 8236 19484 8245
rect 19616 8236 19668 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 3424 8032 3476 8084
rect 6552 8032 6604 8084
rect 12440 8032 12492 8084
rect 14372 8032 14424 8084
rect 15016 8075 15068 8084
rect 15016 8041 15025 8075
rect 15025 8041 15059 8075
rect 15059 8041 15068 8075
rect 15016 8032 15068 8041
rect 15200 8032 15252 8084
rect 10232 7964 10284 8016
rect 11060 7964 11112 8016
rect 11428 7964 11480 8016
rect 12256 7964 12308 8016
rect 13360 7964 13412 8016
rect 2596 7939 2648 7948
rect 2596 7905 2630 7939
rect 2630 7905 2648 7939
rect 2596 7896 2648 7905
rect 2964 7896 3016 7948
rect 5448 7939 5500 7948
rect 5448 7905 5457 7939
rect 5457 7905 5491 7939
rect 5491 7905 5500 7939
rect 5448 7896 5500 7905
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 1860 7692 1912 7744
rect 4160 7760 4212 7812
rect 4712 7828 4764 7880
rect 5908 7828 5960 7880
rect 7656 7828 7708 7880
rect 5540 7760 5592 7812
rect 3976 7692 4028 7744
rect 4068 7692 4120 7744
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 7656 7692 7708 7744
rect 8024 7896 8076 7948
rect 8208 7939 8260 7948
rect 8208 7905 8242 7939
rect 8242 7905 8260 7939
rect 8208 7896 8260 7905
rect 9128 7896 9180 7948
rect 10692 7896 10744 7948
rect 14096 7964 14148 8016
rect 9220 7828 9272 7880
rect 10416 7828 10468 7880
rect 8944 7760 8996 7812
rect 9404 7760 9456 7812
rect 10048 7760 10100 7812
rect 10232 7760 10284 7812
rect 12992 7828 13044 7880
rect 13636 7896 13688 7948
rect 14648 7896 14700 7948
rect 15016 7896 15068 7948
rect 17040 7896 17092 7948
rect 17868 8032 17920 8084
rect 18052 8032 18104 8084
rect 18328 8032 18380 8084
rect 17960 7964 18012 8016
rect 15752 7871 15804 7880
rect 15752 7837 15761 7871
rect 15761 7837 15795 7871
rect 15795 7837 15804 7871
rect 15752 7828 15804 7837
rect 17224 7896 17276 7948
rect 17684 7896 17736 7948
rect 19340 7964 19392 8016
rect 19892 8032 19944 8084
rect 20168 8032 20220 8084
rect 8852 7692 8904 7744
rect 9220 7692 9272 7744
rect 9680 7692 9732 7744
rect 10600 7692 10652 7744
rect 10876 7692 10928 7744
rect 13084 7760 13136 7812
rect 11980 7735 12032 7744
rect 11980 7701 11989 7735
rect 11989 7701 12023 7735
rect 12023 7701 12032 7735
rect 11980 7692 12032 7701
rect 12256 7735 12308 7744
rect 12256 7701 12265 7735
rect 12265 7701 12299 7735
rect 12299 7701 12308 7735
rect 12256 7692 12308 7701
rect 12440 7692 12492 7744
rect 12900 7692 12952 7744
rect 16212 7760 16264 7812
rect 14740 7692 14792 7744
rect 15936 7692 15988 7744
rect 18696 7760 18748 7812
rect 19984 7896 20036 7948
rect 20352 7964 20404 8016
rect 21088 7964 21140 8016
rect 20536 7896 20588 7948
rect 20352 7871 20404 7880
rect 20352 7837 20361 7871
rect 20361 7837 20395 7871
rect 20395 7837 20404 7871
rect 20352 7828 20404 7837
rect 20720 7760 20772 7812
rect 18604 7692 18656 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 2688 7488 2740 7540
rect 4712 7488 4764 7540
rect 5172 7531 5224 7540
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 5448 7531 5500 7540
rect 5448 7497 5457 7531
rect 5457 7497 5491 7531
rect 5491 7497 5500 7531
rect 5448 7488 5500 7497
rect 6276 7488 6328 7540
rect 8576 7488 8628 7540
rect 6644 7420 6696 7472
rect 7104 7420 7156 7472
rect 8208 7420 8260 7472
rect 9220 7420 9272 7472
rect 9588 7488 9640 7540
rect 16396 7531 16448 7540
rect 10232 7420 10284 7472
rect 10968 7420 11020 7472
rect 12256 7420 12308 7472
rect 14188 7420 14240 7472
rect 5172 7352 5224 7404
rect 6920 7352 6972 7404
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 10508 7395 10560 7404
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 11612 7352 11664 7404
rect 1860 7284 1912 7336
rect 2044 7327 2096 7336
rect 2044 7293 2078 7327
rect 2078 7293 2096 7327
rect 2044 7284 2096 7293
rect 3884 7284 3936 7336
rect 6092 7284 6144 7336
rect 7932 7284 7984 7336
rect 8300 7284 8352 7336
rect 10968 7284 11020 7336
rect 3332 7216 3384 7268
rect 4712 7216 4764 7268
rect 4896 7216 4948 7268
rect 8208 7216 8260 7268
rect 8944 7216 8996 7268
rect 9496 7216 9548 7268
rect 9680 7216 9732 7268
rect 10416 7216 10468 7268
rect 11520 7284 11572 7336
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 12532 7284 12584 7336
rect 14372 7352 14424 7404
rect 13728 7284 13780 7336
rect 16396 7497 16405 7531
rect 16405 7497 16439 7531
rect 16439 7497 16448 7531
rect 16396 7488 16448 7497
rect 17960 7488 18012 7540
rect 19156 7488 19208 7540
rect 19616 7488 19668 7540
rect 14740 7420 14792 7472
rect 14648 7395 14700 7404
rect 14648 7361 14657 7395
rect 14657 7361 14691 7395
rect 14691 7361 14700 7395
rect 14648 7352 14700 7361
rect 15108 7352 15160 7404
rect 15844 7395 15896 7404
rect 15844 7361 15853 7395
rect 15853 7361 15887 7395
rect 15887 7361 15896 7395
rect 15844 7352 15896 7361
rect 16028 7395 16080 7404
rect 16028 7361 16037 7395
rect 16037 7361 16071 7395
rect 16071 7361 16080 7395
rect 16028 7352 16080 7361
rect 16212 7352 16264 7404
rect 17684 7352 17736 7404
rect 11612 7216 11664 7268
rect 13544 7216 13596 7268
rect 2044 7148 2096 7200
rect 2412 7148 2464 7200
rect 3792 7148 3844 7200
rect 7748 7148 7800 7200
rect 8852 7148 8904 7200
rect 9588 7148 9640 7200
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 10232 7191 10284 7200
rect 10232 7157 10241 7191
rect 10241 7157 10275 7191
rect 10275 7157 10284 7191
rect 10232 7148 10284 7157
rect 10876 7191 10928 7200
rect 10876 7157 10885 7191
rect 10885 7157 10919 7191
rect 10919 7157 10928 7191
rect 10876 7148 10928 7157
rect 10968 7148 11020 7200
rect 11428 7148 11480 7200
rect 13820 7191 13872 7200
rect 13820 7157 13829 7191
rect 13829 7157 13863 7191
rect 13863 7157 13872 7191
rect 13820 7148 13872 7157
rect 17500 7284 17552 7336
rect 19340 7352 19392 7404
rect 19432 7352 19484 7404
rect 20352 7420 20404 7472
rect 19800 7352 19852 7404
rect 18512 7284 18564 7336
rect 21088 7284 21140 7336
rect 19800 7216 19852 7268
rect 15660 7148 15712 7200
rect 15936 7148 15988 7200
rect 16212 7148 16264 7200
rect 18052 7191 18104 7200
rect 18052 7157 18061 7191
rect 18061 7157 18095 7191
rect 18095 7157 18104 7191
rect 18052 7148 18104 7157
rect 19248 7148 19300 7200
rect 19616 7148 19668 7200
rect 21640 7148 21692 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 1400 6944 1452 6996
rect 3608 6987 3660 6996
rect 3608 6953 3617 6987
rect 3617 6953 3651 6987
rect 3651 6953 3660 6987
rect 3608 6944 3660 6953
rect 5816 6944 5868 6996
rect 1676 6808 1728 6860
rect 2228 6672 2280 6724
rect 3700 6876 3752 6928
rect 7196 6876 7248 6928
rect 7288 6876 7340 6928
rect 7748 6876 7800 6928
rect 2504 6808 2556 6860
rect 2596 6740 2648 6792
rect 4252 6808 4304 6860
rect 5540 6808 5592 6860
rect 6368 6808 6420 6860
rect 8576 6808 8628 6860
rect 9220 6944 9272 6996
rect 9864 6944 9916 6996
rect 10876 6944 10928 6996
rect 11244 6987 11296 6996
rect 11244 6953 11253 6987
rect 11253 6953 11287 6987
rect 11287 6953 11296 6987
rect 11244 6944 11296 6953
rect 11520 6944 11572 6996
rect 11612 6944 11664 6996
rect 11152 6876 11204 6928
rect 12808 6944 12860 6996
rect 13360 6944 13412 6996
rect 13728 6944 13780 6996
rect 14464 6944 14516 6996
rect 15108 6944 15160 6996
rect 15660 6987 15712 6996
rect 15660 6953 15669 6987
rect 15669 6953 15703 6987
rect 15703 6953 15712 6987
rect 15660 6944 15712 6953
rect 12164 6876 12216 6928
rect 15476 6876 15528 6928
rect 5172 6740 5224 6792
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6736 6783 6788 6792
rect 6552 6740 6604 6749
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 7472 6740 7524 6792
rect 7288 6715 7340 6724
rect 7288 6681 7297 6715
rect 7297 6681 7331 6715
rect 7331 6681 7340 6715
rect 7288 6672 7340 6681
rect 2964 6604 3016 6656
rect 5540 6604 5592 6656
rect 5632 6604 5684 6656
rect 6368 6604 6420 6656
rect 6920 6604 6972 6656
rect 8116 6740 8168 6792
rect 8944 6740 8996 6792
rect 9312 6740 9364 6792
rect 7840 6672 7892 6724
rect 11888 6808 11940 6860
rect 14280 6851 14332 6860
rect 10324 6740 10376 6792
rect 11428 6740 11480 6792
rect 11612 6740 11664 6792
rect 11980 6740 12032 6792
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 10232 6604 10284 6656
rect 10416 6604 10468 6656
rect 10968 6604 11020 6656
rect 12624 6672 12676 6724
rect 12992 6672 13044 6724
rect 14280 6817 14289 6851
rect 14289 6817 14323 6851
rect 14323 6817 14332 6851
rect 14280 6808 14332 6817
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 15752 6783 15804 6792
rect 15752 6749 15761 6783
rect 15761 6749 15795 6783
rect 15795 6749 15804 6783
rect 15752 6740 15804 6749
rect 16028 6740 16080 6792
rect 16304 6851 16356 6860
rect 16304 6817 16313 6851
rect 16313 6817 16347 6851
rect 16347 6817 16356 6851
rect 18052 6944 18104 6996
rect 19340 6944 19392 6996
rect 16304 6808 16356 6817
rect 19248 6808 19300 6860
rect 19432 6851 19484 6860
rect 19432 6817 19466 6851
rect 19466 6817 19484 6851
rect 19432 6808 19484 6817
rect 17040 6740 17092 6792
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 18604 6740 18656 6792
rect 19156 6783 19208 6792
rect 19156 6749 19165 6783
rect 19165 6749 19199 6783
rect 19199 6749 19208 6783
rect 19156 6740 19208 6749
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 17684 6672 17736 6724
rect 15200 6604 15252 6656
rect 15384 6604 15436 6656
rect 16304 6604 16356 6656
rect 17408 6604 17460 6656
rect 17868 6604 17920 6656
rect 20168 6672 20220 6724
rect 19432 6604 19484 6656
rect 20444 6604 20496 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 1952 6400 2004 6452
rect 5080 6400 5132 6452
rect 6644 6400 6696 6452
rect 3332 6375 3384 6384
rect 3332 6341 3341 6375
rect 3341 6341 3375 6375
rect 3375 6341 3384 6375
rect 3332 6332 3384 6341
rect 4896 6375 4948 6384
rect 4896 6341 4905 6375
rect 4905 6341 4939 6375
rect 4939 6341 4948 6375
rect 4896 6332 4948 6341
rect 3516 6264 3568 6316
rect 4620 6264 4672 6316
rect 5448 6264 5500 6316
rect 6368 6264 6420 6316
rect 8668 6400 8720 6452
rect 9680 6400 9732 6452
rect 8484 6332 8536 6384
rect 9128 6332 9180 6384
rect 9312 6332 9364 6384
rect 1584 6196 1636 6248
rect 1860 6196 1912 6248
rect 4804 6196 4856 6248
rect 4896 6196 4948 6248
rect 5264 6196 5316 6248
rect 5632 6239 5684 6248
rect 5632 6205 5641 6239
rect 5641 6205 5675 6239
rect 5675 6205 5684 6239
rect 5632 6196 5684 6205
rect 6460 6196 6512 6248
rect 8392 6307 8444 6316
rect 8392 6273 8401 6307
rect 8401 6273 8435 6307
rect 8435 6273 8444 6307
rect 8392 6264 8444 6273
rect 8668 6264 8720 6316
rect 8300 6196 8352 6248
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 9404 6307 9456 6316
rect 9404 6273 9413 6307
rect 9413 6273 9447 6307
rect 9447 6273 9456 6307
rect 9404 6264 9456 6273
rect 11980 6400 12032 6452
rect 12164 6400 12216 6452
rect 10876 6332 10928 6384
rect 14464 6400 14516 6452
rect 18788 6400 18840 6452
rect 19524 6400 19576 6452
rect 20444 6400 20496 6452
rect 14004 6375 14056 6384
rect 14004 6341 14013 6375
rect 14013 6341 14047 6375
rect 14047 6341 14056 6375
rect 14004 6332 14056 6341
rect 16028 6332 16080 6384
rect 9680 6196 9732 6248
rect 12348 6196 12400 6248
rect 12440 6196 12492 6248
rect 12624 6239 12676 6248
rect 12624 6205 12633 6239
rect 12633 6205 12667 6239
rect 12667 6205 12676 6239
rect 12624 6196 12676 6205
rect 13728 6264 13780 6316
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 17684 6264 17736 6316
rect 18420 6264 18472 6316
rect 18604 6307 18656 6316
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 18604 6264 18656 6273
rect 18788 6264 18840 6316
rect 19156 6264 19208 6316
rect 14280 6196 14332 6248
rect 14464 6239 14516 6248
rect 2412 6128 2464 6180
rect 7104 6128 7156 6180
rect 3332 6060 3384 6112
rect 5632 6060 5684 6112
rect 6184 6060 6236 6112
rect 7288 6060 7340 6112
rect 7748 6103 7800 6112
rect 7748 6069 7757 6103
rect 7757 6069 7791 6103
rect 7791 6069 7800 6103
rect 7748 6060 7800 6069
rect 9128 6103 9180 6112
rect 9128 6069 9137 6103
rect 9137 6069 9171 6103
rect 9171 6069 9180 6103
rect 9128 6060 9180 6069
rect 11612 6128 11664 6180
rect 13820 6128 13872 6180
rect 14188 6128 14240 6180
rect 14464 6205 14473 6239
rect 14473 6205 14507 6239
rect 14507 6205 14516 6239
rect 14464 6196 14516 6205
rect 15844 6196 15896 6248
rect 15384 6128 15436 6180
rect 15936 6128 15988 6180
rect 10968 6060 11020 6112
rect 12532 6060 12584 6112
rect 12808 6060 12860 6112
rect 15660 6060 15712 6112
rect 17868 6060 17920 6112
rect 18052 6103 18104 6112
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 19432 6128 19484 6180
rect 20168 6128 20220 6180
rect 21824 6060 21876 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 1768 5899 1820 5908
rect 1768 5865 1777 5899
rect 1777 5865 1811 5899
rect 1811 5865 1820 5899
rect 1768 5856 1820 5865
rect 3976 5856 4028 5908
rect 5448 5899 5500 5908
rect 5448 5865 5457 5899
rect 5457 5865 5491 5899
rect 5491 5865 5500 5899
rect 5448 5856 5500 5865
rect 4252 5788 4304 5840
rect 7196 5899 7248 5908
rect 7196 5865 7205 5899
rect 7205 5865 7239 5899
rect 7239 5865 7248 5899
rect 7196 5856 7248 5865
rect 7472 5856 7524 5908
rect 12348 5856 12400 5908
rect 12440 5856 12492 5908
rect 14096 5856 14148 5908
rect 14188 5856 14240 5908
rect 15016 5856 15068 5908
rect 16212 5856 16264 5908
rect 8576 5831 8628 5840
rect 8576 5797 8585 5831
rect 8585 5797 8619 5831
rect 8619 5797 8628 5831
rect 8576 5788 8628 5797
rect 5080 5720 5132 5772
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 6552 5720 6604 5729
rect 7288 5720 7340 5772
rect 10508 5788 10560 5840
rect 10968 5788 11020 5840
rect 11888 5788 11940 5840
rect 6828 5695 6880 5704
rect 1860 5516 1912 5568
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 8944 5720 8996 5772
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 9772 5720 9824 5772
rect 11704 5763 11756 5772
rect 6736 5584 6788 5636
rect 7472 5584 7524 5636
rect 8392 5652 8444 5704
rect 7748 5584 7800 5636
rect 8300 5584 8352 5636
rect 9312 5652 9364 5704
rect 10968 5652 11020 5704
rect 11152 5652 11204 5704
rect 11704 5729 11713 5763
rect 11713 5729 11747 5763
rect 11747 5729 11756 5763
rect 11704 5720 11756 5729
rect 12992 5788 13044 5840
rect 14004 5788 14056 5840
rect 12440 5720 12492 5772
rect 16396 5720 16448 5772
rect 17960 5856 18012 5908
rect 18052 5856 18104 5908
rect 19340 5899 19392 5908
rect 19340 5865 19349 5899
rect 19349 5865 19383 5899
rect 19383 5865 19392 5899
rect 19340 5856 19392 5865
rect 19432 5856 19484 5908
rect 12256 5652 12308 5704
rect 14832 5652 14884 5704
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 17500 5720 17552 5772
rect 16028 5652 16080 5661
rect 3516 5516 3568 5568
rect 4068 5516 4120 5568
rect 6092 5516 6144 5568
rect 6920 5516 6972 5568
rect 9680 5584 9732 5636
rect 10692 5584 10744 5636
rect 12440 5584 12492 5636
rect 12532 5584 12584 5636
rect 9588 5516 9640 5568
rect 10324 5516 10376 5568
rect 11152 5516 11204 5568
rect 12348 5516 12400 5568
rect 12808 5516 12860 5568
rect 17960 5652 18012 5704
rect 18144 5720 18196 5772
rect 14556 5516 14608 5568
rect 14648 5516 14700 5568
rect 17868 5584 17920 5636
rect 19708 5584 19760 5636
rect 20996 5720 21048 5772
rect 19984 5695 20036 5704
rect 19984 5661 19993 5695
rect 19993 5661 20027 5695
rect 20027 5661 20036 5695
rect 19984 5652 20036 5661
rect 17684 5516 17736 5568
rect 18696 5516 18748 5568
rect 20076 5516 20128 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 3332 5355 3384 5364
rect 3332 5321 3341 5355
rect 3341 5321 3375 5355
rect 3375 5321 3384 5355
rect 3332 5312 3384 5321
rect 7196 5312 7248 5364
rect 8208 5355 8260 5364
rect 8208 5321 8217 5355
rect 8217 5321 8251 5355
rect 8251 5321 8260 5355
rect 8208 5312 8260 5321
rect 9496 5312 9548 5364
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 2964 5176 3016 5228
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 4620 5176 4672 5228
rect 5080 5176 5132 5228
rect 5264 5176 5316 5228
rect 6828 5244 6880 5296
rect 9772 5312 9824 5364
rect 10140 5312 10192 5364
rect 13544 5312 13596 5364
rect 14832 5312 14884 5364
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 3240 5108 3292 5160
rect 5540 5108 5592 5160
rect 6736 5108 6788 5160
rect 9956 5176 10008 5228
rect 10876 5176 10928 5228
rect 11152 5176 11204 5228
rect 11704 5244 11756 5296
rect 12256 5244 12308 5296
rect 8576 5108 8628 5160
rect 8668 5108 8720 5160
rect 9588 5108 9640 5160
rect 10692 5108 10744 5160
rect 12808 5176 12860 5228
rect 15292 5244 15344 5296
rect 14188 5219 14240 5228
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 14372 5176 14424 5228
rect 15384 5219 15436 5228
rect 15384 5185 15393 5219
rect 15393 5185 15427 5219
rect 15427 5185 15436 5219
rect 15384 5176 15436 5185
rect 15936 5312 15988 5364
rect 16396 5312 16448 5364
rect 17500 5312 17552 5364
rect 18972 5312 19024 5364
rect 19984 5312 20036 5364
rect 20168 5355 20220 5364
rect 20168 5321 20177 5355
rect 20177 5321 20211 5355
rect 20211 5321 20220 5355
rect 20168 5312 20220 5321
rect 16948 5244 17000 5296
rect 18788 5219 18840 5228
rect 18788 5185 18797 5219
rect 18797 5185 18831 5219
rect 18831 5185 18840 5219
rect 18788 5176 18840 5185
rect 19800 5176 19852 5228
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 2504 5015 2556 5024
rect 2504 4981 2513 5015
rect 2513 4981 2547 5015
rect 2547 4981 2556 5015
rect 2504 4972 2556 4981
rect 2596 5015 2648 5024
rect 2596 4981 2605 5015
rect 2605 4981 2639 5015
rect 2639 4981 2648 5015
rect 2596 4972 2648 4981
rect 4068 4972 4120 5024
rect 5724 5040 5776 5092
rect 4712 5015 4764 5024
rect 4712 4981 4721 5015
rect 4721 4981 4755 5015
rect 4755 4981 4764 5015
rect 4712 4972 4764 4981
rect 6184 5015 6236 5024
rect 6184 4981 6193 5015
rect 6193 4981 6227 5015
rect 6227 4981 6236 5015
rect 6184 4972 6236 4981
rect 7564 5040 7616 5092
rect 8576 4972 8628 5024
rect 9220 5040 9272 5092
rect 10232 5040 10284 5092
rect 10508 5040 10560 5092
rect 11888 5108 11940 5160
rect 12256 5108 12308 5160
rect 15016 5108 15068 5160
rect 16028 5151 16080 5160
rect 16028 5117 16062 5151
rect 16062 5117 16080 5151
rect 16028 5108 16080 5117
rect 11980 5040 12032 5092
rect 12992 5040 13044 5092
rect 9864 4972 9916 5024
rect 9956 4972 10008 5024
rect 11428 4972 11480 5024
rect 12440 5015 12492 5024
rect 12440 4981 12449 5015
rect 12449 4981 12483 5015
rect 12483 4981 12492 5015
rect 12440 4972 12492 4981
rect 12900 4972 12952 5024
rect 13820 4972 13872 5024
rect 14372 5040 14424 5092
rect 15292 5040 15344 5092
rect 17224 5108 17276 5160
rect 17408 5151 17460 5160
rect 17408 5117 17417 5151
rect 17417 5117 17451 5151
rect 17451 5117 17460 5151
rect 17408 5108 17460 5117
rect 20444 5151 20496 5160
rect 16304 5040 16356 5092
rect 20444 5117 20453 5151
rect 20453 5117 20487 5151
rect 20487 5117 20496 5151
rect 20444 5108 20496 5117
rect 15844 4972 15896 5024
rect 19892 5040 19944 5092
rect 19248 4972 19300 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 2412 4768 2464 4820
rect 2688 4768 2740 4820
rect 3424 4768 3476 4820
rect 4068 4811 4120 4820
rect 4068 4777 4077 4811
rect 4077 4777 4111 4811
rect 4111 4777 4120 4811
rect 4068 4768 4120 4777
rect 6644 4768 6696 4820
rect 6828 4768 6880 4820
rect 7288 4811 7340 4820
rect 7288 4777 7297 4811
rect 7297 4777 7331 4811
rect 7331 4777 7340 4811
rect 7288 4768 7340 4777
rect 7656 4811 7708 4820
rect 7656 4777 7665 4811
rect 7665 4777 7699 4811
rect 7699 4777 7708 4811
rect 7656 4768 7708 4777
rect 8576 4768 8628 4820
rect 10508 4768 10560 4820
rect 10692 4768 10744 4820
rect 11428 4768 11480 4820
rect 12440 4768 12492 4820
rect 13820 4811 13872 4820
rect 13820 4777 13829 4811
rect 13829 4777 13863 4811
rect 13863 4777 13872 4811
rect 13820 4768 13872 4777
rect 15752 4768 15804 4820
rect 16580 4768 16632 4820
rect 2964 4632 3016 4684
rect 3424 4675 3476 4684
rect 3424 4641 3433 4675
rect 3433 4641 3467 4675
rect 3467 4641 3476 4675
rect 3424 4632 3476 4641
rect 2872 4564 2924 4616
rect 3976 4564 4028 4616
rect 5724 4632 5776 4684
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 9680 4632 9732 4684
rect 1860 4428 1912 4480
rect 8392 4564 8444 4616
rect 10508 4632 10560 4684
rect 11612 4700 11664 4752
rect 17960 4768 18012 4820
rect 19340 4768 19392 4820
rect 19800 4768 19852 4820
rect 17684 4700 17736 4752
rect 18512 4700 18564 4752
rect 21180 4700 21232 4752
rect 10876 4632 10928 4684
rect 6644 4496 6696 4548
rect 9496 4496 9548 4548
rect 11520 4632 11572 4684
rect 11704 4564 11756 4616
rect 12164 4632 12216 4684
rect 13636 4632 13688 4684
rect 14556 4632 14608 4684
rect 14648 4675 14700 4684
rect 14648 4641 14657 4675
rect 14657 4641 14691 4675
rect 14691 4641 14700 4675
rect 14648 4632 14700 4641
rect 12072 4564 12124 4616
rect 14372 4564 14424 4616
rect 9864 4428 9916 4480
rect 10048 4471 10100 4480
rect 10048 4437 10057 4471
rect 10057 4437 10091 4471
rect 10091 4437 10100 4471
rect 10048 4428 10100 4437
rect 11612 4428 11664 4480
rect 12900 4428 12952 4480
rect 13268 4428 13320 4480
rect 15384 4564 15436 4616
rect 15568 4564 15620 4616
rect 16028 4564 16080 4616
rect 15200 4496 15252 4548
rect 16396 4632 16448 4684
rect 17132 4675 17184 4684
rect 17132 4641 17141 4675
rect 17141 4641 17175 4675
rect 17175 4641 17184 4675
rect 17132 4632 17184 4641
rect 19432 4675 19484 4684
rect 19432 4641 19441 4675
rect 19441 4641 19475 4675
rect 19475 4641 19484 4675
rect 19432 4632 19484 4641
rect 19984 4632 20036 4684
rect 20812 4632 20864 4684
rect 16580 4607 16632 4616
rect 16580 4573 16589 4607
rect 16589 4573 16623 4607
rect 16623 4573 16632 4607
rect 16580 4564 16632 4573
rect 19340 4564 19392 4616
rect 19892 4564 19944 4616
rect 20352 4607 20404 4616
rect 20352 4573 20361 4607
rect 20361 4573 20395 4607
rect 20395 4573 20404 4607
rect 20352 4564 20404 4573
rect 20536 4564 20588 4616
rect 16212 4428 16264 4480
rect 18972 4428 19024 4480
rect 20076 4428 20128 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 3424 4224 3476 4276
rect 4712 4224 4764 4276
rect 7104 4224 7156 4276
rect 7564 4224 7616 4276
rect 8208 4224 8260 4276
rect 10048 4224 10100 4276
rect 13268 4224 13320 4276
rect 13360 4224 13412 4276
rect 6828 4156 6880 4208
rect 2964 4088 3016 4140
rect 3424 4131 3476 4140
rect 3424 4097 3433 4131
rect 3433 4097 3467 4131
rect 3467 4097 3476 4131
rect 3424 4088 3476 4097
rect 4436 4088 4488 4140
rect 5080 4088 5132 4140
rect 6920 4088 6972 4140
rect 8116 4088 8168 4140
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 9588 4088 9640 4140
rect 10968 4156 11020 4208
rect 14372 4224 14424 4276
rect 14556 4224 14608 4276
rect 14924 4224 14976 4276
rect 11612 4131 11664 4140
rect 4712 4020 4764 4072
rect 5264 4063 5316 4072
rect 3148 3952 3200 4004
rect 5264 4029 5273 4063
rect 5273 4029 5307 4063
rect 5307 4029 5316 4063
rect 5264 4020 5316 4029
rect 6276 4020 6328 4072
rect 7196 4063 7248 4072
rect 7196 4029 7205 4063
rect 7205 4029 7239 4063
rect 7239 4029 7248 4063
rect 7196 4020 7248 4029
rect 8024 4063 8076 4072
rect 8024 4029 8033 4063
rect 8033 4029 8067 4063
rect 8067 4029 8076 4063
rect 8024 4020 8076 4029
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 3332 3927 3384 3936
rect 3332 3893 3341 3927
rect 3341 3893 3375 3927
rect 3375 3893 3384 3927
rect 3332 3884 3384 3893
rect 4160 3884 4212 3936
rect 4252 3884 4304 3936
rect 5172 3952 5224 4004
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 11612 4097 11621 4131
rect 11621 4097 11655 4131
rect 11655 4097 11664 4131
rect 11612 4088 11664 4097
rect 14188 4156 14240 4208
rect 12072 4088 12124 4140
rect 10508 4063 10560 4072
rect 10508 4029 10517 4063
rect 10517 4029 10551 4063
rect 10551 4029 10560 4063
rect 10508 4020 10560 4029
rect 10784 4020 10836 4072
rect 12624 4088 12676 4140
rect 15016 4088 15068 4140
rect 15476 4224 15528 4276
rect 16856 4224 16908 4276
rect 17040 4156 17092 4208
rect 17132 4156 17184 4208
rect 19616 4224 19668 4276
rect 20444 4224 20496 4276
rect 16396 4131 16448 4140
rect 12532 4063 12584 4072
rect 12532 4029 12541 4063
rect 12541 4029 12575 4063
rect 12575 4029 12584 4063
rect 12532 4020 12584 4029
rect 10600 3952 10652 4004
rect 11428 3952 11480 4004
rect 12440 3952 12492 4004
rect 16396 4097 16405 4131
rect 16405 4097 16439 4131
rect 16439 4097 16448 4131
rect 16396 4088 16448 4097
rect 13360 3995 13412 4004
rect 13360 3961 13394 3995
rect 13394 3961 13412 3995
rect 13360 3952 13412 3961
rect 13820 3952 13872 4004
rect 14924 3952 14976 4004
rect 15016 3952 15068 4004
rect 9220 3884 9272 3936
rect 10232 3884 10284 3936
rect 11796 3884 11848 3936
rect 12532 3884 12584 3936
rect 12992 3884 13044 3936
rect 13084 3884 13136 3936
rect 14464 3884 14516 3936
rect 15476 3884 15528 3936
rect 15752 3927 15804 3936
rect 15752 3893 15761 3927
rect 15761 3893 15795 3927
rect 15795 3893 15804 3927
rect 15752 3884 15804 3893
rect 15844 3884 15896 3936
rect 17132 3927 17184 3936
rect 17132 3893 17141 3927
rect 17141 3893 17175 3927
rect 17175 3893 17184 3927
rect 17132 3884 17184 3893
rect 17684 4088 17736 4140
rect 20168 4156 20220 4208
rect 19156 4020 19208 4072
rect 19524 4020 19576 4072
rect 20076 4063 20128 4072
rect 20076 4029 20085 4063
rect 20085 4029 20119 4063
rect 20119 4029 20128 4063
rect 20076 4020 20128 4029
rect 20812 4020 20864 4072
rect 17408 3952 17460 4004
rect 17684 3884 17736 3936
rect 18696 3952 18748 4004
rect 19708 3952 19760 4004
rect 19892 3884 19944 3936
rect 20444 3884 20496 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 940 3680 992 3732
rect 2872 3680 2924 3732
rect 3332 3680 3384 3732
rect 4252 3723 4304 3732
rect 4252 3689 4261 3723
rect 4261 3689 4295 3723
rect 4295 3689 4304 3723
rect 4252 3680 4304 3689
rect 4712 3680 4764 3732
rect 8300 3680 8352 3732
rect 3332 3544 3384 3596
rect 4160 3544 4212 3596
rect 1492 3519 1544 3528
rect 1492 3485 1501 3519
rect 1501 3485 1535 3519
rect 1535 3485 1544 3519
rect 1492 3476 1544 3485
rect 1952 3519 2004 3528
rect 1952 3485 1961 3519
rect 1961 3485 1995 3519
rect 1995 3485 2004 3519
rect 1952 3476 2004 3485
rect 3148 3476 3200 3528
rect 2964 3340 3016 3392
rect 4252 3476 4304 3528
rect 5540 3544 5592 3596
rect 6920 3544 6972 3596
rect 7748 3612 7800 3664
rect 8116 3655 8168 3664
rect 8116 3621 8125 3655
rect 8125 3621 8159 3655
rect 8159 3621 8168 3655
rect 8116 3612 8168 3621
rect 7564 3544 7616 3596
rect 9128 3680 9180 3732
rect 9680 3723 9732 3732
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 10324 3680 10376 3732
rect 10876 3680 10928 3732
rect 11336 3680 11388 3732
rect 11520 3680 11572 3732
rect 12440 3723 12492 3732
rect 12440 3689 12449 3723
rect 12449 3689 12483 3723
rect 12483 3689 12492 3723
rect 12440 3680 12492 3689
rect 13912 3723 13964 3732
rect 13912 3689 13921 3723
rect 13921 3689 13955 3723
rect 13955 3689 13964 3723
rect 13912 3680 13964 3689
rect 15752 3680 15804 3732
rect 9220 3612 9272 3664
rect 12900 3655 12952 3664
rect 8668 3544 8720 3596
rect 9404 3544 9456 3596
rect 11888 3544 11940 3596
rect 12900 3621 12909 3655
rect 12909 3621 12943 3655
rect 12943 3621 12952 3655
rect 12900 3612 12952 3621
rect 13544 3612 13596 3664
rect 13636 3544 13688 3596
rect 14464 3587 14516 3596
rect 5172 3476 5224 3528
rect 5264 3476 5316 3528
rect 7104 3519 7156 3528
rect 7104 3485 7113 3519
rect 7113 3485 7147 3519
rect 7147 3485 7156 3519
rect 7104 3476 7156 3485
rect 7196 3476 7248 3528
rect 8392 3476 8444 3528
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10784 3519 10836 3528
rect 10232 3476 10284 3485
rect 10784 3485 10793 3519
rect 10793 3485 10827 3519
rect 10827 3485 10836 3519
rect 10784 3476 10836 3485
rect 12164 3476 12216 3528
rect 6368 3408 6420 3460
rect 6276 3340 6328 3392
rect 7656 3383 7708 3392
rect 7656 3349 7665 3383
rect 7665 3349 7699 3383
rect 7699 3349 7708 3383
rect 7656 3340 7708 3349
rect 8208 3340 8260 3392
rect 8852 3340 8904 3392
rect 8944 3340 8996 3392
rect 10416 3340 10468 3392
rect 12624 3408 12676 3460
rect 14464 3553 14473 3587
rect 14473 3553 14507 3587
rect 14507 3553 14516 3587
rect 14464 3544 14516 3553
rect 16580 3612 16632 3664
rect 17960 3680 18012 3732
rect 18604 3680 18656 3732
rect 19340 3680 19392 3732
rect 19524 3723 19576 3732
rect 19524 3689 19533 3723
rect 19533 3689 19567 3723
rect 19567 3689 19576 3723
rect 19524 3680 19576 3689
rect 19800 3680 19852 3732
rect 20168 3680 20220 3732
rect 15936 3544 15988 3596
rect 16396 3544 16448 3596
rect 17316 3544 17368 3596
rect 14372 3476 14424 3528
rect 16856 3476 16908 3528
rect 18696 3519 18748 3528
rect 18696 3485 18705 3519
rect 18705 3485 18739 3519
rect 18739 3485 18748 3519
rect 19800 3519 19852 3528
rect 18696 3476 18748 3485
rect 19800 3485 19809 3519
rect 19809 3485 19843 3519
rect 19843 3485 19852 3519
rect 19800 3476 19852 3485
rect 12164 3383 12216 3392
rect 12164 3349 12173 3383
rect 12173 3349 12207 3383
rect 12207 3349 12216 3383
rect 12164 3340 12216 3349
rect 12900 3340 12952 3392
rect 13268 3340 13320 3392
rect 14556 3340 14608 3392
rect 15476 3383 15528 3392
rect 15476 3349 15485 3383
rect 15485 3349 15519 3383
rect 15519 3349 15528 3383
rect 15476 3340 15528 3349
rect 17408 3340 17460 3392
rect 17868 3340 17920 3392
rect 19708 3340 19760 3392
rect 20076 3340 20128 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 2504 3136 2556 3188
rect 2596 3136 2648 3188
rect 3332 3136 3384 3188
rect 5264 3179 5316 3188
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 6184 3136 6236 3188
rect 8392 3136 8444 3188
rect 8852 3136 8904 3188
rect 10968 3136 11020 3188
rect 12348 3136 12400 3188
rect 12624 3136 12676 3188
rect 13268 3136 13320 3188
rect 13728 3179 13780 3188
rect 13728 3145 13737 3179
rect 13737 3145 13771 3179
rect 13771 3145 13780 3179
rect 13728 3136 13780 3145
rect 14004 3136 14056 3188
rect 14372 3136 14424 3188
rect 14740 3136 14792 3188
rect 15016 3136 15068 3188
rect 12072 3111 12124 3120
rect 12072 3077 12081 3111
rect 12081 3077 12115 3111
rect 12115 3077 12124 3111
rect 12072 3068 12124 3077
rect 16120 3136 16172 3188
rect 17132 3136 17184 3188
rect 17224 3136 17276 3188
rect 3332 3043 3384 3052
rect 3332 3009 3341 3043
rect 3341 3009 3375 3043
rect 3375 3009 3384 3043
rect 3332 3000 3384 3009
rect 5724 3000 5776 3052
rect 6368 3000 6420 3052
rect 1492 2932 1544 2984
rect 3792 2932 3844 2984
rect 1676 2864 1728 2916
rect 5816 2932 5868 2984
rect 6736 2932 6788 2984
rect 8576 2932 8628 2984
rect 10232 3000 10284 3052
rect 11980 3000 12032 3052
rect 13084 3043 13136 3052
rect 10140 2975 10192 2984
rect 10140 2941 10149 2975
rect 10149 2941 10183 2975
rect 10183 2941 10192 2975
rect 10140 2932 10192 2941
rect 10784 2932 10836 2984
rect 12164 2932 12216 2984
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 13360 3000 13412 3052
rect 13728 3000 13780 3052
rect 14004 3000 14056 3052
rect 14464 3043 14516 3052
rect 14464 3009 14473 3043
rect 14473 3009 14507 3043
rect 14507 3009 14516 3043
rect 14464 3000 14516 3009
rect 14740 3000 14792 3052
rect 17776 3068 17828 3120
rect 18512 3136 18564 3188
rect 19432 3179 19484 3188
rect 19432 3145 19441 3179
rect 19441 3145 19475 3179
rect 19475 3145 19484 3179
rect 19432 3136 19484 3145
rect 19616 3136 19668 3188
rect 20444 3136 20496 3188
rect 20720 3136 20772 3188
rect 20076 3068 20128 3120
rect 16396 3000 16448 3052
rect 17132 3000 17184 3052
rect 17500 3000 17552 3052
rect 13544 2932 13596 2984
rect 15108 2932 15160 2984
rect 15384 2932 15436 2984
rect 16764 2975 16816 2984
rect 16764 2941 16773 2975
rect 16773 2941 16807 2975
rect 16807 2941 16816 2975
rect 16764 2932 16816 2941
rect 16856 2975 16908 2984
rect 16856 2941 16865 2975
rect 16865 2941 16899 2975
rect 16899 2941 16908 2975
rect 17408 2975 17460 2984
rect 16856 2932 16908 2941
rect 17408 2941 17417 2975
rect 17417 2941 17451 2975
rect 17451 2941 17460 2975
rect 17408 2932 17460 2941
rect 4160 2907 4212 2916
rect 4160 2873 4194 2907
rect 4194 2873 4212 2907
rect 6092 2907 6144 2916
rect 4160 2864 4212 2873
rect 6092 2873 6101 2907
rect 6101 2873 6135 2907
rect 6135 2873 6144 2907
rect 6092 2864 6144 2873
rect 7196 2864 7248 2916
rect 2044 2796 2096 2848
rect 2780 2796 2832 2848
rect 3148 2839 3200 2848
rect 3148 2805 3157 2839
rect 3157 2805 3191 2839
rect 3191 2805 3200 2839
rect 3148 2796 3200 2805
rect 4252 2796 4304 2848
rect 5356 2796 5408 2848
rect 6920 2796 6972 2848
rect 8392 2796 8444 2848
rect 9588 2864 9640 2916
rect 9864 2864 9916 2916
rect 11244 2864 11296 2916
rect 8760 2796 8812 2848
rect 9312 2796 9364 2848
rect 10048 2796 10100 2848
rect 10232 2796 10284 2848
rect 18328 2864 18380 2916
rect 18604 2907 18656 2916
rect 18604 2873 18613 2907
rect 18613 2873 18647 2907
rect 18647 2873 18656 2907
rect 18604 2864 18656 2873
rect 11428 2796 11480 2848
rect 11980 2796 12032 2848
rect 18420 2796 18472 2848
rect 18696 2839 18748 2848
rect 18696 2805 18705 2839
rect 18705 2805 18739 2839
rect 18739 2805 18748 2839
rect 18696 2796 18748 2805
rect 18972 3000 19024 3052
rect 19800 3000 19852 3052
rect 19248 2932 19300 2984
rect 19340 2932 19392 2984
rect 20444 2975 20496 2984
rect 20444 2941 20453 2975
rect 20453 2941 20487 2975
rect 20487 2941 20496 2975
rect 20444 2932 20496 2941
rect 22560 2932 22612 2984
rect 20536 2864 20588 2916
rect 20628 2864 20680 2916
rect 22192 2864 22244 2916
rect 19248 2796 19300 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 1400 2592 1452 2644
rect 2136 2592 2188 2644
rect 3148 2592 3200 2644
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 4712 2592 4764 2644
rect 5632 2592 5684 2644
rect 6552 2592 6604 2644
rect 6920 2635 6972 2644
rect 6920 2601 6929 2635
rect 6929 2601 6963 2635
rect 6963 2601 6972 2635
rect 6920 2592 6972 2601
rect 7196 2592 7248 2644
rect 1860 2524 1912 2576
rect 1952 2456 2004 2508
rect 3240 2524 3292 2576
rect 7656 2524 7708 2576
rect 8116 2524 8168 2576
rect 8484 2524 8536 2576
rect 9312 2524 9364 2576
rect 3792 2456 3844 2508
rect 4160 2456 4212 2508
rect 5080 2456 5132 2508
rect 5816 2456 5868 2508
rect 8208 2456 8260 2508
rect 8392 2499 8444 2508
rect 8392 2465 8401 2499
rect 8401 2465 8435 2499
rect 8435 2465 8444 2499
rect 8392 2456 8444 2465
rect 2688 2388 2740 2440
rect 3424 2431 3476 2440
rect 3424 2397 3433 2431
rect 3433 2397 3467 2431
rect 3467 2397 3476 2431
rect 3424 2388 3476 2397
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 8852 2456 8904 2508
rect 9128 2499 9180 2508
rect 9128 2465 9137 2499
rect 9137 2465 9171 2499
rect 9171 2465 9180 2499
rect 9128 2456 9180 2465
rect 9956 2456 10008 2508
rect 6368 2388 6420 2397
rect 8668 2388 8720 2440
rect 8300 2320 8352 2372
rect 11060 2592 11112 2644
rect 14280 2592 14332 2644
rect 12256 2524 12308 2576
rect 13176 2524 13228 2576
rect 13360 2524 13412 2576
rect 10968 2456 11020 2508
rect 11336 2456 11388 2508
rect 11796 2499 11848 2508
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 13452 2456 13504 2508
rect 13912 2456 13964 2508
rect 11704 2388 11756 2440
rect 14096 2524 14148 2576
rect 16304 2592 16356 2644
rect 16672 2635 16724 2644
rect 16672 2601 16681 2635
rect 16681 2601 16715 2635
rect 16715 2601 16724 2635
rect 16672 2592 16724 2601
rect 17132 2592 17184 2644
rect 17500 2592 17552 2644
rect 17684 2592 17736 2644
rect 17868 2592 17920 2644
rect 18236 2592 18288 2644
rect 19156 2592 19208 2644
rect 19524 2592 19576 2644
rect 19708 2635 19760 2644
rect 19708 2601 19717 2635
rect 19717 2601 19751 2635
rect 19751 2601 19760 2635
rect 19708 2592 19760 2601
rect 14740 2499 14792 2508
rect 14740 2465 14749 2499
rect 14749 2465 14783 2499
rect 14783 2465 14792 2499
rect 14740 2456 14792 2465
rect 14832 2499 14884 2508
rect 14832 2465 14841 2499
rect 14841 2465 14875 2499
rect 14875 2465 14884 2499
rect 14832 2456 14884 2465
rect 15292 2456 15344 2508
rect 19064 2524 19116 2576
rect 19248 2524 19300 2576
rect 20628 2567 20680 2576
rect 20628 2533 20637 2567
rect 20637 2533 20671 2567
rect 20671 2533 20680 2567
rect 20628 2524 20680 2533
rect 16488 2388 16540 2440
rect 17868 2431 17920 2440
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 3424 2252 3476 2304
rect 4804 2252 4856 2304
rect 5908 2252 5960 2304
rect 9128 2252 9180 2304
rect 9680 2252 9732 2304
rect 10784 2295 10836 2304
rect 10784 2261 10793 2295
rect 10793 2261 10827 2295
rect 10827 2261 10836 2295
rect 10784 2252 10836 2261
rect 12716 2252 12768 2304
rect 17224 2295 17276 2304
rect 17224 2261 17233 2295
rect 17233 2261 17267 2295
rect 17267 2261 17276 2295
rect 17224 2252 17276 2261
rect 17316 2252 17368 2304
rect 20076 2456 20128 2508
rect 18972 2431 19024 2440
rect 18972 2397 18981 2431
rect 18981 2397 19015 2431
rect 19015 2397 19024 2431
rect 18972 2388 19024 2397
rect 19892 2431 19944 2440
rect 19892 2397 19901 2431
rect 19901 2397 19935 2431
rect 19935 2397 19944 2431
rect 19892 2388 19944 2397
rect 18328 2320 18380 2372
rect 21456 2320 21508 2372
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 5080 2048 5132 2100
rect 9956 2048 10008 2100
rect 10784 2048 10836 2100
rect 204 1980 256 2032
rect 8392 1980 8444 2032
rect 2044 1912 2096 1964
rect 7196 1912 7248 1964
rect 14740 2048 14792 2100
rect 20904 2048 20956 2100
rect 14280 1980 14332 2032
rect 18972 1980 19024 2032
rect 20260 1912 20312 1964
rect 1308 1844 1360 1896
rect 7564 1844 7616 1896
rect 7748 1844 7800 1896
rect 14832 1844 14884 1896
rect 15476 1844 15528 1896
rect 17408 1844 17460 1896
rect 5356 1776 5408 1828
rect 7380 1776 7432 1828
rect 17316 1776 17368 1828
rect 572 1708 624 1760
rect 8116 1708 8168 1760
rect 12992 1708 13044 1760
rect 15476 1708 15528 1760
rect 2412 1640 2464 1692
rect 7104 1640 7156 1692
rect 2780 1572 2832 1624
rect 6828 1572 6880 1624
rect 9680 1368 9732 1420
rect 15108 1368 15160 1420
rect 16764 1300 16816 1352
rect 17960 1300 18012 1352
rect 12808 1232 12860 1284
rect 14372 1232 14424 1284
rect 16580 1096 16632 1148
rect 17132 1096 17184 1148
<< metal2 >>
rect 202 22320 258 22800
rect 570 22320 626 22800
rect 938 22320 994 22800
rect 1306 22320 1362 22800
rect 1674 22320 1730 22800
rect 2042 22320 2098 22800
rect 2410 22320 2466 22800
rect 2778 22320 2834 22800
rect 3238 22320 3294 22800
rect 3606 22320 3662 22800
rect 3974 22320 4030 22800
rect 4342 22320 4398 22800
rect 4710 22320 4766 22800
rect 5078 22320 5134 22800
rect 5446 22320 5502 22800
rect 5906 22320 5962 22800
rect 6274 22320 6330 22800
rect 6642 22320 6698 22800
rect 7010 22320 7066 22800
rect 7378 22320 7434 22800
rect 7746 22320 7802 22800
rect 8114 22320 8170 22800
rect 8482 22320 8538 22800
rect 8942 22320 8998 22800
rect 9310 22320 9366 22800
rect 9678 22320 9734 22800
rect 10046 22320 10102 22800
rect 10414 22320 10470 22800
rect 10782 22320 10838 22800
rect 11150 22320 11206 22800
rect 11610 22320 11666 22800
rect 11978 22320 12034 22800
rect 12346 22320 12402 22800
rect 12714 22320 12770 22800
rect 13082 22320 13138 22800
rect 13450 22320 13506 22800
rect 13818 22320 13874 22800
rect 14186 22320 14242 22800
rect 14646 22320 14702 22800
rect 15014 22320 15070 22800
rect 15382 22320 15438 22800
rect 15750 22320 15806 22800
rect 16118 22320 16174 22800
rect 16486 22320 16542 22800
rect 16854 22320 16910 22800
rect 17314 22320 17370 22800
rect 17682 22320 17738 22800
rect 18050 22320 18106 22800
rect 18418 22320 18474 22800
rect 18786 22320 18842 22800
rect 19154 22320 19210 22800
rect 19522 22320 19578 22800
rect 19890 22320 19946 22800
rect 20350 22320 20406 22800
rect 20718 22320 20774 22800
rect 20810 22672 20866 22681
rect 20810 22607 20866 22616
rect 216 17882 244 22320
rect 584 20330 612 22320
rect 572 20324 624 20330
rect 572 20266 624 20272
rect 204 17876 256 17882
rect 204 17818 256 17824
rect 952 17746 980 22320
rect 1320 19242 1348 22320
rect 1688 19786 1716 22320
rect 1950 21040 2006 21049
rect 1950 20975 2006 20984
rect 1858 20632 1914 20641
rect 1858 20567 1914 20576
rect 1676 19780 1728 19786
rect 1676 19722 1728 19728
rect 1872 19310 1900 20567
rect 1964 19990 1992 20975
rect 1952 19984 2004 19990
rect 1952 19926 2004 19932
rect 1950 19408 2006 19417
rect 1950 19343 2006 19352
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 1308 19236 1360 19242
rect 1308 19178 1360 19184
rect 1688 18057 1716 19246
rect 1964 18902 1992 19343
rect 2056 19310 2084 22320
rect 2318 19952 2374 19961
rect 2318 19887 2320 19896
rect 2372 19887 2374 19896
rect 2320 19858 2372 19864
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 2424 19258 2452 22320
rect 2792 19938 2820 22320
rect 2792 19910 3096 19938
rect 2780 19848 2832 19854
rect 2778 19816 2780 19825
rect 2832 19816 2834 19825
rect 2778 19751 2834 19760
rect 2424 19230 3004 19258
rect 2976 19174 3004 19230
rect 2780 19168 2832 19174
rect 2964 19168 3016 19174
rect 2832 19128 2912 19156
rect 2780 19110 2832 19116
rect 1952 18896 2004 18902
rect 1952 18838 2004 18844
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2228 18760 2280 18766
rect 1950 18728 2006 18737
rect 2228 18702 2280 18708
rect 1950 18663 2006 18672
rect 1964 18426 1992 18663
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 2240 18290 2268 18702
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 1674 18048 1730 18057
rect 1674 17983 1730 17992
rect 1490 17912 1546 17921
rect 1490 17847 1546 17856
rect 1860 17876 1912 17882
rect 940 17740 992 17746
rect 940 17682 992 17688
rect 1504 16250 1532 17847
rect 1860 17818 1912 17824
rect 1872 17785 1900 17818
rect 1858 17776 1914 17785
rect 1768 17740 1820 17746
rect 1858 17711 1914 17720
rect 1768 17682 1820 17688
rect 1780 17649 1808 17682
rect 1766 17640 1822 17649
rect 1766 17575 1822 17584
rect 2044 17332 2096 17338
rect 2044 17274 2096 17280
rect 1582 17096 1638 17105
rect 1582 17031 1638 17040
rect 1676 17060 1728 17066
rect 1492 16244 1544 16250
rect 1492 16186 1544 16192
rect 1492 16040 1544 16046
rect 1492 15982 1544 15988
rect 1400 15972 1452 15978
rect 1400 15914 1452 15920
rect 1412 15570 1440 15914
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1504 12889 1532 15982
rect 1596 15706 1624 17031
rect 1676 17002 1728 17008
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1582 14376 1638 14385
rect 1582 14311 1638 14320
rect 1596 14074 1624 14311
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1688 13870 1716 17002
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1780 16794 1808 16934
rect 2056 16794 2084 17274
rect 2240 17066 2268 18226
rect 2228 17060 2280 17066
rect 2228 17002 2280 17008
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1584 13796 1636 13802
rect 1584 13738 1636 13744
rect 1596 12986 1624 13738
rect 1674 13560 1730 13569
rect 1674 13495 1730 13504
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1490 12880 1546 12889
rect 1490 12815 1546 12824
rect 1492 12368 1544 12374
rect 1492 12310 1544 12316
rect 1400 11620 1452 11626
rect 1400 11562 1452 11568
rect 1412 9042 1440 11562
rect 1504 11354 1532 12310
rect 1492 11348 1544 11354
rect 1492 11290 1544 11296
rect 1582 11248 1638 11257
rect 1582 11183 1638 11192
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 7002 1440 8230
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1596 6458 1624 11183
rect 1688 10266 1716 13495
rect 1780 12306 1808 15438
rect 1768 12300 1820 12306
rect 1768 12242 1820 12248
rect 1780 10810 1808 12242
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1872 10577 1900 16594
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 2044 14884 2096 14890
rect 2044 14826 2096 14832
rect 2056 14414 2084 14826
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 2044 13728 2096 13734
rect 2044 13670 2096 13676
rect 1964 12753 1992 13670
rect 2056 13530 2084 13670
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 1950 12744 2006 12753
rect 1950 12679 2006 12688
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1858 10568 1914 10577
rect 1858 10503 1914 10512
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1872 10130 1900 10503
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1872 9353 1900 9454
rect 1858 9344 1914 9353
rect 1858 9279 1914 9288
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1674 7440 1730 7449
rect 1674 7375 1730 7384
rect 1688 6866 1716 7375
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1596 5234 1624 6190
rect 1780 5914 1808 8298
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1872 7342 1900 7686
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1872 6254 1900 7278
rect 1964 6458 1992 12174
rect 2056 9217 2084 13466
rect 2148 12238 2176 15982
rect 2240 14890 2268 17002
rect 2332 16046 2360 18770
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2412 17060 2464 17066
rect 2412 17002 2464 17008
rect 2424 16522 2452 17002
rect 2412 16516 2464 16522
rect 2412 16458 2464 16464
rect 2410 16144 2466 16153
rect 2410 16079 2466 16088
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2424 15706 2452 16079
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2516 15586 2544 17614
rect 2608 16794 2636 17682
rect 2792 17513 2820 18566
rect 2884 17882 2912 19128
rect 2964 19110 3016 19116
rect 2964 18148 3016 18154
rect 2964 18090 3016 18096
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2976 17678 3004 18090
rect 3068 17882 3096 19910
rect 3252 18329 3280 22320
rect 3516 19916 3568 19922
rect 3516 19858 3568 19864
rect 3528 19378 3556 19858
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3528 19174 3556 19314
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3238 18320 3294 18329
rect 3238 18255 3294 18264
rect 3146 18184 3202 18193
rect 3330 18184 3386 18193
rect 3146 18119 3202 18128
rect 3252 18142 3330 18170
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2778 17504 2834 17513
rect 2778 17439 2834 17448
rect 2780 17332 2832 17338
rect 2976 17320 3004 17614
rect 3160 17542 3188 18119
rect 3252 17882 3280 18142
rect 3330 18119 3386 18128
rect 3436 17882 3464 18702
rect 3516 18692 3568 18698
rect 3516 18634 3568 18640
rect 3528 18290 3556 18634
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3620 18057 3648 22320
rect 3882 22264 3938 22273
rect 3882 22199 3938 22208
rect 3698 21856 3754 21865
rect 3698 21791 3754 21800
rect 3712 18068 3740 21791
rect 3896 21282 3924 22199
rect 3884 21276 3936 21282
rect 3884 21218 3936 21224
rect 3792 20664 3844 20670
rect 3792 20606 3844 20612
rect 3804 19786 3832 20606
rect 3882 20224 3938 20233
rect 3882 20159 3938 20168
rect 3792 19780 3844 19786
rect 3792 19722 3844 19728
rect 3792 19168 3844 19174
rect 3792 19110 3844 19116
rect 3804 18222 3832 19110
rect 3896 18873 3924 20159
rect 3882 18864 3938 18873
rect 3882 18799 3938 18808
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3606 18048 3662 18057
rect 3712 18040 3924 18068
rect 3606 17983 3662 17992
rect 3240 17876 3292 17882
rect 3240 17818 3292 17824
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3056 17332 3108 17338
rect 2976 17292 3056 17320
rect 2780 17274 2832 17280
rect 3056 17274 3108 17280
rect 2792 17105 2820 17274
rect 2872 17128 2924 17134
rect 2778 17096 2834 17105
rect 2872 17070 2924 17076
rect 2778 17031 2834 17040
rect 2596 16788 2648 16794
rect 2596 16730 2648 16736
rect 2780 16720 2832 16726
rect 2780 16662 2832 16668
rect 2792 16538 2820 16662
rect 2700 16510 2820 16538
rect 2594 15600 2650 15609
rect 2516 15558 2594 15586
rect 2594 15535 2650 15544
rect 2608 15502 2636 15535
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2228 14884 2280 14890
rect 2228 14826 2280 14832
rect 2700 14385 2728 16510
rect 2778 16280 2834 16289
rect 2778 16215 2834 16224
rect 2686 14376 2742 14385
rect 2686 14311 2742 14320
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2332 12782 2360 13262
rect 2424 12850 2452 13330
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2042 9208 2098 9217
rect 2042 9143 2098 9152
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2056 7342 2084 8434
rect 2044 7336 2096 7342
rect 2044 7278 2096 7284
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1872 5574 1900 6190
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 940 3732 992 3738
rect 940 3674 992 3680
rect 204 2032 256 2038
rect 204 1974 256 1980
rect 216 480 244 1974
rect 572 1760 624 1766
rect 572 1702 624 1708
rect 584 480 612 1702
rect 952 480 980 3674
rect 1412 2650 1440 5102
rect 1872 4486 1900 5510
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1872 4026 1900 4422
rect 1872 3998 1992 4026
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1504 2990 1532 3470
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1676 2916 1728 2922
rect 1676 2858 1728 2864
rect 1400 2644 1452 2650
rect 1400 2586 1452 2592
rect 1308 1896 1360 1902
rect 1308 1838 1360 1844
rect 1320 480 1348 1838
rect 1688 480 1716 2858
rect 1872 2582 1900 3878
rect 1964 3534 1992 3998
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1860 2576 1912 2582
rect 1860 2518 1912 2524
rect 1964 2514 1992 3470
rect 2056 2854 2084 7142
rect 2148 7018 2176 12038
rect 2608 11694 2636 12718
rect 2792 12442 2820 16215
rect 2884 14618 2912 17070
rect 3252 16726 3280 17818
rect 3424 17740 3476 17746
rect 3424 17682 3476 17688
rect 3436 17241 3464 17682
rect 3422 17232 3478 17241
rect 3422 17167 3478 17176
rect 3896 17134 3924 18040
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3988 16969 4016 22320
rect 4356 22250 4384 22320
rect 4172 22222 4384 22250
rect 4066 21448 4122 21457
rect 4066 21383 4122 21392
rect 4080 21010 4108 21383
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4080 19514 4108 19654
rect 4068 19508 4120 19514
rect 4172 19496 4200 22222
rect 4724 20890 4752 22320
rect 4724 20862 4844 20890
rect 4710 19816 4766 19825
rect 4710 19751 4766 19760
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4172 19468 4476 19496
rect 4068 19450 4120 19456
rect 4066 19408 4122 19417
rect 4066 19343 4122 19352
rect 4252 19372 4304 19378
rect 4080 19310 4108 19343
rect 4252 19314 4304 19320
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4172 18834 4200 19246
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 4264 17320 4292 19314
rect 4448 19281 4476 19468
rect 4434 19272 4490 19281
rect 4344 19236 4396 19242
rect 4434 19207 4490 19216
rect 4344 19178 4396 19184
rect 4356 19145 4384 19178
rect 4342 19136 4398 19145
rect 4342 19071 4398 19080
rect 4724 18970 4752 19751
rect 4816 18970 4844 20862
rect 4988 20460 5040 20466
rect 4988 20402 5040 20408
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 4908 19174 4936 19858
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4436 18352 4488 18358
rect 4434 18320 4436 18329
rect 4488 18320 4490 18329
rect 4434 18255 4490 18264
rect 4712 18284 4764 18290
rect 4712 18226 4764 18232
rect 4344 18216 4396 18222
rect 4396 18176 4476 18204
rect 4344 18158 4396 18164
rect 4448 18086 4476 18176
rect 4528 18148 4580 18154
rect 4528 18090 4580 18096
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4356 17882 4384 18022
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4540 17678 4568 18090
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4264 17292 4568 17320
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 3974 16960 4030 16969
rect 3974 16895 4030 16904
rect 3988 16782 4200 16810
rect 3988 16726 4016 16782
rect 3240 16720 3292 16726
rect 3240 16662 3292 16668
rect 3976 16720 4028 16726
rect 3976 16662 4028 16668
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 3344 16114 3372 16526
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3252 15745 3280 15846
rect 3238 15736 3294 15745
rect 3238 15671 3294 15680
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2884 13841 2912 13942
rect 2870 13832 2926 13841
rect 2870 13767 2926 13776
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2976 13462 3004 13670
rect 2964 13456 3016 13462
rect 2964 13398 3016 13404
rect 2870 13152 2926 13161
rect 2870 13087 2926 13096
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2332 10010 2360 11494
rect 2608 11286 2636 11630
rect 2596 11280 2648 11286
rect 2596 11222 2648 11228
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2596 10532 2648 10538
rect 2596 10474 2648 10480
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2240 9982 2360 10010
rect 2240 9178 2268 9982
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2332 9110 2360 9862
rect 2516 9722 2544 10066
rect 2608 10062 2636 10474
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2608 9602 2636 9998
rect 2424 9586 2636 9602
rect 2412 9580 2636 9586
rect 2464 9574 2636 9580
rect 2412 9522 2464 9528
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2424 9178 2452 9318
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2424 7206 2452 8978
rect 2516 8634 2544 9318
rect 2608 9178 2636 9386
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2700 8974 2728 11154
rect 2792 10538 2820 12174
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2884 10266 2912 13087
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2976 12442 3004 12582
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 3054 12336 3110 12345
rect 2964 12300 3016 12306
rect 3054 12271 3110 12280
rect 2964 12242 3016 12248
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2780 10192 2832 10198
rect 2976 10146 3004 12242
rect 2780 10134 2832 10140
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2792 8838 2820 10134
rect 2884 10118 3004 10146
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2884 8498 2912 10118
rect 3068 9654 3096 12271
rect 3252 12170 3280 15506
rect 3330 14920 3386 14929
rect 3330 14855 3386 14864
rect 3344 14006 3372 14855
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 3436 13530 3464 16594
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 3514 16008 3570 16017
rect 3514 15943 3570 15952
rect 3528 15706 3556 15943
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3608 15496 3660 15502
rect 3608 15438 3660 15444
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3528 14414 3556 14758
rect 3620 14482 3648 15438
rect 3792 15156 3844 15162
rect 3896 15144 3924 16458
rect 4172 16046 4200 16782
rect 4264 16114 4292 17138
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 4448 16794 4476 16934
rect 4540 16794 4568 17292
rect 4724 17202 4752 18226
rect 4816 18154 4844 18770
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4908 17134 4936 19110
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 4344 16720 4396 16726
rect 4342 16688 4344 16697
rect 4396 16688 4398 16697
rect 4342 16623 4398 16632
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4724 16250 4752 16934
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 4712 15972 4764 15978
rect 4712 15914 4764 15920
rect 4066 15872 4122 15881
rect 4066 15807 4122 15816
rect 4080 15706 4108 15807
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 3974 15464 4030 15473
rect 3974 15399 4030 15408
rect 4160 15428 4212 15434
rect 3844 15116 3924 15144
rect 3792 15098 3844 15104
rect 3790 14784 3846 14793
rect 3790 14719 3846 14728
rect 3608 14476 3660 14482
rect 3608 14418 3660 14424
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3240 12164 3292 12170
rect 3240 12106 3292 12112
rect 3252 12073 3280 12106
rect 3238 12064 3294 12073
rect 3238 11999 3294 12008
rect 3146 11928 3202 11937
rect 3146 11863 3202 11872
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 9042 3004 9318
rect 3054 9208 3110 9217
rect 3054 9143 3110 9152
rect 3068 9042 3096 9143
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2596 7948 2648 7954
rect 2596 7890 2648 7896
rect 2608 7562 2636 7890
rect 2608 7546 2728 7562
rect 2608 7540 2740 7546
rect 2608 7534 2688 7540
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2148 6990 2544 7018
rect 2226 6896 2282 6905
rect 2516 6866 2544 6990
rect 2226 6831 2282 6840
rect 2504 6860 2556 6866
rect 2240 6730 2268 6831
rect 2504 6802 2556 6808
rect 2608 6798 2636 7534
rect 2688 7482 2740 7488
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2412 6180 2464 6186
rect 2412 6122 2464 6128
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 2056 2553 2084 2790
rect 2148 2650 2176 4966
rect 2424 4826 2452 6122
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2410 3904 2466 3913
rect 2410 3839 2466 3848
rect 2424 3369 2452 3839
rect 2410 3360 2466 3369
rect 2410 3295 2466 3304
rect 2516 3194 2544 4966
rect 2608 3194 2636 4966
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2042 2544 2098 2553
rect 1952 2508 2004 2514
rect 2042 2479 2098 2488
rect 1952 2450 2004 2456
rect 2700 2446 2728 4762
rect 2884 4622 2912 8434
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 6662 3004 7890
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2976 4690 3004 5170
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2976 4146 3004 4626
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2884 3505 2912 3674
rect 2870 3496 2926 3505
rect 2870 3431 2926 3440
rect 2976 3398 3004 4082
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2792 2689 2820 2790
rect 2778 2680 2834 2689
rect 2778 2615 2834 2624
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 2044 1964 2096 1970
rect 2044 1906 2096 1912
rect 2056 480 2084 1906
rect 2792 1737 2820 2615
rect 2778 1728 2834 1737
rect 2412 1692 2464 1698
rect 2778 1663 2834 1672
rect 2412 1634 2464 1640
rect 2424 480 2452 1634
rect 2780 1624 2832 1630
rect 2780 1566 2832 1572
rect 2792 480 2820 1566
rect 3068 513 3096 8978
rect 3160 8906 3188 11863
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3252 11354 3280 11698
rect 3344 11354 3372 12242
rect 3528 12238 3556 12650
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3252 10810 3280 11018
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3252 10130 3280 10542
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3252 8922 3280 9522
rect 3344 9110 3372 10406
rect 3436 9364 3464 12174
rect 3620 11778 3648 14214
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 3712 13530 3740 13874
rect 3700 13524 3752 13530
rect 3700 13466 3752 13472
rect 3528 11750 3648 11778
rect 3528 9654 3556 11750
rect 3606 11656 3662 11665
rect 3606 11591 3662 11600
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3436 9336 3556 9364
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3252 8906 3372 8922
rect 3148 8900 3200 8906
rect 3252 8900 3384 8906
rect 3252 8894 3332 8900
rect 3148 8842 3200 8848
rect 3332 8842 3384 8848
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 8566 3280 8774
rect 3240 8560 3292 8566
rect 3146 8528 3202 8537
rect 3240 8502 3292 8508
rect 3146 8463 3202 8472
rect 3160 4185 3188 8463
rect 3252 5166 3280 8502
rect 3344 8498 3372 8842
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3436 8090 3464 8366
rect 3528 8362 3556 9336
rect 3620 8634 3648 11591
rect 3698 11520 3754 11529
rect 3698 11455 3754 11464
rect 3712 10849 3740 11455
rect 3698 10840 3754 10849
rect 3804 10810 3832 14719
rect 3896 13870 3924 15116
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3896 12782 3924 13806
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3882 12608 3938 12617
rect 3882 12543 3938 12552
rect 3896 11286 3924 12543
rect 3988 12442 4016 15399
rect 4160 15370 4212 15376
rect 4066 15192 4122 15201
rect 4066 15127 4122 15136
rect 4080 14278 4108 15127
rect 4172 14618 4200 15370
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4264 14550 4292 15302
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4172 13530 4200 14010
rect 4250 13968 4306 13977
rect 4250 13903 4306 13912
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4080 12918 4108 13262
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 3974 12200 4030 12209
rect 3974 12135 4030 12144
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 3988 10962 4016 12135
rect 4264 11626 4292 13903
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4448 12306 4476 12718
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4632 11626 4660 11766
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4080 11354 4108 11494
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 3896 10934 4016 10962
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 3698 10775 3754 10784
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3804 9500 3832 9590
rect 3712 9472 3832 9500
rect 3712 9382 3740 9472
rect 3896 9450 3924 10934
rect 3976 10532 4028 10538
rect 3976 10474 4028 10480
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3422 7848 3478 7857
rect 3422 7783 3478 7792
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 3344 6390 3372 7210
rect 3332 6384 3384 6390
rect 3332 6326 3384 6332
rect 3344 6225 3372 6326
rect 3330 6216 3386 6225
rect 3330 6151 3386 6160
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3344 5370 3372 6054
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3146 4176 3202 4185
rect 3146 4111 3202 4120
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3160 3534 3188 3946
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 3252 2961 3280 5102
rect 3436 4826 3464 7783
rect 3528 6610 3556 8298
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3620 6769 3648 6938
rect 3712 6934 3740 9318
rect 3988 9160 4016 10474
rect 4080 10441 4108 10950
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 3804 9132 4016 9160
rect 3804 7206 3832 9132
rect 4080 9092 4108 10066
rect 4172 9654 4200 11154
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4264 10810 4292 11086
rect 4724 11082 4752 15914
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4816 14958 4844 15438
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4816 14414 4844 14894
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 5000 14260 5028 20402
rect 5092 18986 5120 22320
rect 5356 20324 5408 20330
rect 5356 20266 5408 20272
rect 5368 19922 5396 20266
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5172 19780 5224 19786
rect 5172 19722 5224 19728
rect 5184 19174 5212 19722
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5170 19000 5226 19009
rect 5092 18958 5170 18986
rect 5170 18935 5226 18944
rect 5080 18896 5132 18902
rect 5080 18838 5132 18844
rect 5092 17882 5120 18838
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 5184 16590 5212 18702
rect 5276 17785 5304 19790
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 5368 19310 5396 19722
rect 5356 19304 5408 19310
rect 5356 19246 5408 19252
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5368 18748 5396 19110
rect 5460 18816 5488 22320
rect 5538 19408 5594 19417
rect 5538 19343 5594 19352
rect 5552 18884 5580 19343
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5724 18896 5776 18902
rect 5552 18856 5724 18884
rect 5724 18838 5776 18844
rect 5460 18788 5672 18816
rect 5368 18720 5580 18748
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5368 18222 5396 18566
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5262 17776 5318 17785
rect 5262 17711 5318 17720
rect 5276 17202 5304 17711
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5368 16658 5396 18022
rect 5552 17796 5580 18720
rect 5644 18306 5672 18788
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5736 18426 5764 18566
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5644 18278 5764 18306
rect 5552 17768 5672 17796
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5184 16114 5212 16526
rect 5368 16250 5396 16594
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5460 16182 5488 17682
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5552 17338 5580 17614
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5644 17218 5672 17768
rect 5552 17190 5672 17218
rect 5552 16658 5580 17190
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5262 16008 5318 16017
rect 5552 15994 5580 16594
rect 5644 16114 5672 16934
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5552 15966 5672 15994
rect 5262 15943 5318 15952
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 15366 5212 15846
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5092 14346 5120 14894
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 4816 14232 5028 14260
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 4264 9586 4292 10134
rect 4356 9908 4384 10678
rect 4325 9880 4384 9908
rect 4325 9704 4353 9880
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4325 9676 4384 9704
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4160 9104 4212 9110
rect 3988 9064 4160 9092
rect 3988 8498 4016 9064
rect 4160 9046 4212 9052
rect 4356 8820 4384 9676
rect 4710 9480 4766 9489
rect 4710 9415 4766 9424
rect 4724 9178 4752 9415
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4264 8792 4384 8820
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3988 7750 4016 8434
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4264 8344 4292 8792
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4710 8392 4766 8401
rect 4344 8356 4396 8362
rect 4264 8316 4344 8344
rect 4172 7818 4200 8298
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 3976 7744 4028 7750
rect 4068 7744 4120 7750
rect 3976 7686 4028 7692
rect 4066 7712 4068 7721
rect 4120 7712 4122 7721
rect 4264 7698 4292 8316
rect 4710 8327 4712 8336
rect 4344 8298 4396 8304
rect 4764 8327 4766 8336
rect 4712 8298 4764 8304
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 3884 7336 3936 7342
rect 3988 7324 4016 7686
rect 4066 7647 4122 7656
rect 4172 7670 4292 7698
rect 3936 7296 4016 7324
rect 3884 7278 3936 7284
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3700 6928 3752 6934
rect 3700 6870 3752 6876
rect 3606 6760 3662 6769
rect 3606 6695 3662 6704
rect 3528 6582 3648 6610
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3528 5574 3556 6258
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3436 4282 3464 4626
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3344 3738 3372 3878
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3436 3618 3464 4082
rect 3344 3602 3464 3618
rect 3332 3596 3464 3602
rect 3384 3590 3464 3596
rect 3332 3538 3384 3544
rect 3344 3194 3372 3538
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3344 3058 3372 3130
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3238 2952 3294 2961
rect 3238 2887 3294 2896
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 3160 2650 3188 2790
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 3252 1306 3280 2518
rect 3160 1278 3280 1306
rect 3054 504 3110 513
rect 202 0 258 480
rect 570 0 626 480
rect 938 0 994 480
rect 1306 0 1362 480
rect 1674 0 1730 480
rect 2042 0 2098 480
rect 2410 0 2466 480
rect 2778 0 2834 480
rect 3160 480 3188 1278
rect 3344 921 3372 2586
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3436 2310 3464 2382
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3330 912 3386 921
rect 3330 847 3386 856
rect 3054 439 3110 448
rect 3146 0 3202 480
rect 3436 241 3464 2246
rect 3528 480 3556 5510
rect 3620 2689 3648 6582
rect 3606 2680 3662 2689
rect 3606 2615 3662 2624
rect 3712 2145 3740 6870
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3988 5234 4016 5850
rect 4172 5692 4200 7670
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4724 7546 4752 7822
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4264 5846 4292 6802
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4618 6352 4674 6361
rect 4618 6287 4620 6296
rect 4672 6287 4674 6296
rect 4620 6258 4672 6264
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 4066 5672 4122 5681
rect 4172 5664 4292 5692
rect 4066 5607 4122 5616
rect 4080 5574 4108 5607
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4068 5024 4120 5030
rect 3974 4992 4030 5001
rect 4068 4966 4120 4972
rect 3974 4927 4030 4936
rect 3988 4706 4016 4927
rect 4080 4826 4108 4966
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 3988 4678 4108 4706
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 3882 2952 3938 2961
rect 3804 2514 3832 2926
rect 3882 2887 3938 2896
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3698 2136 3754 2145
rect 3698 2071 3754 2080
rect 3896 480 3924 2887
rect 3988 1329 4016 4558
rect 4080 4049 4108 4678
rect 4066 4040 4122 4049
rect 4066 3975 4122 3984
rect 4264 3942 4292 5664
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4632 4622 4660 5170
rect 4724 5114 4752 7210
rect 4816 6254 4844 14232
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4894 13016 4950 13025
rect 4894 12951 4950 12960
rect 4908 12782 4936 12951
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 4896 11824 4948 11830
rect 5000 11812 5028 12242
rect 4948 11784 5028 11812
rect 4896 11766 4948 11772
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4894 10840 4950 10849
rect 4894 10775 4950 10784
rect 4908 9042 4936 10775
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4908 7274 4936 8978
rect 4896 7268 4948 7274
rect 4896 7210 4948 7216
rect 4896 6384 4948 6390
rect 4894 6352 4896 6361
rect 4948 6352 4950 6361
rect 4894 6287 4950 6296
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4724 5086 4844 5114
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4724 4282 4752 4966
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4448 4049 4476 4082
rect 4712 4072 4764 4078
rect 4434 4040 4490 4049
rect 4712 4014 4764 4020
rect 4434 3975 4490 3984
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4172 3602 4200 3878
rect 4250 3768 4306 3777
rect 4250 3703 4252 3712
rect 4304 3703 4306 3712
rect 4252 3674 4304 3680
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4264 3534 4292 3674
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4448 3380 4476 3975
rect 4724 3738 4752 4014
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4448 3352 4752 3380
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4724 3176 4752 3352
rect 4632 3148 4752 3176
rect 4160 2916 4212 2922
rect 4160 2858 4212 2864
rect 4172 2514 4200 2858
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 3974 1320 4030 1329
rect 3974 1255 4030 1264
rect 4264 480 4292 2790
rect 4632 2292 4660 3148
rect 4816 3074 4844 5086
rect 4724 3046 4844 3074
rect 4724 2650 4752 3046
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4804 2304 4856 2310
rect 4632 2264 4752 2292
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4724 2088 4752 2264
rect 4908 2292 4936 6190
rect 4856 2264 4936 2292
rect 4804 2246 4856 2252
rect 4632 2060 4752 2088
rect 4632 480 4660 2060
rect 5000 480 5028 11630
rect 5092 11218 5120 13126
rect 5184 12617 5212 15302
rect 5170 12608 5226 12617
rect 5170 12543 5226 12552
rect 5170 12336 5226 12345
rect 5170 12271 5226 12280
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 5078 11112 5134 11121
rect 5078 11047 5134 11056
rect 5092 8945 5120 11047
rect 5184 9081 5212 12271
rect 5276 10985 5304 15943
rect 5644 15609 5672 15966
rect 5736 15706 5764 18278
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5630 15600 5686 15609
rect 5540 15564 5592 15570
rect 5630 15535 5686 15544
rect 5724 15564 5776 15570
rect 5540 15506 5592 15512
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5368 14074 5396 14826
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5460 14657 5488 14758
rect 5446 14648 5502 14657
rect 5446 14583 5502 14592
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5460 13802 5488 14214
rect 5552 14074 5580 15506
rect 5644 15042 5672 15535
rect 5724 15506 5776 15512
rect 5736 15162 5764 15506
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5644 15014 5764 15042
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5644 14550 5672 14894
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5630 14376 5686 14385
rect 5630 14311 5686 14320
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5644 13954 5672 14311
rect 5552 13926 5672 13954
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5460 12986 5488 13330
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5262 10976 5318 10985
rect 5262 10911 5318 10920
rect 5460 10826 5488 12650
rect 5368 10798 5488 10826
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5276 9994 5304 10678
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5276 9654 5304 9930
rect 5264 9648 5316 9654
rect 5264 9590 5316 9596
rect 5264 9376 5316 9382
rect 5368 9364 5396 10798
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5460 9926 5488 10610
rect 5552 10010 5580 13926
rect 5630 13560 5686 13569
rect 5630 13495 5632 13504
rect 5684 13495 5686 13504
rect 5632 13466 5684 13472
rect 5736 13433 5764 15014
rect 5722 13424 5778 13433
rect 5722 13359 5778 13368
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5644 11898 5672 13262
rect 5736 12850 5764 13262
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5736 12442 5764 12786
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5828 11354 5856 18906
rect 5920 18630 5948 22320
rect 6000 21004 6052 21010
rect 6000 20946 6052 20952
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 6012 18426 6040 20946
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6104 19825 6132 19858
rect 6090 19816 6146 19825
rect 6090 19751 6146 19760
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 6196 18970 6224 19654
rect 6288 19360 6316 22320
rect 6656 20210 6684 22320
rect 6564 20182 6684 20210
rect 6288 19332 6500 19360
rect 6472 19292 6500 19332
rect 6380 19264 6500 19292
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6104 17649 6132 18770
rect 6288 18766 6316 19110
rect 6276 18760 6328 18766
rect 6276 18702 6328 18708
rect 6380 18442 6408 19264
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6472 18601 6500 19110
rect 6458 18592 6514 18601
rect 6458 18527 6514 18536
rect 6288 18414 6408 18442
rect 6288 18034 6316 18414
rect 6460 18080 6512 18086
rect 6288 18006 6408 18034
rect 6460 18022 6512 18028
rect 6090 17640 6146 17649
rect 6090 17575 6092 17584
rect 6144 17575 6146 17584
rect 6092 17546 6144 17552
rect 6104 17515 6132 17546
rect 6090 17096 6146 17105
rect 6090 17031 6146 17040
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6012 16250 6040 16662
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6104 15892 6132 17031
rect 6276 16516 6328 16522
rect 6276 16458 6328 16464
rect 6288 16046 6316 16458
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6104 15864 6316 15892
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6092 15632 6144 15638
rect 6092 15574 6144 15580
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5920 14822 5948 15438
rect 6104 15094 6132 15574
rect 6092 15088 6144 15094
rect 6092 15030 6144 15036
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5920 14618 5948 14758
rect 6090 14648 6146 14657
rect 5908 14612 5960 14618
rect 6090 14583 6146 14592
rect 5908 14554 5960 14560
rect 5920 13938 5948 14554
rect 6104 14550 6132 14583
rect 6092 14544 6144 14550
rect 6092 14486 6144 14492
rect 6090 14376 6146 14385
rect 6090 14311 6146 14320
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5920 13190 5948 13738
rect 5998 13560 6054 13569
rect 5998 13495 6054 13504
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5920 12170 5948 12582
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 5906 11792 5962 11801
rect 5906 11727 5962 11736
rect 5920 11694 5948 11727
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5644 10130 5672 11086
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5736 10538 5764 11018
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5920 10577 5948 10610
rect 5906 10568 5962 10577
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5828 10526 5906 10554
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5722 10024 5778 10033
rect 5552 9982 5672 10010
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5460 9586 5488 9862
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5552 9518 5580 9862
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5644 9382 5672 9982
rect 5722 9959 5778 9968
rect 5736 9722 5764 9959
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 5316 9336 5396 9364
rect 5632 9376 5684 9382
rect 5264 9318 5316 9324
rect 5632 9318 5684 9324
rect 5170 9072 5226 9081
rect 5170 9007 5226 9016
rect 5078 8936 5134 8945
rect 5078 8871 5134 8880
rect 5092 6644 5120 8871
rect 5184 8401 5212 9007
rect 5170 8392 5226 8401
rect 5170 8327 5226 8336
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7546 5212 8230
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5184 7410 5212 7482
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5184 6798 5212 7346
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5092 6616 5212 6644
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5092 5778 5120 6394
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 5092 5234 5120 5714
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5092 3482 5120 4082
rect 5184 4010 5212 6616
rect 5276 6254 5304 9318
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5368 8634 5396 8978
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5354 8528 5410 8537
rect 5354 8463 5410 8472
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5262 6080 5318 6089
rect 5262 6015 5318 6024
rect 5276 5234 5304 6015
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5262 4176 5318 4185
rect 5262 4111 5318 4120
rect 5276 4078 5304 4111
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5172 3528 5224 3534
rect 5092 3476 5172 3482
rect 5092 3470 5224 3476
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5092 3454 5212 3470
rect 5092 2514 5120 3454
rect 5276 3194 5304 3470
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5368 2854 5396 8463
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5460 7546 5488 7890
rect 5552 7818 5580 9046
rect 5630 8800 5686 8809
rect 5630 8735 5686 8744
rect 5644 8498 5672 8735
rect 5736 8634 5764 9386
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5828 8514 5856 10526
rect 5906 10503 5962 10512
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5920 9926 5948 10066
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5920 9489 5948 9862
rect 5906 9480 5962 9489
rect 5906 9415 5962 9424
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5736 8486 5856 8514
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5538 7032 5594 7041
rect 5538 6967 5594 6976
rect 5552 6866 5580 6967
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5460 5914 5488 6258
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5552 5166 5580 6598
rect 5644 6254 5672 6598
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5538 4856 5594 4865
rect 5538 4791 5594 4800
rect 5552 4185 5580 4791
rect 5538 4176 5594 4185
rect 5538 4111 5594 4120
rect 5538 3632 5594 3641
rect 5538 3567 5540 3576
rect 5592 3567 5594 3576
rect 5540 3538 5592 3544
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5644 2650 5672 6054
rect 5736 5098 5764 8486
rect 5920 7886 5948 9318
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5814 7304 5870 7313
rect 5814 7239 5870 7248
rect 5828 7002 5856 7239
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 5724 4684 5776 4690
rect 5828 4672 5856 6734
rect 5776 4644 5856 4672
rect 5724 4626 5776 4632
rect 5736 3058 5764 4626
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 5722 2816 5778 2825
rect 5722 2751 5778 2760
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 5092 2106 5120 2450
rect 5080 2100 5132 2106
rect 5080 2042 5132 2048
rect 5356 1828 5408 1834
rect 5356 1770 5408 1776
rect 5368 480 5396 1770
rect 5736 480 5764 2751
rect 5828 2514 5856 2926
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5920 2310 5948 7822
rect 6012 2802 6040 13495
rect 6104 12889 6132 14311
rect 6090 12880 6146 12889
rect 6090 12815 6146 12824
rect 6104 11626 6132 12815
rect 6196 12238 6224 15642
rect 6288 14074 6316 15864
rect 6380 14618 6408 18006
rect 6472 17202 6500 18022
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6472 16130 6500 17138
rect 6564 16697 6592 20182
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6656 19378 6684 19790
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6656 18766 6684 19314
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6656 17202 6684 18702
rect 6840 17882 6868 19450
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6550 16688 6606 16697
rect 6550 16623 6606 16632
rect 6472 16102 6592 16130
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6472 15065 6500 15982
rect 6458 15056 6514 15065
rect 6458 14991 6514 15000
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6380 12866 6408 13738
rect 6472 12986 6500 14991
rect 6564 14550 6592 16102
rect 6656 16046 6684 17138
rect 6840 16794 6868 17682
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6932 16454 6960 17818
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6656 15473 6684 15982
rect 6932 15978 6960 16390
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6642 15464 6698 15473
rect 6642 15399 6698 15408
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6656 14278 6684 15399
rect 6748 15337 6776 15846
rect 6734 15328 6790 15337
rect 6734 15263 6790 15272
rect 6644 14272 6696 14278
rect 6564 14232 6644 14260
rect 6564 13326 6592 14232
rect 6644 14214 6696 14220
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6656 12918 6684 14010
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6748 13841 6776 13874
rect 6734 13832 6790 13841
rect 6734 13767 6790 13776
rect 6840 13530 6868 15846
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6932 15162 6960 15302
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 6748 13190 6776 13398
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6644 12912 6696 12918
rect 6380 12838 6500 12866
rect 6748 12889 6776 13126
rect 6644 12854 6696 12860
rect 6734 12880 6790 12889
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6276 12708 6328 12714
rect 6276 12650 6328 12656
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6288 11898 6316 12650
rect 6380 12442 6408 12718
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6472 12186 6500 12838
rect 6734 12815 6790 12824
rect 6840 12714 6868 13262
rect 6932 13002 6960 14758
rect 7024 13190 7052 22320
rect 7392 19009 7420 22320
rect 7760 20482 7788 22320
rect 7484 20454 7788 20482
rect 7378 19000 7434 19009
rect 7378 18935 7434 18944
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7194 18456 7250 18465
rect 7194 18391 7250 18400
rect 7208 18057 7236 18391
rect 7194 18048 7250 18057
rect 7194 17983 7250 17992
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7116 17678 7144 17818
rect 7196 17740 7248 17746
rect 7196 17682 7248 17688
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 16794 7144 17478
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7208 15706 7236 17682
rect 7300 16776 7328 18566
rect 7392 17882 7420 18770
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7484 17218 7512 20454
rect 8128 20346 8156 22320
rect 8300 21276 8352 21282
rect 8300 21218 8352 21224
rect 7564 20324 7616 20330
rect 8128 20318 8248 20346
rect 7564 20266 7616 20272
rect 7576 20058 7604 20266
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7562 19000 7618 19009
rect 7562 18935 7618 18944
rect 7576 17320 7604 18935
rect 7668 18426 7696 19994
rect 8024 19984 8076 19990
rect 8024 19926 8076 19932
rect 8036 19378 8064 19926
rect 8220 19394 8248 20318
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 8128 19366 8248 19394
rect 8128 19242 8156 19366
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 7760 18630 7788 19178
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7760 18290 7788 18566
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8312 17898 8340 21218
rect 8496 20346 8524 22320
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 8496 20318 8616 20346
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8404 19514 8432 19858
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 8390 19408 8446 19417
rect 8390 19343 8446 19352
rect 8404 18578 8432 19343
rect 8496 18698 8524 20198
rect 8588 19145 8616 20318
rect 8668 20256 8720 20262
rect 8668 20198 8720 20204
rect 8574 19136 8630 19145
rect 8574 19071 8630 19080
rect 8484 18692 8536 18698
rect 8484 18634 8536 18640
rect 8404 18550 8524 18578
rect 8390 18456 8446 18465
rect 8390 18391 8446 18400
rect 8404 18057 8432 18391
rect 8390 18048 8446 18057
rect 8390 17983 8446 17992
rect 8312 17870 8432 17898
rect 8404 17746 8432 17870
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 7852 17338 7880 17478
rect 8312 17338 8340 17614
rect 7840 17332 7892 17338
rect 7576 17292 7788 17320
rect 7484 17190 7604 17218
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7300 16748 7420 16776
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7300 15706 7328 16594
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7286 15600 7342 15609
rect 7286 15535 7342 15544
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7116 14346 7144 15438
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7208 14074 7236 14962
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7116 13569 7144 13670
rect 7102 13560 7158 13569
rect 7102 13495 7158 13504
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 6932 12974 7052 13002
rect 6828 12708 6880 12714
rect 6748 12668 6828 12696
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6380 12158 6500 12186
rect 6552 12164 6604 12170
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6380 11626 6408 12158
rect 6552 12106 6604 12112
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6368 11620 6420 11626
rect 6368 11562 6420 11568
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6104 7342 6132 10406
rect 6182 10296 6238 10305
rect 6182 10231 6238 10240
rect 6196 10062 6224 10231
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6196 8537 6224 9998
rect 6182 8528 6238 8537
rect 6182 8463 6238 8472
rect 6182 8392 6238 8401
rect 6182 8327 6238 8336
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6196 7154 6224 8327
rect 6288 8072 6316 11290
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6380 10266 6408 10610
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6368 9648 6420 9654
rect 6366 9616 6368 9625
rect 6420 9616 6422 9625
rect 6366 9551 6422 9560
rect 6366 9480 6422 9489
rect 6366 9415 6422 9424
rect 6380 8265 6408 9415
rect 6366 8256 6422 8265
rect 6366 8191 6422 8200
rect 6288 8044 6408 8072
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6288 7546 6316 7890
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6104 7126 6224 7154
rect 6104 5574 6132 7126
rect 6182 7032 6238 7041
rect 6380 7018 6408 8044
rect 6472 7585 6500 12038
rect 6564 11830 6592 12106
rect 6552 11824 6604 11830
rect 6552 11766 6604 11772
rect 6656 11098 6684 12378
rect 6748 12322 6776 12668
rect 6828 12650 6880 12656
rect 7024 12322 7052 12974
rect 7116 12481 7144 13330
rect 7102 12472 7158 12481
rect 7102 12407 7158 12416
rect 6748 12294 6960 12322
rect 7024 12294 7236 12322
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6748 11286 6776 11630
rect 6840 11286 6868 12174
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 6932 11218 6960 12294
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7012 11620 7064 11626
rect 7012 11562 7064 11568
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7024 11150 7052 11562
rect 7116 11354 7144 12038
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 6564 11070 6684 11098
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 6564 10062 6592 11070
rect 6642 10976 6698 10985
rect 6642 10911 6698 10920
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6564 8090 6592 9862
rect 6656 8809 6684 10911
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6748 10690 6776 10746
rect 6826 10704 6882 10713
rect 6748 10662 6826 10690
rect 6826 10639 6882 10648
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6642 8800 6698 8809
rect 6642 8735 6698 8744
rect 6748 8537 6776 10474
rect 6840 9654 6868 10542
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6932 10169 6960 10406
rect 6918 10160 6974 10169
rect 6918 10095 6974 10104
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6826 9480 6882 9489
rect 6826 9415 6882 9424
rect 6840 9081 6868 9415
rect 6826 9072 6882 9081
rect 6826 9007 6828 9016
rect 6880 9007 6882 9016
rect 6828 8978 6880 8984
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6734 8528 6790 8537
rect 6656 8486 6734 8514
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6458 7576 6514 7585
rect 6458 7511 6514 7520
rect 6182 6967 6238 6976
rect 6288 6990 6408 7018
rect 6196 6118 6224 6967
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6196 5409 6224 6054
rect 6182 5400 6238 5409
rect 6182 5335 6238 5344
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6196 3194 6224 4966
rect 6288 4457 6316 6990
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6380 6662 6408 6802
rect 6472 6780 6500 7511
rect 6564 7313 6592 7686
rect 6656 7478 6684 8486
rect 6840 8498 6868 8842
rect 6734 8463 6790 8472
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6826 8256 6882 8265
rect 6826 8191 6882 8200
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6550 7304 6606 7313
rect 6550 7239 6606 7248
rect 6734 7032 6790 7041
rect 6734 6967 6790 6976
rect 6748 6798 6776 6967
rect 6552 6792 6604 6798
rect 6472 6752 6552 6780
rect 6736 6792 6788 6798
rect 6552 6734 6604 6740
rect 6656 6752 6736 6780
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6458 6624 6514 6633
rect 6458 6559 6514 6568
rect 6366 6488 6422 6497
rect 6366 6423 6422 6432
rect 6380 6322 6408 6423
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6472 6254 6500 6559
rect 6656 6458 6684 6752
rect 6736 6734 6788 6740
rect 6840 6610 6868 8191
rect 6932 7410 6960 9998
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6748 6582 6868 6610
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6748 5930 6776 6582
rect 6472 5902 6776 5930
rect 6274 4448 6330 4457
rect 6274 4383 6330 4392
rect 6288 4078 6316 4383
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6380 3466 6408 3878
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6092 2916 6144 2922
rect 6288 2904 6316 3334
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6144 2876 6316 2904
rect 6092 2858 6144 2864
rect 6012 2774 6224 2802
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 6196 480 6224 2774
rect 6380 2446 6408 2994
rect 6472 2825 6500 5902
rect 6932 5817 6960 6598
rect 6918 5808 6974 5817
rect 6552 5772 6604 5778
rect 6918 5743 6974 5752
rect 6552 5714 6604 5720
rect 6458 2816 6514 2825
rect 6458 2751 6514 2760
rect 6564 2650 6592 5714
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6748 5273 6776 5578
rect 6840 5302 6868 5646
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6828 5296 6880 5302
rect 6734 5264 6790 5273
rect 6828 5238 6880 5244
rect 6734 5199 6790 5208
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6656 4554 6684 4762
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6642 4040 6698 4049
rect 6642 3975 6698 3984
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6656 1034 6684 3975
rect 6748 2990 6776 5102
rect 6840 4826 6868 5238
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6840 3369 6868 4150
rect 6932 4146 6960 5510
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6826 3360 6882 3369
rect 6826 3295 6882 3304
rect 6932 3210 6960 3538
rect 6840 3182 6960 3210
rect 6840 3097 6868 3182
rect 6826 3088 6882 3097
rect 6826 3023 6882 3032
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6840 1630 6868 3023
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6932 2650 6960 2790
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 6828 1624 6880 1630
rect 6828 1566 6880 1572
rect 7024 1034 7052 11086
rect 7116 8362 7144 11290
rect 7208 10713 7236 12294
rect 7300 12073 7328 15535
rect 7392 14414 7420 16748
rect 7484 16590 7512 17002
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7484 16250 7512 16526
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7484 15502 7512 16186
rect 7576 15745 7604 17190
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7668 16590 7696 17070
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7562 15736 7618 15745
rect 7668 15706 7696 15846
rect 7562 15671 7618 15680
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7470 15192 7526 15201
rect 7470 15127 7526 15136
rect 7484 14822 7512 15127
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7576 14634 7604 15506
rect 7654 15464 7710 15473
rect 7654 15399 7710 15408
rect 7668 14822 7696 15399
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7484 14606 7604 14634
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7484 14278 7512 14606
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7392 13462 7420 14214
rect 7470 13968 7526 13977
rect 7470 13903 7472 13912
rect 7524 13903 7526 13912
rect 7472 13874 7524 13880
rect 7472 13796 7524 13802
rect 7472 13738 7524 13744
rect 7380 13456 7432 13462
rect 7380 13398 7432 13404
rect 7380 13320 7432 13326
rect 7378 13288 7380 13297
rect 7432 13288 7434 13297
rect 7378 13223 7434 13232
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7286 12064 7342 12073
rect 7286 11999 7342 12008
rect 7392 10810 7420 12582
rect 7484 12209 7512 13738
rect 7576 12442 7604 14418
rect 7668 13938 7696 14758
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7760 13512 7788 17292
rect 7840 17274 7892 17280
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8022 17232 8078 17241
rect 8022 17167 8024 17176
rect 8076 17167 8078 17176
rect 8024 17138 8076 17144
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8312 16726 8340 17274
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 8392 15972 8444 15978
rect 8392 15914 8444 15920
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8220 15502 8248 15914
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8114 15056 8170 15065
rect 8114 14991 8116 15000
rect 8168 14991 8170 15000
rect 8298 15056 8354 15065
rect 8298 14991 8354 15000
rect 8116 14962 8168 14968
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8024 14544 8076 14550
rect 8024 14486 8076 14492
rect 8036 13852 8064 14486
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8128 14074 8156 14350
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8116 13864 8168 13870
rect 8036 13824 8116 13852
rect 8116 13806 8168 13812
rect 8312 13802 8340 14991
rect 8300 13796 8352 13802
rect 8300 13738 8352 13744
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7668 13484 7788 13512
rect 8208 13524 8260 13530
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7668 12306 7696 13484
rect 8208 13466 8260 13472
rect 7840 13456 7892 13462
rect 7840 13398 7892 13404
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7656 12300 7708 12306
rect 7576 12260 7656 12288
rect 7470 12200 7526 12209
rect 7470 12135 7526 12144
rect 7576 12073 7604 12260
rect 7656 12242 7708 12248
rect 7562 12064 7618 12073
rect 7562 11999 7618 12008
rect 7760 11914 7788 13126
rect 7852 12782 7880 13398
rect 8220 13297 8248 13466
rect 8300 13320 8352 13326
rect 8206 13288 8262 13297
rect 8300 13262 8352 13268
rect 8206 13223 8262 13232
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 8114 12336 8170 12345
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7668 11886 7788 11914
rect 7852 11898 7880 12174
rect 7944 11898 7972 12310
rect 8114 12271 8170 12280
rect 8128 12170 8156 12271
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 7840 11892 7892 11898
rect 7470 11656 7526 11665
rect 7470 11591 7526 11600
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7194 10704 7250 10713
rect 7194 10639 7250 10648
rect 7288 10532 7340 10538
rect 7288 10474 7340 10480
rect 7300 9994 7328 10474
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 7208 9081 7236 9590
rect 7194 9072 7250 9081
rect 7194 9007 7250 9016
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 7116 6186 7144 7414
rect 7208 7018 7236 9007
rect 7300 7154 7328 9930
rect 7392 9926 7420 10066
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7392 8809 7420 9862
rect 7378 8800 7434 8809
rect 7378 8735 7434 8744
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7392 8294 7420 8366
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7484 7449 7512 11591
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 10538 7604 10610
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7668 9654 7696 11886
rect 7840 11834 7892 11840
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 7760 11218 7788 11766
rect 8220 11694 8248 13126
rect 8312 12986 8340 13262
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8298 12336 8354 12345
rect 8298 12271 8354 12280
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 8128 10742 8156 11222
rect 8116 10736 8168 10742
rect 8116 10678 8168 10684
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8220 10470 8248 10542
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7760 10266 7788 10406
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 8114 10160 8170 10169
rect 8114 10095 8116 10104
rect 8168 10095 8170 10104
rect 8116 10066 8168 10072
rect 7748 9920 7800 9926
rect 8220 9897 8248 10406
rect 7748 9862 7800 9868
rect 8206 9888 8262 9897
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7576 9110 7604 9522
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7470 7440 7526 7449
rect 7470 7375 7526 7384
rect 7300 7126 7420 7154
rect 7208 6990 7328 7018
rect 7300 6934 7328 6990
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 7102 6080 7158 6089
rect 7102 6015 7158 6024
rect 7116 5273 7144 6015
rect 7208 5914 7236 6870
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7300 6633 7328 6666
rect 7286 6624 7342 6633
rect 7286 6559 7342 6568
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7300 5953 7328 6054
rect 7286 5944 7342 5953
rect 7196 5908 7248 5914
rect 7286 5879 7342 5888
rect 7196 5850 7248 5856
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7102 5264 7158 5273
rect 7102 5199 7158 5208
rect 7116 4282 7144 5199
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7208 4078 7236 5306
rect 7300 4826 7328 5714
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7286 4584 7342 4593
rect 7286 4519 7342 4528
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 7116 1698 7144 3470
rect 7208 2922 7236 3470
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7208 2417 7236 2586
rect 7194 2408 7250 2417
rect 7194 2343 7250 2352
rect 7208 1970 7236 2343
rect 7196 1964 7248 1970
rect 7196 1906 7248 1912
rect 7104 1692 7156 1698
rect 7104 1634 7156 1640
rect 6564 1006 6684 1034
rect 6932 1006 7052 1034
rect 6564 480 6592 1006
rect 6932 480 6960 1006
rect 7300 480 7328 4519
rect 7392 1834 7420 7126
rect 7576 7041 7604 8230
rect 7668 7886 7696 8978
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7656 7744 7708 7750
rect 7654 7712 7656 7721
rect 7708 7712 7710 7721
rect 7654 7647 7710 7656
rect 7760 7206 7788 9862
rect 8206 9823 8262 9832
rect 7932 9444 7984 9450
rect 8312 9432 8340 12271
rect 8404 11286 8432 15914
rect 8496 15609 8524 18550
rect 8680 18329 8708 20198
rect 8772 19961 8800 20538
rect 8758 19952 8814 19961
rect 8956 19938 8984 22320
rect 9324 20262 9352 22320
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 8956 19910 9352 19938
rect 8758 19887 8814 19896
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 8944 19780 8996 19786
rect 8944 19722 8996 19728
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8772 18834 8800 19450
rect 8852 18896 8904 18902
rect 8852 18838 8904 18844
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8666 18320 8722 18329
rect 8666 18255 8722 18264
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8588 17882 8616 18090
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8772 17746 8800 18770
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8588 16454 8616 17002
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 8482 15600 8538 15609
rect 8588 15570 8616 16390
rect 8482 15535 8538 15544
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8484 15428 8536 15434
rect 8484 15370 8536 15376
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 8496 11098 8524 15370
rect 8680 14498 8708 17682
rect 8864 17134 8892 18838
rect 8956 18290 8984 19722
rect 9048 18426 9076 19790
rect 9220 19236 9272 19242
rect 9220 19178 9272 19184
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 9034 18048 9090 18057
rect 9034 17983 9090 17992
rect 9048 17762 9076 17983
rect 9140 17882 9168 18702
rect 9232 18630 9260 19178
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9232 18290 9260 18566
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 9048 17734 9168 17762
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8942 16688 8998 16697
rect 8942 16623 8998 16632
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8760 16040 8812 16046
rect 8864 16017 8892 16390
rect 8760 15982 8812 15988
rect 8850 16008 8906 16017
rect 8772 15638 8800 15982
rect 8850 15943 8906 15952
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8864 15706 8892 15846
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8588 14470 8708 14498
rect 8588 13190 8616 14470
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8680 12918 8708 13262
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8588 12073 8616 12242
rect 8680 12170 8708 12854
rect 8772 12481 8800 14554
rect 8758 12472 8814 12481
rect 8758 12407 8814 12416
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8574 12064 8630 12073
rect 8574 11999 8630 12008
rect 8574 11928 8630 11937
rect 8574 11863 8630 11872
rect 8404 11070 8524 11098
rect 8404 10690 8432 11070
rect 8588 10962 8616 11863
rect 8680 11830 8708 12106
rect 8668 11824 8720 11830
rect 8668 11766 8720 11772
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8668 11620 8720 11626
rect 8668 11562 8720 11568
rect 8680 11121 8708 11562
rect 8772 11354 8800 11698
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8666 11112 8722 11121
rect 8666 11047 8722 11056
rect 8496 10934 8616 10962
rect 8496 10849 8524 10934
rect 8482 10840 8538 10849
rect 8482 10775 8538 10784
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8404 10662 8524 10690
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8404 10062 8432 10474
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 7984 9404 8340 9432
rect 7932 9386 7984 9392
rect 8312 9353 8340 9404
rect 8298 9344 8354 9353
rect 7820 9276 8116 9296
rect 8298 9279 8354 9288
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8206 9208 8262 9217
rect 8206 9143 8208 9152
rect 8260 9143 8262 9152
rect 8208 9114 8260 9120
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 8022 8800 8078 8809
rect 8022 8735 8078 8744
rect 8036 8430 8064 8735
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8128 8276 8156 9046
rect 8298 8936 8354 8945
rect 8404 8906 8432 9998
rect 8298 8871 8354 8880
rect 8392 8900 8444 8906
rect 8312 8430 8340 8871
rect 8392 8842 8444 8848
rect 8300 8424 8352 8430
rect 8496 8378 8524 10662
rect 8588 10130 8616 10746
rect 8760 10532 8812 10538
rect 8760 10474 8812 10480
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8300 8366 8352 8372
rect 8404 8350 8524 8378
rect 8128 8248 8248 8276
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8220 8072 8248 8248
rect 8036 8044 8248 8072
rect 8036 7954 8064 8044
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 7932 7336 7984 7342
rect 8036 7324 8064 7890
rect 8220 7478 8248 7890
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 7984 7296 8064 7324
rect 8300 7336 8352 7342
rect 7932 7278 7984 7284
rect 8300 7278 8352 7284
rect 8208 7268 8260 7274
rect 8208 7210 8260 7216
rect 7748 7200 7800 7206
rect 7654 7168 7710 7177
rect 7748 7142 7800 7148
rect 7654 7103 7710 7112
rect 7562 7032 7618 7041
rect 7562 6967 7618 6976
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7484 5914 7512 6734
rect 7576 6712 7604 6967
rect 7668 6916 7696 7103
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7748 6928 7800 6934
rect 7668 6888 7748 6916
rect 7748 6870 7800 6876
rect 8022 6896 8078 6905
rect 8022 6831 8078 6840
rect 7840 6724 7892 6730
rect 7576 6684 7840 6712
rect 7840 6666 7892 6672
rect 8036 6633 8064 6831
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8022 6624 8078 6633
rect 8022 6559 8078 6568
rect 8128 6474 8156 6734
rect 7576 6446 8156 6474
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7470 5672 7526 5681
rect 7470 5607 7472 5616
rect 7524 5607 7526 5616
rect 7472 5578 7524 5584
rect 7576 5522 7604 6446
rect 8220 6168 8248 7210
rect 8312 6662 8340 7278
rect 8404 6746 8432 8350
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8496 7993 8524 8230
rect 8482 7984 8538 7993
rect 8482 7919 8538 7928
rect 8588 7546 8616 9862
rect 8680 9761 8708 10202
rect 8666 9752 8722 9761
rect 8772 9722 8800 10474
rect 8864 10266 8892 15506
rect 8956 14006 8984 16623
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8956 13025 8984 13942
rect 8942 13016 8998 13025
rect 8942 12951 8998 12960
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8956 11694 8984 12582
rect 8944 11688 8996 11694
rect 9048 11665 9076 17614
rect 9140 15065 9168 17734
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 9324 15586 9352 19910
rect 9496 19916 9548 19922
rect 9496 19858 9548 19864
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9416 18902 9444 19246
rect 9404 18896 9456 18902
rect 9404 18838 9456 18844
rect 9508 18426 9536 19858
rect 9692 19802 9720 22320
rect 10060 22250 10088 22320
rect 10060 22222 10180 22250
rect 9864 19984 9916 19990
rect 9864 19926 9916 19932
rect 9692 19774 9812 19802
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9692 19310 9720 19654
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9600 18426 9628 18566
rect 9692 18426 9720 18770
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9784 18306 9812 19774
rect 9508 18278 9812 18306
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9416 17338 9444 17682
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9508 15688 9536 18278
rect 9588 18216 9640 18222
rect 9772 18216 9824 18222
rect 9588 18158 9640 18164
rect 9770 18184 9772 18193
rect 9824 18184 9826 18193
rect 9600 17202 9628 18158
rect 9680 18148 9732 18154
rect 9770 18119 9826 18128
rect 9680 18090 9732 18096
rect 9692 17882 9720 18090
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9784 17338 9812 18022
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9600 16794 9628 17138
rect 9680 16992 9732 16998
rect 9732 16952 9812 16980
rect 9680 16934 9732 16940
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9600 16114 9628 16730
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9508 15660 9628 15688
rect 9126 15056 9182 15065
rect 9126 14991 9182 15000
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 9140 14278 9168 14826
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9140 14074 9168 14214
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9140 13394 9168 13738
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 8944 11630 8996 11636
rect 9034 11656 9090 11665
rect 9034 11591 9090 11600
rect 9048 11354 9076 11591
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9034 10976 9090 10985
rect 9034 10911 9090 10920
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8956 10606 8984 10746
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 9048 10130 9076 10911
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9034 10024 9090 10033
rect 9034 9959 9090 9968
rect 8666 9687 8722 9696
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8772 9178 8800 9386
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8680 8129 8708 8298
rect 8666 8120 8722 8129
rect 8666 8055 8722 8064
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8588 6866 8616 7482
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8404 6718 8616 6746
rect 8300 6656 8352 6662
rect 8352 6616 8524 6644
rect 8300 6598 8352 6604
rect 8496 6390 8524 6616
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8211 6140 8248 6168
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 8211 6066 8239 6140
rect 8312 6089 8340 6190
rect 8298 6080 8354 6089
rect 7760 5896 7788 6054
rect 8211 6038 8248 6066
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 7484 5494 7604 5522
rect 7668 5868 7788 5896
rect 7380 1828 7432 1834
rect 7380 1770 7432 1776
rect 7484 1748 7512 5494
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7576 5001 7604 5034
rect 7562 4992 7618 5001
rect 7562 4927 7618 4936
rect 7668 4826 7696 5868
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7576 3913 7604 4218
rect 7562 3904 7618 3913
rect 7562 3839 7618 3848
rect 7760 3670 7788 5578
rect 8220 5370 8248 6038
rect 8298 6015 8354 6024
rect 8404 5710 8432 6258
rect 8588 5846 8616 6718
rect 8666 6624 8722 6633
rect 8666 6559 8722 6568
rect 8680 6458 8708 6559
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 8220 4434 8248 5306
rect 8128 4406 8248 4434
rect 8022 4312 8078 4321
rect 8022 4247 8078 4256
rect 8036 4078 8064 4247
rect 8128 4146 8156 4406
rect 8208 4276 8260 4282
rect 8312 4264 8340 5578
rect 8404 4622 8432 5646
rect 8588 5166 8616 5782
rect 8680 5166 8708 6258
rect 8772 5953 8800 8910
rect 8864 7750 8892 9386
rect 8956 9042 8984 9522
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8956 7818 8984 8978
rect 9048 8265 9076 9959
rect 9034 8256 9090 8265
rect 9034 8191 9090 8200
rect 9140 8072 9168 13330
rect 9232 12345 9260 15574
rect 9324 15558 9444 15586
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9324 14414 9352 15438
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9324 12782 9352 13126
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9218 12336 9274 12345
rect 9218 12271 9274 12280
rect 9220 12096 9272 12102
rect 9416 12050 9444 15558
rect 9600 15201 9628 15660
rect 9586 15192 9642 15201
rect 9586 15127 9642 15136
rect 9588 14884 9640 14890
rect 9588 14826 9640 14832
rect 9600 14618 9628 14826
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9600 13462 9628 14418
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9600 12345 9628 13398
rect 9586 12336 9642 12345
rect 9586 12271 9642 12280
rect 9692 12170 9720 15846
rect 9784 14550 9812 16952
rect 9876 16538 9904 19926
rect 10152 19378 10180 22222
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9968 16658 9996 19178
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10060 19009 10088 19110
rect 10046 19000 10102 19009
rect 10244 18970 10272 19790
rect 10336 19514 10364 19790
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10046 18935 10102 18944
rect 10232 18964 10284 18970
rect 10060 18902 10088 18935
rect 10232 18906 10284 18912
rect 10048 18896 10100 18902
rect 10336 18850 10364 19314
rect 10048 18838 10100 18844
rect 10244 18822 10364 18850
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10060 18578 10088 18702
rect 10060 18550 10180 18578
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 10060 18086 10088 18362
rect 10152 18154 10180 18550
rect 10140 18148 10192 18154
rect 10140 18090 10192 18096
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10060 17882 10088 18022
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 10060 16538 10088 16934
rect 9876 16510 10088 16538
rect 9862 15600 9918 15609
rect 9862 15535 9918 15544
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9220 12038 9272 12044
rect 9232 11830 9260 12038
rect 9324 12022 9444 12050
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9324 11676 9352 12022
rect 9402 11928 9458 11937
rect 9600 11898 9628 12038
rect 9402 11863 9458 11872
rect 9588 11892 9640 11898
rect 9416 11812 9444 11863
rect 9588 11834 9640 11840
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9416 11784 9536 11812
rect 9508 11694 9536 11784
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9232 11648 9352 11676
rect 9496 11688 9548 11694
rect 9232 10418 9260 11648
rect 9600 11665 9628 11698
rect 9496 11630 9548 11636
rect 9586 11656 9642 11665
rect 9586 11591 9642 11600
rect 9404 11552 9456 11558
rect 9588 11552 9640 11558
rect 9456 11512 9588 11540
rect 9404 11494 9456 11500
rect 9588 11494 9640 11500
rect 9692 11354 9720 11834
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9784 11234 9812 14350
rect 9876 14074 9904 15535
rect 10060 14482 10088 16510
rect 10152 16250 10180 17614
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9862 13832 9918 13841
rect 9862 13767 9918 13776
rect 9876 12730 9904 13767
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9968 13258 9996 13466
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9876 12702 9996 12730
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9876 12306 9904 12582
rect 9968 12306 9996 12702
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9692 11206 9812 11234
rect 9312 10736 9364 10742
rect 9310 10704 9312 10713
rect 9364 10704 9366 10713
rect 9310 10639 9366 10648
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9232 10390 9352 10418
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9232 10169 9260 10202
rect 9218 10160 9274 10169
rect 9218 10095 9274 10104
rect 9324 9926 9352 10390
rect 9508 10266 9536 10542
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9416 9874 9444 10066
rect 9508 10010 9536 10202
rect 9600 10130 9628 10542
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9508 9982 9628 10010
rect 9692 9994 9720 11206
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9218 9616 9274 9625
rect 9218 9551 9274 9560
rect 9232 9178 9260 9551
rect 9324 9382 9352 9862
rect 9416 9846 9536 9874
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9218 8936 9274 8945
rect 9218 8871 9274 8880
rect 9048 8044 9168 8072
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8758 5944 8814 5953
rect 8758 5879 8814 5888
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8482 4856 8538 4865
rect 8588 4826 8616 4966
rect 8482 4791 8538 4800
rect 8576 4820 8628 4826
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8260 4236 8340 4264
rect 8208 4218 8260 4224
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7576 1902 7604 3538
rect 8128 3505 8156 3606
rect 8114 3496 8170 3505
rect 8114 3431 8170 3440
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 7668 2582 7696 3334
rect 7746 3224 7802 3233
rect 7746 3159 7802 3168
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7760 1902 7788 3159
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8116 2576 8168 2582
rect 8022 2544 8078 2553
rect 8116 2518 8168 2524
rect 8022 2479 8078 2488
rect 7564 1896 7616 1902
rect 7564 1838 7616 1844
rect 7748 1896 7800 1902
rect 7748 1838 7800 1844
rect 7484 1720 7696 1748
rect 7668 480 7696 1720
rect 8036 480 8064 2479
rect 8128 1766 8156 2518
rect 8220 2514 8248 3334
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8312 2378 8340 3674
rect 8404 3534 8432 4558
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8404 3194 8432 3470
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8496 3097 8524 4791
rect 8576 4762 8628 4768
rect 8576 4140 8628 4146
rect 8680 4128 8708 5102
rect 8628 4100 8708 4128
rect 8576 4082 8628 4088
rect 8482 3088 8538 3097
rect 8482 3023 8538 3032
rect 8588 2990 8616 4082
rect 8666 3904 8722 3913
rect 8666 3839 8722 3848
rect 8680 3602 8708 3839
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8576 2984 8628 2990
rect 8482 2952 8538 2961
rect 8772 2972 8800 5879
rect 8864 3398 8892 7142
rect 8956 6798 8984 7210
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 9048 5930 9076 8044
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9140 6497 9168 7890
rect 9232 7886 9260 8871
rect 9324 8634 9352 8978
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9312 8492 9364 8498
rect 9416 8480 9444 9658
rect 9508 9518 9536 9846
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9508 9178 9536 9318
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9494 9072 9550 9081
rect 9494 9007 9550 9016
rect 9364 8452 9444 8480
rect 9312 8434 9364 8440
rect 9508 8378 9536 9007
rect 9416 8350 9536 8378
rect 9416 7936 9444 8350
rect 9600 8276 9628 9982
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9784 9722 9812 10066
rect 9876 9897 9904 12106
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9968 11558 9996 11698
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9954 11384 10010 11393
rect 9954 11319 10010 11328
rect 9968 11218 9996 11319
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9954 10568 10010 10577
rect 9954 10503 10010 10512
rect 9862 9888 9918 9897
rect 9862 9823 9918 9832
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9324 7908 9444 7936
rect 9508 8248 9628 8276
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9232 7478 9260 7686
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 9324 7177 9352 7908
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9416 7410 9444 7754
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9508 7274 9536 8248
rect 9692 7750 9720 9590
rect 9862 9480 9918 9489
rect 9862 9415 9918 9424
rect 9876 9081 9904 9415
rect 9968 9382 9996 10503
rect 10060 9489 10088 14282
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10152 12889 10180 13738
rect 10244 13394 10272 18822
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10336 16250 10364 18158
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10428 15745 10456 22320
rect 10600 18828 10652 18834
rect 10652 18788 10732 18816
rect 10600 18770 10652 18776
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10612 18222 10640 18634
rect 10600 18216 10652 18222
rect 10704 18193 10732 18788
rect 10600 18158 10652 18164
rect 10690 18184 10746 18193
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10520 16182 10548 16934
rect 10612 16658 10640 18158
rect 10690 18119 10746 18128
rect 10796 17270 10824 22320
rect 11164 18850 11192 22320
rect 11624 20670 11652 22320
rect 11612 20664 11664 20670
rect 11612 20606 11664 20612
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11072 18822 11192 18850
rect 11520 18828 11572 18834
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 10784 17264 10836 17270
rect 10784 17206 10836 17212
rect 10980 17202 11008 17682
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10966 16960 11022 16969
rect 10966 16895 11022 16904
rect 10980 16726 11008 16895
rect 11072 16794 11100 18822
rect 11572 18788 11744 18816
rect 11520 18770 11572 18776
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11164 17134 11192 18702
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 11256 17746 11284 18090
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11624 17202 11652 17478
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10508 16176 10560 16182
rect 10508 16118 10560 16124
rect 10612 16046 10640 16594
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10414 15736 10470 15745
rect 10414 15671 10470 15680
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10428 14074 10456 15506
rect 10508 15496 10560 15502
rect 10692 15496 10744 15502
rect 10508 15438 10560 15444
rect 10598 15464 10654 15473
rect 10520 14618 10548 15438
rect 10692 15438 10744 15444
rect 10598 15399 10654 15408
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10612 14362 10640 15399
rect 10704 14890 10732 15438
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10692 14544 10744 14550
rect 10692 14486 10744 14492
rect 10520 14334 10640 14362
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10520 13530 10548 14334
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10612 13938 10640 14214
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10704 13530 10732 14486
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10796 13938 10824 14350
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10796 13462 10824 13874
rect 10784 13456 10836 13462
rect 10598 13424 10654 13433
rect 10232 13388 10284 13394
rect 10784 13398 10836 13404
rect 10598 13359 10654 13368
rect 10692 13388 10744 13394
rect 10232 13330 10284 13336
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10230 13016 10286 13025
rect 10230 12951 10286 12960
rect 10138 12880 10194 12889
rect 10244 12850 10272 12951
rect 10520 12850 10548 13262
rect 10138 12815 10194 12824
rect 10232 12844 10284 12850
rect 10152 12730 10180 12815
rect 10232 12786 10284 12792
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10152 12702 10364 12730
rect 10232 12640 10284 12646
rect 10138 12608 10194 12617
rect 10232 12582 10284 12588
rect 10138 12543 10194 12552
rect 10046 9480 10102 9489
rect 10046 9415 10102 9424
rect 9956 9376 10008 9382
rect 10152 9364 10180 12543
rect 10244 12442 10272 12582
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10244 11354 10272 12038
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10336 10554 10364 12702
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10428 12209 10456 12582
rect 10612 12481 10640 13359
rect 10692 13330 10744 13336
rect 10598 12472 10654 12481
rect 10598 12407 10654 12416
rect 10414 12200 10470 12209
rect 10414 12135 10470 12144
rect 10704 11744 10732 13330
rect 10796 12850 10824 13398
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10888 12424 10916 15846
rect 11256 15570 11284 15982
rect 11348 15638 11376 15982
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10980 12782 11008 14554
rect 11334 14512 11390 14521
rect 11152 14476 11204 14482
rect 11334 14447 11336 14456
rect 11152 14418 11204 14424
rect 11388 14447 11390 14456
rect 11336 14418 11388 14424
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 11072 13734 11100 14350
rect 11164 14074 11192 14418
rect 11428 14408 11480 14414
rect 11426 14376 11428 14385
rect 11520 14408 11572 14414
rect 11480 14376 11482 14385
rect 11520 14350 11572 14356
rect 11426 14311 11482 14320
rect 11532 14260 11560 14350
rect 11532 14232 11652 14260
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11152 14068 11204 14074
rect 11624 14056 11652 14232
rect 11152 14010 11204 14016
rect 11532 14028 11652 14056
rect 11150 13968 11206 13977
rect 11532 13938 11560 14028
rect 11150 13903 11206 13912
rect 11520 13932 11572 13938
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11164 13530 11192 13903
rect 11520 13874 11572 13880
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11520 13728 11572 13734
rect 11518 13696 11520 13705
rect 11572 13696 11574 13705
rect 11518 13631 11574 13640
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11058 13152 11114 13161
rect 11058 13087 11114 13096
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10888 12396 11008 12424
rect 10876 12300 10928 12306
rect 10612 11716 10732 11744
rect 10796 12260 10876 12288
rect 10414 11656 10470 11665
rect 10414 11591 10470 11600
rect 10428 11286 10456 11591
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10244 10526 10364 10554
rect 10244 9704 10272 10526
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 10033 10364 10406
rect 10322 10024 10378 10033
rect 10322 9959 10378 9968
rect 10416 9716 10468 9722
rect 10244 9676 10364 9704
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 9956 9318 10008 9324
rect 10060 9336 10180 9364
rect 9862 9072 9918 9081
rect 9968 9042 9996 9318
rect 9862 9007 9918 9016
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9496 7268 9548 7274
rect 9496 7210 9548 7216
rect 9600 7206 9628 7482
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9588 7200 9640 7206
rect 9310 7168 9366 7177
rect 9588 7142 9640 7148
rect 9310 7103 9366 7112
rect 9218 7032 9274 7041
rect 9218 6967 9220 6976
rect 9272 6967 9274 6976
rect 9220 6938 9272 6944
rect 9312 6792 9364 6798
rect 9364 6752 9444 6780
rect 9312 6734 9364 6740
rect 9126 6488 9182 6497
rect 9126 6423 9182 6432
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9140 6118 9168 6326
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9048 5902 9168 5930
rect 9140 5828 9168 5902
rect 8942 5808 8998 5817
rect 8942 5743 8944 5752
rect 8996 5743 8998 5752
rect 9048 5800 9168 5828
rect 8944 5714 8996 5720
rect 8956 3641 8984 5714
rect 8942 3632 8998 3641
rect 8942 3567 8998 3576
rect 8942 3496 8998 3505
rect 8942 3431 8998 3440
rect 8956 3398 8984 3431
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8576 2926 8628 2932
rect 8680 2944 8800 2972
rect 8482 2887 8538 2896
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8404 2514 8432 2790
rect 8496 2582 8524 2887
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8404 2038 8432 2450
rect 8680 2446 8708 2944
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8392 2032 8444 2038
rect 8392 1974 8444 1980
rect 8116 1760 8168 1766
rect 8680 1714 8708 2382
rect 8772 2281 8800 2790
rect 8864 2514 8892 3130
rect 9048 3097 9076 5800
rect 9232 5098 9260 6190
rect 9324 5710 9352 6326
rect 9416 6322 9444 6752
rect 9692 6458 9720 7210
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9680 6248 9732 6254
rect 9784 6225 9812 8910
rect 10060 8809 10088 9336
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10046 8800 10102 8809
rect 10046 8735 10102 8744
rect 10060 8480 10088 8735
rect 9968 8452 10088 8480
rect 9862 8120 9918 8129
rect 9862 8055 9918 8064
rect 9876 7290 9904 8055
rect 9968 7698 9996 8452
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 10060 7818 10088 8298
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 9968 7670 10088 7698
rect 9876 7262 9996 7290
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 7002 9904 7142
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9862 6488 9918 6497
rect 9862 6423 9918 6432
rect 9680 6190 9732 6196
rect 9770 6216 9826 6225
rect 9402 5808 9458 5817
rect 9692 5778 9720 6190
rect 9770 6151 9826 6160
rect 9784 5778 9812 6151
rect 9402 5743 9458 5752
rect 9680 5772 9732 5778
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 9232 4865 9260 5034
rect 9218 4856 9274 4865
rect 9218 4791 9274 4800
rect 9126 4312 9182 4321
rect 9126 4247 9182 4256
rect 9140 3738 9168 4247
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9310 3904 9366 3913
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9232 3670 9260 3878
rect 9310 3839 9366 3848
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9034 3088 9090 3097
rect 9034 3023 9090 3032
rect 9324 2854 9352 3839
rect 9416 3602 9444 5743
rect 9680 5714 9732 5720
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9680 5636 9732 5642
rect 9732 5596 9812 5624
rect 9680 5578 9732 5584
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9508 4865 9536 5306
rect 9600 5166 9628 5510
rect 9784 5370 9812 5596
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9494 4856 9550 4865
rect 9494 4791 9550 4800
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 9126 2680 9182 2689
rect 9126 2615 9182 2624
rect 8942 2544 8998 2553
rect 8852 2508 8904 2514
rect 9140 2514 9168 2615
rect 9312 2576 9364 2582
rect 9312 2518 9364 2524
rect 8942 2479 8998 2488
rect 9128 2508 9180 2514
rect 8852 2450 8904 2456
rect 8758 2272 8814 2281
rect 8758 2207 8814 2216
rect 8116 1702 8168 1708
rect 8404 1686 8708 1714
rect 8404 480 8432 1686
rect 8772 480 8800 2207
rect 8956 2145 8984 2479
rect 9128 2450 9180 2456
rect 9128 2304 9180 2310
rect 9324 2292 9352 2518
rect 9180 2264 9352 2292
rect 9128 2246 9180 2252
rect 8942 2136 8998 2145
rect 8942 2071 8998 2080
rect 9140 480 9168 2246
rect 9508 480 9536 4490
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9600 2922 9628 4082
rect 9692 3738 9720 4626
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9784 2802 9812 5306
rect 9876 5030 9904 6423
rect 9968 5234 9996 7262
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9876 2922 9904 4422
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 9784 2774 9904 2802
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 1426 9720 2246
rect 9680 1420 9732 1426
rect 9680 1362 9732 1368
rect 9876 480 9904 2774
rect 9968 2514 9996 4966
rect 10060 4593 10088 7670
rect 10152 5370 10180 9114
rect 10244 9058 10272 9522
rect 10336 9178 10364 9676
rect 10416 9658 10468 9664
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10244 9030 10364 9058
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10244 8498 10272 8910
rect 10336 8820 10364 9030
rect 10428 8945 10456 9658
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10414 8936 10470 8945
rect 10414 8871 10470 8880
rect 10336 8792 10456 8820
rect 10322 8664 10378 8673
rect 10322 8599 10378 8608
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10244 8022 10272 8298
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10336 7857 10364 8599
rect 10428 8498 10456 8792
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10414 8392 10470 8401
rect 10414 8327 10416 8336
rect 10468 8327 10470 8336
rect 10416 8298 10468 8304
rect 10520 8129 10548 9114
rect 10612 8294 10640 11716
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10704 11354 10732 11562
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10704 9382 10732 11290
rect 10796 10742 10824 12260
rect 10876 12242 10928 12248
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 10888 11626 10916 12106
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 10874 11384 10930 11393
rect 10874 11319 10930 11328
rect 10784 10736 10836 10742
rect 10784 10678 10836 10684
rect 10796 10248 10824 10678
rect 10888 10606 10916 11319
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10796 10220 10916 10248
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10796 9761 10824 10066
rect 10888 10062 10916 10220
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10782 9752 10838 9761
rect 10782 9687 10838 9696
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10704 9178 10732 9318
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10796 8974 10824 9114
rect 10784 8968 10836 8974
rect 10704 8916 10784 8922
rect 10704 8910 10836 8916
rect 10704 8894 10824 8910
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10506 8120 10562 8129
rect 10506 8055 10562 8064
rect 10416 7880 10468 7886
rect 10322 7848 10378 7857
rect 10232 7812 10284 7818
rect 10612 7857 10640 8230
rect 10704 7954 10732 8894
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10416 7822 10468 7828
rect 10598 7848 10654 7857
rect 10322 7783 10378 7792
rect 10232 7754 10284 7760
rect 10244 7478 10272 7754
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 10428 7274 10456 7822
rect 10598 7783 10654 7792
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10416 7268 10468 7274
rect 10416 7210 10468 7216
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10244 6662 10272 7142
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10336 5574 10364 6734
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10138 5128 10194 5137
rect 10322 5128 10378 5137
rect 10138 5063 10194 5072
rect 10232 5092 10284 5098
rect 10046 4584 10102 4593
rect 10046 4519 10102 4528
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10060 4282 10088 4422
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10152 4162 10180 5063
rect 10284 5072 10322 5080
rect 10284 5063 10378 5072
rect 10284 5052 10364 5063
rect 10232 5034 10284 5040
rect 10322 4584 10378 4593
rect 10322 4519 10378 4528
rect 10060 4134 10180 4162
rect 10060 2854 10088 4134
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10244 3534 10272 3878
rect 10336 3738 10364 4519
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10140 3528 10192 3534
rect 10138 3496 10140 3505
rect 10232 3528 10284 3534
rect 10192 3496 10194 3505
rect 10232 3470 10284 3476
rect 10138 3431 10194 3440
rect 10138 3088 10194 3097
rect 10244 3058 10272 3470
rect 10428 3398 10456 6598
rect 10520 5846 10548 7346
rect 10508 5840 10560 5846
rect 10508 5782 10560 5788
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10520 4826 10548 5034
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10520 4078 10548 4626
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10612 4010 10640 7686
rect 10690 7576 10746 7585
rect 10690 7511 10746 7520
rect 10704 7041 10732 7511
rect 10690 7032 10746 7041
rect 10690 6967 10746 6976
rect 10690 6624 10746 6633
rect 10690 6559 10746 6568
rect 10704 6089 10732 6559
rect 10690 6080 10746 6089
rect 10690 6015 10746 6024
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 10704 5545 10732 5578
rect 10690 5536 10746 5545
rect 10690 5471 10746 5480
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10704 4826 10732 5102
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10704 4321 10732 4762
rect 10690 4312 10746 4321
rect 10690 4247 10746 4256
rect 10796 4162 10824 8774
rect 10888 7750 10916 9590
rect 10980 9450 11008 12396
rect 11072 10606 11100 13087
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11428 12912 11480 12918
rect 11428 12854 11480 12860
rect 11518 12880 11574 12889
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11060 10600 11112 10606
rect 11164 10577 11192 12718
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11348 12238 11376 12582
rect 11440 12238 11468 12854
rect 11518 12815 11574 12824
rect 11532 12345 11560 12815
rect 11624 12424 11652 13806
rect 11716 13530 11744 18788
rect 11808 18154 11836 19110
rect 11796 18148 11848 18154
rect 11796 18090 11848 18096
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11900 17678 11928 17750
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11796 17128 11848 17134
rect 11794 17096 11796 17105
rect 11848 17096 11850 17105
rect 11794 17031 11850 17040
rect 11900 16658 11928 17614
rect 11992 16794 12020 22320
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12268 19990 12296 20402
rect 12164 19984 12216 19990
rect 12164 19926 12216 19932
rect 12256 19984 12308 19990
rect 12256 19926 12308 19932
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 12084 19378 12112 19790
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 12084 18834 12112 19314
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12084 18426 12112 18770
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 12084 16833 12112 17682
rect 12070 16824 12126 16833
rect 11980 16788 12032 16794
rect 12070 16759 12126 16768
rect 11980 16730 12032 16736
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 16182 11836 16390
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11796 15972 11848 15978
rect 11796 15914 11848 15920
rect 11808 15162 11836 15914
rect 11900 15910 11928 16594
rect 11992 16153 12020 16594
rect 11978 16144 12034 16153
rect 11978 16079 12034 16088
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11808 13394 11836 15098
rect 11900 15026 11928 15846
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11992 14822 12020 15506
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11900 14414 11928 14758
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11624 12396 11744 12424
rect 11518 12336 11574 12345
rect 11518 12271 11574 12280
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11532 12084 11560 12271
rect 11532 12056 11652 12084
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11532 11082 11560 11222
rect 11520 11076 11572 11082
rect 11520 11018 11572 11024
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11060 10542 11112 10548
rect 11150 10568 11206 10577
rect 11256 10538 11284 10610
rect 11150 10503 11206 10512
rect 11244 10532 11296 10538
rect 11244 10474 11296 10480
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10980 8634 11008 8774
rect 11072 8673 11100 10406
rect 11152 9920 11204 9926
rect 11256 9908 11284 10474
rect 11348 10266 11376 10678
rect 11624 10606 11652 12056
rect 11716 11354 11744 12396
rect 11808 11762 11836 13194
rect 11900 12617 11928 13942
rect 11992 13530 12020 14214
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 11978 13152 12034 13161
rect 11978 13087 12034 13096
rect 11886 12608 11942 12617
rect 11886 12543 11942 12552
rect 11900 12442 11928 12543
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11900 11626 11928 11766
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11808 10810 11836 11018
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11518 10432 11574 10441
rect 11518 10367 11574 10376
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11532 9994 11560 10367
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11204 9880 11284 9908
rect 11152 9862 11204 9868
rect 11058 8664 11114 8673
rect 10968 8628 11020 8634
rect 11058 8599 11114 8608
rect 11164 8616 11192 9862
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11334 9480 11390 9489
rect 11334 9415 11390 9424
rect 11520 9444 11572 9450
rect 11348 8945 11376 9415
rect 11520 9386 11572 9392
rect 11532 9194 11560 9386
rect 11624 9330 11652 10542
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11716 10266 11744 10474
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11716 9897 11744 10066
rect 11702 9888 11758 9897
rect 11702 9823 11758 9832
rect 11794 9752 11850 9761
rect 11794 9687 11850 9696
rect 11702 9480 11758 9489
rect 11808 9450 11836 9687
rect 11900 9586 11928 11562
rect 11992 11558 12020 13087
rect 12084 12782 12112 16662
rect 12176 16250 12204 19926
rect 12254 19136 12310 19145
rect 12254 19071 12310 19080
rect 12268 18834 12296 19071
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12268 17270 12296 17614
rect 12360 17338 12388 22320
rect 12728 20058 12756 22320
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12452 19514 12480 19858
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12544 18170 12572 19246
rect 12636 18426 12664 19858
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12728 18426 12756 19110
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12452 18142 12572 18170
rect 12716 18216 12768 18222
rect 12820 18204 12848 19654
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12768 18176 12848 18204
rect 12716 18158 12768 18164
rect 12452 17338 12480 18142
rect 12532 18080 12584 18086
rect 12530 18048 12532 18057
rect 12584 18048 12586 18057
rect 12530 17983 12586 17992
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12544 17134 12572 17682
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12714 17096 12770 17105
rect 12912 17066 12940 18702
rect 13004 18290 13032 18838
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13096 17882 13124 22320
rect 13464 19786 13492 22320
rect 13832 20058 13860 22320
rect 14004 20256 14056 20262
rect 14004 20198 14056 20204
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13266 19000 13322 19009
rect 13266 18935 13322 18944
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12714 17031 12716 17040
rect 12768 17031 12770 17040
rect 12900 17060 12952 17066
rect 12716 17002 12768 17008
rect 12900 17002 12952 17008
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 12176 13530 12204 15302
rect 12728 14929 12756 15846
rect 12820 15162 12848 16934
rect 12912 16590 12940 17002
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 12912 15502 12940 16526
rect 13004 16454 13032 17138
rect 13096 16969 13124 17682
rect 13188 17542 13216 18090
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13082 16960 13138 16969
rect 13082 16895 13138 16904
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 13004 16114 13032 16390
rect 13280 16114 13308 18935
rect 13464 18601 13492 19110
rect 13450 18592 13506 18601
rect 13450 18527 13506 18536
rect 13556 17785 13584 19110
rect 13648 18290 13676 19314
rect 13832 18630 13860 19654
rect 13924 19009 13952 19858
rect 13910 19000 13966 19009
rect 13910 18935 13966 18944
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13912 18352 13964 18358
rect 13726 18320 13782 18329
rect 13636 18284 13688 18290
rect 13912 18294 13964 18300
rect 13726 18255 13782 18264
rect 13636 18226 13688 18232
rect 13542 17776 13598 17785
rect 13542 17711 13598 17720
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13358 16824 13414 16833
rect 13358 16759 13414 16768
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12714 14920 12770 14929
rect 12440 14884 12492 14890
rect 12714 14855 12770 14864
rect 12440 14826 12492 14832
rect 12452 14249 12480 14826
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12438 14240 12494 14249
rect 12438 14175 12494 14184
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 12162 12472 12218 12481
rect 12162 12407 12164 12416
rect 12216 12407 12218 12416
rect 12164 12378 12216 12384
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12176 11665 12204 11834
rect 12162 11656 12218 11665
rect 12162 11591 12218 11600
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12162 11520 12218 11529
rect 12084 11354 12112 11494
rect 12162 11455 12218 11464
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11992 10810 12020 11086
rect 12084 11082 12112 11290
rect 12176 11218 12204 11455
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12162 10840 12218 10849
rect 11980 10804 12032 10810
rect 12162 10775 12218 10784
rect 11980 10746 12032 10752
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11702 9415 11704 9424
rect 11756 9415 11758 9424
rect 11796 9444 11848 9450
rect 11704 9386 11756 9392
rect 11796 9386 11848 9392
rect 11992 9382 12020 10542
rect 12070 10296 12126 10305
rect 12070 10231 12126 10240
rect 12084 10033 12112 10231
rect 12070 10024 12126 10033
rect 12070 9959 12126 9968
rect 12072 9920 12124 9926
rect 12176 9908 12204 10775
rect 12360 10606 12388 13126
rect 12440 12776 12492 12782
rect 12544 12764 12572 14758
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12492 12736 12572 12764
rect 12440 12718 12492 12724
rect 12452 11694 12480 12718
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12452 11150 12480 11630
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12544 10742 12572 12174
rect 12636 11014 12664 13398
rect 12728 12442 12756 14350
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12820 11608 12848 14758
rect 12898 14376 12954 14385
rect 12898 14311 12954 14320
rect 12728 11580 12848 11608
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12728 10826 12756 11580
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12636 10798 12756 10826
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12636 10305 12664 10798
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12438 10296 12494 10305
rect 12438 10231 12440 10240
rect 12492 10231 12494 10240
rect 12622 10296 12678 10305
rect 12622 10231 12678 10240
rect 12440 10202 12492 10208
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12124 9880 12204 9908
rect 12072 9862 12124 9868
rect 11980 9376 12032 9382
rect 11624 9302 11744 9330
rect 11980 9318 12032 9324
rect 11532 9166 11652 9194
rect 11334 8936 11390 8945
rect 11334 8871 11390 8880
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11164 8588 11284 8616
rect 10968 8570 11020 8576
rect 11256 8129 11284 8588
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11242 8120 11298 8129
rect 11242 8055 11298 8064
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11072 7868 11100 7958
rect 11348 7868 11376 8434
rect 11440 8401 11468 8502
rect 11426 8392 11482 8401
rect 11426 8327 11482 8336
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11072 7840 11376 7868
rect 11440 7800 11468 7958
rect 11164 7772 11468 7800
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 11058 7712 11114 7721
rect 11058 7647 11114 7656
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10980 7342 11008 7414
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10888 7002 10916 7142
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10980 6662 11008 7142
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 10888 5409 10916 6326
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10980 5846 11008 6054
rect 10968 5840 11020 5846
rect 10968 5782 11020 5788
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10874 5400 10930 5409
rect 10874 5335 10930 5344
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10888 4690 10916 5170
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10980 4214 11008 5646
rect 10968 4208 11020 4214
rect 10796 4134 10916 4162
rect 10968 4150 11020 4156
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10796 3534 10824 4014
rect 10888 3738 10916 4134
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10506 3360 10562 3369
rect 10506 3295 10562 3304
rect 10138 3023 10194 3032
rect 10232 3052 10284 3058
rect 10152 2990 10180 3023
rect 10232 2994 10284 3000
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10232 2848 10284 2854
rect 10520 2836 10548 3295
rect 10796 2990 10824 3470
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10980 3097 11008 3130
rect 10966 3088 11022 3097
rect 10966 3023 11022 3032
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10520 2808 10640 2836
rect 10232 2790 10284 2796
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 9968 2106 9996 2450
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 10244 480 10272 2790
rect 10612 480 10640 2808
rect 11072 2650 11100 7647
rect 11164 7528 11192 7772
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11164 7500 11376 7528
rect 11150 7168 11206 7177
rect 11150 7103 11206 7112
rect 11164 6934 11192 7103
rect 11242 7032 11298 7041
rect 11242 6967 11244 6976
rect 11296 6967 11298 6976
rect 11244 6938 11296 6944
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 11348 6780 11376 7500
rect 11624 7410 11652 9166
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11440 6798 11468 7142
rect 11532 7002 11560 7278
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11624 7002 11652 7210
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11164 6752 11376 6780
rect 11428 6792 11480 6798
rect 11164 5710 11192 6752
rect 11428 6734 11480 6740
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11624 6186 11652 6734
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11716 6066 11744 9302
rect 12084 9194 12112 9862
rect 11992 9166 12112 9194
rect 11992 8480 12020 9166
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 12084 8650 12112 9046
rect 12084 8622 12204 8650
rect 11900 8452 12020 8480
rect 11900 8344 11928 8452
rect 12176 8412 12204 8622
rect 11624 6038 11744 6066
rect 11808 8316 11928 8344
rect 12084 8384 12204 8412
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11164 5234 11192 5510
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11440 4826 11468 4966
rect 11518 4856 11574 4865
rect 11428 4820 11480 4826
rect 11518 4791 11574 4800
rect 11428 4762 11480 4768
rect 11532 4690 11560 4791
rect 11624 4758 11652 6038
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11716 5545 11744 5714
rect 11702 5536 11758 5545
rect 11702 5471 11758 5480
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11612 4752 11664 4758
rect 11612 4694 11664 4700
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11716 4622 11744 5238
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11612 4480 11664 4486
rect 11808 4434 11836 8316
rect 11886 7848 11942 7857
rect 11886 7783 11942 7792
rect 11900 6866 11928 7783
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11992 6798 12020 7686
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11886 6624 11942 6633
rect 11886 6559 11942 6568
rect 11900 5846 11928 6559
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11612 4422 11664 4428
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11624 4146 11652 4422
rect 11716 4406 11836 4434
rect 11900 4604 11928 5102
rect 11992 5098 12020 6394
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 12084 4842 12112 8384
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 7324 12204 8230
rect 12268 8022 12296 10066
rect 12360 9722 12388 10066
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12360 9178 12388 9454
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12452 9110 12480 9862
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12544 8974 12572 9454
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12360 8498 12388 8774
rect 12530 8664 12586 8673
rect 12530 8599 12586 8608
rect 12438 8528 12494 8537
rect 12348 8492 12400 8498
rect 12438 8463 12494 8472
rect 12348 8434 12400 8440
rect 12452 8430 12480 8463
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12544 8362 12572 8599
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 8090 12480 8230
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12256 8016 12308 8022
rect 12544 7970 12572 8298
rect 12256 7958 12308 7964
rect 12360 7942 12572 7970
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12268 7478 12296 7686
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12176 7296 12296 7324
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12176 6458 12204 6870
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12268 6338 12296 7296
rect 12176 6310 12296 6338
rect 12176 4978 12204 6310
rect 12360 6254 12388 7942
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12452 7342 12480 7686
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12452 6254 12480 7278
rect 12544 7177 12572 7278
rect 12530 7168 12586 7177
rect 12530 7103 12586 7112
rect 12636 6730 12664 10134
rect 12728 8922 12756 10406
rect 12820 9450 12848 10950
rect 12912 9761 12940 14311
rect 13004 13394 13032 15642
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 13569 13124 14758
rect 13188 14346 13216 15030
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13176 14340 13228 14346
rect 13176 14282 13228 14288
rect 13082 13560 13138 13569
rect 13082 13495 13138 13504
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13004 13025 13032 13330
rect 12990 13016 13046 13025
rect 12990 12951 13046 12960
rect 13096 11937 13124 13495
rect 13280 13258 13308 14894
rect 13372 14618 13400 16759
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13188 12102 13216 12650
rect 13280 12646 13308 13194
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13372 12442 13400 14418
rect 13464 13530 13492 17206
rect 13648 17202 13676 18226
rect 13740 17338 13768 18255
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13728 17060 13780 17066
rect 13728 17002 13780 17008
rect 13542 16280 13598 16289
rect 13542 16215 13598 16224
rect 13556 16182 13584 16215
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13556 14414 13584 15506
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13544 13864 13596 13870
rect 13648 13852 13676 14758
rect 13596 13824 13676 13852
rect 13544 13806 13596 13812
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13556 13394 13584 13806
rect 13740 13462 13768 17002
rect 13832 16250 13860 18158
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13924 15586 13952 18294
rect 13832 15558 13952 15586
rect 13832 13734 13860 15558
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13924 14958 13952 15438
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13176 12096 13228 12102
rect 13280 12084 13308 12378
rect 13358 12336 13414 12345
rect 13358 12271 13414 12280
rect 13372 12238 13400 12271
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13280 12056 13492 12084
rect 13176 12038 13228 12044
rect 13082 11928 13138 11937
rect 13082 11863 13138 11872
rect 13358 11928 13414 11937
rect 13358 11863 13414 11872
rect 13266 11248 13322 11257
rect 13266 11183 13322 11192
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 13004 9994 13032 10746
rect 13176 10736 13228 10742
rect 13096 10696 13176 10724
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 12898 9752 12954 9761
rect 12898 9687 12954 9696
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 13004 9382 13032 9930
rect 13096 9722 13124 10696
rect 13176 10678 13228 10684
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12728 8894 12848 8922
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12530 6488 12586 6497
rect 12530 6423 12586 6432
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12544 6118 12572 6423
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12636 5930 12664 6190
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12544 5902 12664 5930
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12268 5302 12296 5646
rect 12360 5574 12388 5850
rect 12452 5778 12480 5850
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12544 5642 12572 5902
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12532 5636 12584 5642
rect 12584 5596 12664 5624
rect 12532 5578 12584 5584
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12452 5409 12480 5578
rect 12438 5400 12494 5409
rect 12438 5335 12494 5344
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12256 5160 12308 5166
rect 12254 5128 12256 5137
rect 12308 5128 12310 5137
rect 12254 5063 12310 5072
rect 12440 5024 12492 5030
rect 12176 4950 12388 4978
rect 12440 4966 12492 4972
rect 12084 4814 12296 4842
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12072 4616 12124 4622
rect 11900 4576 12072 4604
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11336 3732 11388 3738
rect 11440 3720 11468 3946
rect 11520 3732 11572 3738
rect 11440 3692 11520 3720
rect 11336 3674 11388 3680
rect 11520 3674 11572 3680
rect 11348 3618 11376 3674
rect 11348 3590 11652 3618
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11256 2922 11468 2938
rect 11244 2916 11468 2922
rect 11296 2910 11468 2916
rect 11244 2858 11296 2864
rect 11440 2854 11468 2910
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11150 2544 11206 2553
rect 10968 2508 11020 2514
rect 11150 2479 11206 2488
rect 11334 2544 11390 2553
rect 11334 2479 11336 2488
rect 10968 2450 11020 2456
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10796 2106 10824 2246
rect 10784 2100 10836 2106
rect 10784 2042 10836 2048
rect 10980 480 11008 2450
rect 11164 1442 11192 2479
rect 11388 2479 11390 2488
rect 11336 2450 11388 2456
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11164 1414 11376 1442
rect 11348 480 11376 1414
rect 11624 762 11652 3590
rect 11716 2446 11744 4406
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 2514 11836 3878
rect 11900 3602 11928 4576
rect 12072 4558 12124 4564
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 11978 4040 12034 4049
rect 11978 3975 12034 3984
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11992 3058 12020 3975
rect 12084 3126 12112 4082
rect 12176 3534 12204 4626
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12176 3398 12204 3470
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12176 2990 12204 3334
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11992 1442 12020 2790
rect 12268 2582 12296 4814
rect 12360 3482 12388 4950
rect 12452 4826 12480 4966
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12530 4312 12586 4321
rect 12530 4247 12586 4256
rect 12544 4078 12572 4247
rect 12636 4146 12664 5596
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12440 4004 12492 4010
rect 12440 3946 12492 3952
rect 12452 3738 12480 3946
rect 12532 3936 12584 3942
rect 12530 3904 12532 3913
rect 12584 3904 12586 3913
rect 12530 3839 12586 3848
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12360 3454 12572 3482
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12360 2961 12388 3130
rect 12346 2952 12402 2961
rect 12346 2887 12402 2896
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 11992 1414 12204 1442
rect 11624 734 11836 762
rect 11808 480 11836 734
rect 12176 480 12204 1414
rect 12544 480 12572 3454
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12636 3194 12664 3402
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12728 2310 12756 8774
rect 12820 8566 12848 8894
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12820 7002 12848 8366
rect 12912 7750 12940 9114
rect 13004 9042 13032 9318
rect 13188 9110 13216 10406
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 13084 8968 13136 8974
rect 13136 8928 13216 8956
rect 13084 8910 13136 8916
rect 12990 8800 13046 8809
rect 12990 8735 13046 8744
rect 13004 8634 13032 8735
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13004 7886 13032 8434
rect 13096 8362 13124 8502
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 13082 8120 13138 8129
rect 13082 8055 13138 8064
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13096 7818 13124 8055
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12898 7576 12954 7585
rect 12898 7511 12954 7520
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12820 6497 12848 6938
rect 12806 6488 12862 6497
rect 12806 6423 12862 6432
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12820 5574 12848 6054
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 12820 1290 12848 5170
rect 12912 5114 12940 7511
rect 13188 7018 13216 8928
rect 13280 8294 13308 11183
rect 13372 8809 13400 11863
rect 13464 11778 13492 12056
rect 13556 11898 13584 13194
rect 13924 12782 13952 14214
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 14016 12424 14044 20198
rect 14096 19168 14148 19174
rect 14096 19110 14148 19116
rect 14108 18902 14136 19110
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 17678 14136 18566
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14108 17134 14136 17614
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14200 17066 14228 22320
rect 14660 20244 14688 22320
rect 15028 20262 15056 22320
rect 15292 20664 15344 20670
rect 15292 20606 15344 20612
rect 15108 20324 15160 20330
rect 15108 20266 15160 20272
rect 14384 20216 14688 20244
rect 15016 20256 15068 20262
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14292 18970 14320 19178
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14384 18193 14412 20216
rect 15016 20198 15068 20204
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 15120 19922 15148 20266
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 14370 18184 14426 18193
rect 14370 18119 14426 18128
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14278 17912 14334 17921
rect 14278 17847 14334 17856
rect 14188 17060 14240 17066
rect 14188 17002 14240 17008
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 14108 16114 14136 16390
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 14108 15638 14136 16050
rect 14186 16008 14242 16017
rect 14186 15943 14242 15952
rect 14096 15632 14148 15638
rect 14096 15574 14148 15580
rect 14108 14414 14136 15574
rect 14096 14408 14148 14414
rect 14094 14376 14096 14385
rect 14148 14376 14150 14385
rect 14094 14311 14150 14320
rect 14200 14074 14228 15943
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 14108 12918 14136 13738
rect 14200 13394 14228 14010
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 13832 12396 14044 12424
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 11937 13768 12174
rect 13726 11928 13782 11937
rect 13544 11892 13596 11898
rect 13596 11852 13676 11880
rect 13726 11863 13782 11872
rect 13544 11834 13596 11840
rect 13464 11750 13584 11778
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13464 9178 13492 10678
rect 13556 10266 13584 11750
rect 13648 10418 13676 11852
rect 13726 11248 13782 11257
rect 13726 11183 13728 11192
rect 13780 11183 13782 11192
rect 13728 11154 13780 11160
rect 13726 11112 13782 11121
rect 13726 11047 13782 11056
rect 13740 10674 13768 11047
rect 13832 10713 13860 12396
rect 14094 12336 14150 12345
rect 14004 12300 14056 12306
rect 14094 12271 14150 12280
rect 14004 12242 14056 12248
rect 14016 11801 14044 12242
rect 14002 11792 14058 11801
rect 14002 11727 14058 11736
rect 14108 11393 14136 12271
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14094 11384 14150 11393
rect 14094 11319 14150 11328
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 13818 10704 13874 10713
rect 13728 10668 13780 10674
rect 13924 10674 13952 11018
rect 13818 10639 13874 10648
rect 13912 10668 13964 10674
rect 13728 10610 13780 10616
rect 13912 10610 13964 10616
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13648 10390 13860 10418
rect 13634 10296 13690 10305
rect 13544 10260 13596 10266
rect 13634 10231 13690 10240
rect 13544 10202 13596 10208
rect 13542 9752 13598 9761
rect 13542 9687 13598 9696
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13556 9058 13584 9687
rect 13648 9081 13676 10231
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13464 9030 13584 9058
rect 13634 9072 13690 9081
rect 13358 8800 13414 8809
rect 13358 8735 13414 8744
rect 13464 8378 13492 9030
rect 13634 9007 13690 9016
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13372 8350 13492 8378
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13096 6990 13216 7018
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 13004 5846 13032 6666
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 12912 5098 13032 5114
rect 12912 5092 13044 5098
rect 12912 5086 12992 5092
rect 12992 5034 13044 5040
rect 12900 5024 12952 5030
rect 12898 4992 12900 5001
rect 12952 4992 12954 5001
rect 12898 4927 12954 4936
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12912 3670 12940 4422
rect 13096 3942 13124 6990
rect 13174 6080 13230 6089
rect 13174 6015 13230 6024
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12808 1284 12860 1290
rect 12808 1226 12860 1232
rect 12912 480 12940 3334
rect 13004 1766 13032 3878
rect 13082 3088 13138 3097
rect 13082 3023 13084 3032
rect 13136 3023 13138 3032
rect 13084 2994 13136 3000
rect 13188 2582 13216 6015
rect 13280 4486 13308 8230
rect 13372 8022 13400 8350
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13358 7576 13414 7585
rect 13358 7511 13414 7520
rect 13372 7002 13400 7511
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13372 4729 13400 6734
rect 13358 4720 13414 4729
rect 13358 4655 13414 4664
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13360 4276 13412 4282
rect 13360 4218 13412 4224
rect 13280 3398 13308 4218
rect 13372 4010 13400 4218
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 12992 1760 13044 1766
rect 12992 1702 13044 1708
rect 13280 480 13308 3130
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13372 2582 13400 2994
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 13464 2514 13492 8230
rect 13556 7274 13584 8774
rect 13648 8430 13676 8910
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13544 7268 13596 7274
rect 13544 7210 13596 7216
rect 13648 6712 13676 7890
rect 13740 7342 13768 9862
rect 13832 9654 13860 10390
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13924 9466 13952 10474
rect 13832 9438 13952 9466
rect 13832 8974 13860 9438
rect 13912 9172 13964 9178
rect 14016 9160 14044 11154
rect 14200 11014 14228 11630
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14108 10606 14136 10950
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14200 10441 14228 10542
rect 14186 10432 14242 10441
rect 14186 10367 14242 10376
rect 14292 10248 14320 17847
rect 14384 16969 14412 18022
rect 14370 16960 14426 16969
rect 14370 16895 14426 16904
rect 14370 16688 14426 16697
rect 14370 16623 14372 16632
rect 14424 16623 14426 16632
rect 14372 16594 14424 16600
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14384 15065 14412 16186
rect 14370 15056 14426 15065
rect 14370 14991 14426 15000
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14384 12889 14412 14418
rect 14476 12986 14504 19858
rect 15304 19786 15332 20606
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 14922 19408 14978 19417
rect 14922 19343 14978 19352
rect 15108 19372 15160 19378
rect 14936 19310 14964 19343
rect 15108 19314 15160 19320
rect 14924 19304 14976 19310
rect 14924 19246 14976 19252
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14554 18184 14610 18193
rect 14554 18119 14610 18128
rect 14568 16658 14596 18119
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14660 17649 14688 17682
rect 14646 17640 14702 17649
rect 14646 17575 14702 17584
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 15028 16250 15056 19110
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14556 15564 14608 15570
rect 15016 15564 15068 15570
rect 14608 15524 14688 15552
rect 14556 15506 14608 15512
rect 14660 15366 14688 15524
rect 15016 15506 15068 15512
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14568 14890 14596 15302
rect 14556 14884 14608 14890
rect 14556 14826 14608 14832
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14370 12880 14426 12889
rect 14568 12850 14596 14826
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14648 14544 14700 14550
rect 14648 14486 14700 14492
rect 14660 13802 14688 14486
rect 15028 14362 15056 15506
rect 15120 14550 15148 19314
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15212 16114 15240 17682
rect 15304 17649 15332 18906
rect 15290 17640 15346 17649
rect 15290 17575 15346 17584
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15304 16114 15332 17070
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15304 15706 15332 15846
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15396 15337 15424 22320
rect 15476 19984 15528 19990
rect 15476 19926 15528 19932
rect 15488 18970 15516 19926
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15672 19514 15700 19858
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15488 17762 15516 18226
rect 15488 17734 15608 17762
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15488 16726 15516 17614
rect 15580 16794 15608 17734
rect 15764 17626 15792 22320
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15856 18465 15884 19790
rect 15934 19544 15990 19553
rect 15934 19479 15990 19488
rect 15948 19378 15976 19479
rect 15936 19372 15988 19378
rect 16132 19360 16160 22320
rect 16500 20890 16528 22320
rect 16316 20862 16528 20890
rect 16212 19440 16264 19446
rect 16212 19382 16264 19388
rect 15936 19314 15988 19320
rect 16040 19332 16160 19360
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15842 18456 15898 18465
rect 15948 18426 15976 19110
rect 15842 18391 15898 18400
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15948 17882 15976 18226
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15764 17598 15884 17626
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 16794 15700 17478
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15476 16720 15528 16726
rect 15476 16662 15528 16668
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15672 16250 15700 16594
rect 15750 16552 15806 16561
rect 15750 16487 15806 16496
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15764 15910 15792 16487
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15382 15328 15438 15337
rect 15382 15263 15438 15272
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 15304 14482 15332 14826
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 15028 14334 15148 14362
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14936 13025 14964 13330
rect 14922 13016 14978 13025
rect 14922 12951 14978 12960
rect 14370 12815 14426 12824
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14462 12608 14518 12617
rect 14462 12543 14518 12552
rect 14476 12238 14504 12543
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11898 14780 12038
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14384 11121 14412 11766
rect 14554 11656 14610 11665
rect 14554 11591 14610 11600
rect 14568 11218 14596 11591
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15028 11336 15056 13466
rect 15120 11937 15148 14334
rect 15384 13864 15436 13870
rect 15198 13832 15254 13841
rect 15384 13806 15436 13812
rect 15198 13767 15254 13776
rect 15292 13796 15344 13802
rect 15212 13326 15240 13767
rect 15292 13738 15344 13744
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15304 13172 15332 13738
rect 15396 13190 15424 13806
rect 15212 13144 15332 13172
rect 15384 13184 15436 13190
rect 15212 12646 15240 13144
rect 15384 13126 15436 13132
rect 15290 13016 15346 13025
rect 15290 12951 15346 12960
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15212 12102 15240 12582
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15106 11928 15162 11937
rect 15106 11863 15162 11872
rect 14936 11308 15056 11336
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14370 11112 14426 11121
rect 14370 11047 14426 11056
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14200 10220 14320 10248
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 9518 14136 9862
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 13964 9132 14044 9160
rect 13912 9114 13964 9120
rect 14108 9024 14136 9318
rect 14200 9178 14228 10220
rect 14384 10169 14412 10746
rect 14936 10538 14964 11308
rect 15120 11257 15148 11863
rect 15212 11694 15240 12038
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15106 11248 15162 11257
rect 15106 11183 15162 11192
rect 15014 10976 15070 10985
rect 15014 10911 15070 10920
rect 14924 10532 14976 10538
rect 14924 10474 14976 10480
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14370 10160 14426 10169
rect 14280 10124 14332 10130
rect 14568 10130 14596 10406
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14646 10160 14702 10169
rect 14370 10095 14426 10104
rect 14556 10124 14608 10130
rect 14280 10066 14332 10072
rect 14646 10095 14702 10104
rect 14556 10066 14608 10072
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 13924 8996 14136 9024
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13832 8430 13860 8774
rect 13924 8650 13952 8996
rect 14292 8838 14320 10066
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14384 9738 14412 9862
rect 14384 9710 14504 9738
rect 14476 9654 14504 9710
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14096 8832 14148 8838
rect 14280 8832 14332 8838
rect 14148 8792 14228 8820
rect 14096 8774 14148 8780
rect 13924 8622 14136 8650
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13818 8256 13874 8265
rect 13818 8191 13874 8200
rect 13832 7721 13860 8191
rect 13818 7712 13874 7721
rect 13818 7647 13874 7656
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13820 7200 13872 7206
rect 13726 7168 13782 7177
rect 13924 7188 13952 8502
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 13872 7160 13952 7188
rect 13820 7142 13872 7148
rect 13726 7103 13782 7112
rect 13740 7002 13768 7103
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13648 6684 13768 6712
rect 13740 6322 13768 6684
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13832 6186 13860 7142
rect 14016 6390 14044 8434
rect 14108 8022 14136 8622
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 14094 7576 14150 7585
rect 14094 7511 14150 7520
rect 14108 7041 14136 7511
rect 14200 7478 14228 8792
rect 14280 8774 14332 8780
rect 14278 8664 14334 8673
rect 14278 8599 14334 8608
rect 14188 7472 14240 7478
rect 14188 7414 14240 7420
rect 14094 7032 14150 7041
rect 14292 7018 14320 8599
rect 14384 8498 14412 9454
rect 14568 9432 14596 10066
rect 14476 9404 14596 9432
rect 14476 8922 14504 9404
rect 14660 9364 14688 10095
rect 14924 9580 14976 9586
rect 15028 9568 15056 10911
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 14976 9540 15056 9568
rect 14924 9522 14976 9528
rect 14568 9336 14688 9364
rect 14568 9160 14596 9336
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14568 9132 14688 9160
rect 14660 9042 14688 9132
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14740 8968 14792 8974
rect 14476 8894 14596 8922
rect 14740 8910 14792 8916
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14568 8430 14596 8894
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14660 8276 14688 8774
rect 14752 8566 14780 8910
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14844 8276 14872 8910
rect 15028 8786 15056 9540
rect 15120 8974 15148 9998
rect 15212 9654 15240 9998
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15304 9568 15332 12951
rect 15488 12442 15516 15438
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15580 11762 15608 14758
rect 15672 13569 15700 15506
rect 15764 14385 15792 15846
rect 15750 14376 15806 14385
rect 15750 14311 15806 14320
rect 15750 14240 15806 14249
rect 15750 14175 15806 14184
rect 15658 13560 15714 13569
rect 15764 13530 15792 14175
rect 15658 13495 15714 13504
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15658 13288 15714 13297
rect 15658 13223 15714 13232
rect 15672 12782 15700 13223
rect 15750 13016 15806 13025
rect 15750 12951 15806 12960
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15384 11552 15436 11558
rect 15580 11529 15608 11562
rect 15384 11494 15436 11500
rect 15566 11520 15622 11529
rect 15396 11286 15424 11494
rect 15566 11455 15622 11464
rect 15474 11384 15530 11393
rect 15474 11319 15530 11328
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15396 10130 15424 10610
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15304 9540 15424 9568
rect 15292 9444 15344 9450
rect 15292 9386 15344 9392
rect 15304 9178 15332 9386
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 14568 8248 14872 8276
rect 14936 8758 15056 8786
rect 14936 8276 14964 8758
rect 15014 8664 15070 8673
rect 15014 8599 15070 8608
rect 15028 8430 15056 8599
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 14936 8248 15056 8276
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14384 7410 14412 8026
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14462 7168 14518 7177
rect 14462 7103 14518 7112
rect 14094 6967 14150 6976
rect 14200 6990 14320 7018
rect 14476 7002 14504 7103
rect 14464 6996 14516 7002
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 14016 5846 14044 6326
rect 14200 6186 14228 6990
rect 14464 6938 14516 6944
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14292 6254 14320 6802
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14384 5953 14412 6734
rect 14476 6458 14504 6734
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14370 5944 14426 5953
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14188 5908 14240 5914
rect 14370 5879 14426 5888
rect 14188 5850 14240 5856
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 13726 5672 13782 5681
rect 13726 5607 13782 5616
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13556 3670 13584 5306
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13648 4185 13676 4626
rect 13634 4176 13690 4185
rect 13634 4111 13690 4120
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13542 3496 13598 3505
rect 13542 3431 13598 3440
rect 13556 2990 13584 3431
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 13648 480 13676 3538
rect 13740 3194 13768 5607
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13832 4826 13860 4966
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13832 3074 13860 3946
rect 13910 3904 13966 3913
rect 13910 3839 13966 3848
rect 13924 3738 13952 3839
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13924 3505 13952 3674
rect 14002 3632 14058 3641
rect 14002 3567 14058 3576
rect 13910 3496 13966 3505
rect 13910 3431 13966 3440
rect 14016 3346 14044 3567
rect 13740 3058 13860 3074
rect 13728 3052 13860 3058
rect 13780 3046 13860 3052
rect 13924 3318 14044 3346
rect 13728 2994 13780 3000
rect 13924 2514 13952 3318
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 14016 3058 14044 3130
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14002 2816 14058 2825
rect 14002 2751 14058 2760
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 14016 480 14044 2751
rect 14108 2582 14136 5850
rect 14200 5234 14228 5850
rect 14384 5234 14412 5879
rect 14476 5817 14504 6190
rect 14462 5808 14518 5817
rect 14462 5743 14518 5752
rect 14568 5574 14596 8248
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 15028 8090 15056 8248
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14660 7410 14688 7890
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7478 14780 7686
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 15028 5914 15056 7890
rect 15120 7410 15148 8910
rect 15212 8090 15240 9046
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15106 7168 15162 7177
rect 15106 7103 15162 7112
rect 15120 7002 15148 7103
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 14832 5704 14884 5710
rect 14646 5672 14702 5681
rect 14832 5646 14884 5652
rect 14646 5607 14702 5616
rect 14660 5574 14688 5607
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14844 5370 14872 5646
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14200 4214 14228 5170
rect 15016 5160 15068 5166
rect 14554 5128 14610 5137
rect 14372 5092 14424 5098
rect 15120 5148 15148 6938
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15068 5120 15148 5148
rect 15016 5102 15068 5108
rect 14554 5063 14610 5072
rect 14372 5034 14424 5040
rect 14384 4865 14412 5034
rect 14370 4856 14426 4865
rect 14370 4791 14426 4800
rect 14568 4808 14596 5063
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14568 4780 14688 4808
rect 14660 4690 14688 4780
rect 15014 4720 15070 4729
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14648 4684 14700 4690
rect 15014 4655 15070 4664
rect 14648 4626 14700 4632
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14384 4282 14412 4558
rect 14568 4282 14596 4626
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 14188 4208 14240 4214
rect 14188 4150 14240 4156
rect 14278 3768 14334 3777
rect 14278 3703 14334 3712
rect 14292 3176 14320 3703
rect 14384 3534 14412 4218
rect 14936 4010 14964 4218
rect 15028 4162 15056 4655
rect 15212 4554 15240 6598
rect 15304 5302 15332 8978
rect 15396 6662 15424 9540
rect 15488 7857 15516 11319
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15580 10266 15608 10610
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15580 9110 15608 9454
rect 15672 9178 15700 12378
rect 15764 10266 15792 12951
rect 15856 12730 15884 17598
rect 15936 17536 15988 17542
rect 16040 17513 16068 19332
rect 16120 19236 16172 19242
rect 16120 19178 16172 19184
rect 16132 18426 16160 19178
rect 16224 18970 16252 19382
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 15936 17478 15988 17484
rect 16026 17504 16082 17513
rect 15948 16998 15976 17478
rect 16026 17439 16082 17448
rect 16028 17060 16080 17066
rect 16028 17002 16080 17008
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15948 14940 15976 16934
rect 16040 16590 16068 17002
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 16040 15502 16068 16526
rect 16224 15994 16252 18566
rect 16316 18329 16344 20862
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16486 19544 16542 19553
rect 16592 19514 16620 19926
rect 16486 19479 16542 19488
rect 16580 19508 16632 19514
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16302 18320 16358 18329
rect 16302 18255 16358 18264
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16316 16794 16344 18090
rect 16408 17241 16436 19110
rect 16500 17542 16528 19479
rect 16580 19450 16632 19456
rect 16592 19310 16620 19450
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16672 19236 16724 19242
rect 16672 19178 16724 19184
rect 16684 17882 16712 19178
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16394 17232 16450 17241
rect 16394 17167 16450 17176
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16396 16788 16448 16794
rect 16396 16730 16448 16736
rect 16302 16416 16358 16425
rect 16302 16351 16358 16360
rect 16132 15966 16252 15994
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 16028 14952 16080 14958
rect 15948 14912 16028 14940
rect 16028 14894 16080 14900
rect 16040 14482 16068 14894
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15948 13802 15976 14282
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15948 13190 15976 13262
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15856 12702 15976 12730
rect 15844 12164 15896 12170
rect 15844 12106 15896 12112
rect 15856 11937 15884 12106
rect 15842 11928 15898 11937
rect 15842 11863 15898 11872
rect 15842 11656 15898 11665
rect 15842 11591 15898 11600
rect 15856 11393 15884 11591
rect 15842 11384 15898 11393
rect 15842 11319 15844 11328
rect 15896 11319 15898 11328
rect 15844 11290 15896 11296
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15842 9888 15898 9897
rect 15842 9823 15898 9832
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15764 9518 15792 9590
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15580 8673 15608 8774
rect 15566 8664 15622 8673
rect 15566 8599 15622 8608
rect 15566 8528 15622 8537
rect 15566 8463 15622 8472
rect 15474 7848 15530 7857
rect 15474 7783 15530 7792
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15384 6180 15436 6186
rect 15384 6122 15436 6128
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15396 5234 15424 6122
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 15028 4146 15148 4162
rect 15016 4140 15148 4146
rect 15068 4134 15148 4140
rect 15016 4082 15068 4088
rect 15028 4051 15056 4082
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14476 3602 14504 3878
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14556 3392 14608 3398
rect 14462 3360 14518 3369
rect 14556 3334 14608 3340
rect 14462 3295 14518 3304
rect 14372 3188 14424 3194
rect 14292 3148 14372 3176
rect 14372 3130 14424 3136
rect 14476 3058 14504 3295
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14096 2576 14148 2582
rect 14096 2518 14148 2524
rect 14292 2038 14320 2586
rect 14280 2032 14332 2038
rect 14280 1974 14332 1980
rect 14568 1442 14596 3334
rect 15028 3194 15056 3946
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 15016 3188 15068 3194
rect 15016 3130 15068 3136
rect 14752 3058 14780 3130
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 15120 2990 15148 4134
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15304 2514 15332 5034
rect 15396 4729 15424 5170
rect 15382 4720 15438 4729
rect 15382 4655 15438 4664
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15396 2990 15424 4558
rect 15488 4282 15516 6870
rect 15580 4622 15608 8463
rect 15672 8265 15700 8978
rect 15764 8430 15792 9454
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15658 8256 15714 8265
rect 15658 8191 15714 8200
rect 15672 7993 15700 8191
rect 15658 7984 15714 7993
rect 15658 7919 15714 7928
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15764 7721 15792 7822
rect 15750 7712 15806 7721
rect 15750 7647 15806 7656
rect 15660 7200 15712 7206
rect 15764 7177 15792 7647
rect 15856 7410 15884 9823
rect 15948 9625 15976 12702
rect 16026 12472 16082 12481
rect 16026 12407 16082 12416
rect 16040 11898 16068 12407
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16026 11384 16082 11393
rect 16026 11319 16082 11328
rect 16040 10810 16068 11319
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15934 9616 15990 9625
rect 15934 9551 15990 9560
rect 15934 9208 15990 9217
rect 15934 9143 15990 9152
rect 15948 9042 15976 9143
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15934 8936 15990 8945
rect 15934 8871 15990 8880
rect 15948 8566 15976 8871
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 16026 8392 16082 8401
rect 15948 7750 15976 8366
rect 16026 8327 16082 8336
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 16040 7585 16068 8327
rect 16026 7576 16082 7585
rect 16026 7511 16082 7520
rect 16040 7410 16068 7511
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 15936 7200 15988 7206
rect 15660 7142 15712 7148
rect 15750 7168 15806 7177
rect 15672 7002 15700 7142
rect 15936 7142 15988 7148
rect 15750 7103 15806 7112
rect 15948 7041 15976 7142
rect 15934 7032 15990 7041
rect 15660 6996 15712 7002
rect 15934 6967 15990 6976
rect 15660 6938 15712 6944
rect 16040 6882 16068 7346
rect 15948 6854 16068 6882
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 15488 3942 15516 4218
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 14832 2508 14884 2514
rect 14832 2450 14884 2456
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 14752 2106 14780 2450
rect 14740 2100 14792 2106
rect 14740 2042 14792 2048
rect 14844 1902 14872 2450
rect 15488 1902 15516 3334
rect 15672 2802 15700 6054
rect 15764 4826 15792 6734
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15856 5545 15884 6190
rect 15948 6186 15976 6854
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16040 6390 16068 6734
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 16040 5710 16068 6326
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 15842 5536 15898 5545
rect 15842 5471 15898 5480
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 15856 4865 15884 4966
rect 15842 4856 15898 4865
rect 15752 4820 15804 4826
rect 15842 4791 15898 4800
rect 15752 4762 15804 4768
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15764 3738 15792 3878
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15856 3233 15884 3878
rect 15948 3602 15976 5306
rect 16040 5166 16068 5646
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 16026 4720 16082 4729
rect 16026 4655 16082 4664
rect 16040 4622 16068 4655
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 15842 3224 15898 3233
rect 16132 3194 16160 15966
rect 16212 15904 16264 15910
rect 16210 15872 16212 15881
rect 16264 15872 16266 15881
rect 16210 15807 16266 15816
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 14550 16252 14758
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16224 13841 16252 14350
rect 16210 13832 16266 13841
rect 16210 13767 16266 13776
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 11898 16252 13670
rect 16316 13025 16344 16351
rect 16408 16046 16436 16730
rect 16500 16658 16528 17478
rect 16592 17338 16620 17682
rect 16776 17610 16804 18226
rect 16764 17604 16816 17610
rect 16764 17546 16816 17552
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16672 17264 16724 17270
rect 16672 17206 16724 17212
rect 16580 17128 16632 17134
rect 16578 17096 16580 17105
rect 16632 17096 16634 17105
rect 16578 17031 16634 17040
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16486 15872 16542 15881
rect 16486 15807 16542 15816
rect 16394 15736 16450 15745
rect 16394 15671 16450 15680
rect 16302 13016 16358 13025
rect 16302 12951 16358 12960
rect 16408 12850 16436 15671
rect 16500 15201 16528 15807
rect 16486 15192 16542 15201
rect 16486 15127 16542 15136
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16500 12986 16528 14350
rect 16592 13818 16620 16594
rect 16684 16046 16712 17206
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16776 16250 16804 16526
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16868 16153 16896 22320
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 17236 19310 17264 19858
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17236 19145 17264 19246
rect 17222 19136 17278 19145
rect 17222 19071 17278 19080
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 17038 18592 17094 18601
rect 17038 18527 17094 18536
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16854 16144 16910 16153
rect 16854 16079 16910 16088
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16684 14346 16712 15506
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16776 14074 16804 15438
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16592 13790 16712 13818
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16592 13530 16620 13670
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16592 12730 16620 13330
rect 16684 13161 16712 13790
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16670 13152 16726 13161
rect 16670 13087 16726 13096
rect 16684 12986 16712 13087
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16776 12850 16804 13262
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16868 12730 16896 15846
rect 16960 13977 16988 18022
rect 16946 13968 17002 13977
rect 16946 13903 17002 13912
rect 16592 12702 16712 12730
rect 16304 12640 16356 12646
rect 16684 12617 16712 12702
rect 16776 12702 16896 12730
rect 16304 12582 16356 12588
rect 16670 12608 16726 12617
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16224 8401 16252 11698
rect 16316 10577 16344 12582
rect 16670 12543 16726 12552
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16486 12336 16542 12345
rect 16486 12271 16542 12280
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 11694 16436 12038
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16302 10568 16358 10577
rect 16302 10503 16358 10512
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 9178 16344 9318
rect 16408 9178 16436 11086
rect 16500 10674 16528 12271
rect 16592 11694 16620 12378
rect 16776 12209 16804 12702
rect 16762 12200 16818 12209
rect 16762 12135 16818 12144
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16776 11064 16804 12135
rect 16854 11928 16910 11937
rect 16854 11863 16910 11872
rect 16868 11286 16896 11863
rect 16960 11694 16988 13903
rect 17052 13394 17080 18527
rect 17144 16153 17172 18838
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17236 18601 17264 18770
rect 17222 18592 17278 18601
rect 17222 18527 17278 18536
rect 17130 16144 17186 16153
rect 17130 16079 17186 16088
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17052 13297 17080 13330
rect 17038 13288 17094 13297
rect 17038 13223 17094 13232
rect 17144 13025 17172 15846
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17236 14278 17264 14826
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17236 13462 17264 13670
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17130 13016 17186 13025
rect 17130 12951 17186 12960
rect 17236 12782 17264 13126
rect 17224 12776 17276 12782
rect 17038 12744 17094 12753
rect 17224 12718 17276 12724
rect 17038 12679 17040 12688
rect 17092 12679 17094 12688
rect 17040 12650 17092 12656
rect 17328 12594 17356 22320
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17512 17882 17540 19722
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17408 17604 17460 17610
rect 17408 17546 17460 17552
rect 17420 14385 17448 17546
rect 17512 16697 17540 17818
rect 17498 16688 17554 16697
rect 17498 16623 17554 16632
rect 17696 16425 17724 22320
rect 18064 19802 18092 22320
rect 18432 20074 18460 22320
rect 18602 21448 18658 21457
rect 18602 21383 18658 21392
rect 18432 20046 18552 20074
rect 17788 19774 18092 19802
rect 17788 19174 17816 19774
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18524 19496 18552 20046
rect 18432 19468 18552 19496
rect 18142 19408 18198 19417
rect 18142 19343 18198 19352
rect 18156 19310 18184 19343
rect 17960 19304 18012 19310
rect 17880 19264 17960 19292
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17788 18193 17816 18770
rect 17774 18184 17830 18193
rect 17774 18119 17830 18128
rect 17880 18068 17908 19264
rect 17960 19246 18012 19252
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18432 18986 18460 19468
rect 18616 19378 18644 21383
rect 18694 21040 18750 21049
rect 18694 20975 18750 20984
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18708 19258 18736 20975
rect 18800 19922 18828 22320
rect 19168 20754 19196 22320
rect 19246 22264 19302 22273
rect 19246 22199 19302 22208
rect 19076 20726 19196 20754
rect 19076 20058 19104 20726
rect 19154 20632 19210 20641
rect 19154 20567 19210 20576
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 19168 19990 19196 20567
rect 19156 19984 19208 19990
rect 19156 19926 19208 19932
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18524 19242 18736 19258
rect 18512 19236 18736 19242
rect 18564 19230 18736 19236
rect 18512 19178 18564 19184
rect 18432 18958 18644 18986
rect 18144 18896 18196 18902
rect 18142 18864 18144 18873
rect 18196 18864 18198 18873
rect 18142 18799 18198 18808
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 18329 18000 18566
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18512 18352 18564 18358
rect 17958 18320 18014 18329
rect 18512 18294 18564 18300
rect 17958 18255 18014 18264
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18432 18086 18460 18158
rect 17788 18040 17908 18068
rect 18420 18080 18472 18086
rect 18418 18048 18420 18057
rect 18472 18048 18474 18057
rect 17788 16658 17816 18040
rect 18418 17983 18474 17992
rect 18524 17513 18552 18294
rect 18616 18222 18644 18958
rect 18696 18828 18748 18834
rect 18800 18816 18828 19858
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18748 18788 18828 18816
rect 18696 18770 18748 18776
rect 18708 18426 18736 18770
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18892 17921 18920 19654
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19168 19417 19196 19450
rect 19154 19408 19210 19417
rect 18972 19372 19024 19378
rect 19154 19343 19210 19352
rect 18972 19314 19024 19320
rect 18984 19281 19012 19314
rect 18970 19272 19026 19281
rect 18970 19207 19026 19216
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18984 18737 19012 19110
rect 19260 18902 19288 22199
rect 19536 20670 19564 22320
rect 19524 20664 19576 20670
rect 19524 20606 19576 20612
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19352 20233 19380 20538
rect 19338 20224 19394 20233
rect 19338 20159 19394 20168
rect 19352 19378 19380 20159
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19720 19825 19748 19858
rect 19706 19816 19762 19825
rect 19706 19751 19762 19760
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 19352 18834 19380 19314
rect 19524 19236 19576 19242
rect 19524 19178 19576 19184
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19248 18760 19300 18766
rect 18970 18728 19026 18737
rect 19248 18702 19300 18708
rect 18970 18663 19026 18672
rect 18972 18624 19024 18630
rect 19260 18601 19288 18702
rect 18972 18566 19024 18572
rect 19246 18592 19302 18601
rect 18878 17912 18934 17921
rect 18878 17847 18934 17856
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18510 17504 18566 17513
rect 18116 17436 18412 17456
rect 18510 17439 18566 17448
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 17960 16992 18012 16998
rect 18420 16992 18472 16998
rect 17960 16934 18012 16940
rect 18326 16960 18382 16969
rect 17972 16697 18000 16934
rect 18420 16934 18472 16940
rect 18326 16895 18382 16904
rect 18340 16794 18368 16895
rect 18432 16833 18460 16934
rect 18418 16824 18474 16833
rect 18328 16788 18380 16794
rect 18418 16759 18474 16768
rect 18328 16730 18380 16736
rect 18052 16720 18104 16726
rect 17958 16688 18014 16697
rect 17776 16652 17828 16658
rect 18052 16662 18104 16668
rect 17958 16623 18014 16632
rect 17776 16594 17828 16600
rect 17682 16416 17738 16425
rect 17682 16351 17738 16360
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17512 14929 17540 15098
rect 17498 14920 17554 14929
rect 17498 14855 17554 14864
rect 17604 14804 17632 16186
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17512 14776 17632 14804
rect 17406 14376 17462 14385
rect 17406 14311 17462 14320
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17420 13938 17448 14214
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17420 13326 17448 13874
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17512 13190 17540 14776
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17604 13870 17632 14418
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17500 12708 17552 12714
rect 17500 12650 17552 12656
rect 17052 12566 17356 12594
rect 17406 12608 17462 12617
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16776 11036 16988 11064
rect 16672 11008 16724 11014
rect 16672 10950 16724 10956
rect 16762 10976 16818 10985
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16500 9926 16528 9998
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16500 9450 16528 9862
rect 16684 9450 16712 10950
rect 16762 10911 16818 10920
rect 16488 9444 16540 9450
rect 16488 9386 16540 9392
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16394 9072 16450 9081
rect 16394 9007 16396 9016
rect 16448 9007 16450 9016
rect 16396 8978 16448 8984
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16210 8392 16266 8401
rect 16210 8327 16266 8336
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 16224 7410 16252 7754
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16316 7290 16344 8298
rect 16408 7546 16436 8842
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16224 7262 16344 7290
rect 16224 7206 16252 7262
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 5914 16252 7142
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16316 6662 16344 6802
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16316 5098 16344 6598
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16408 5370 16436 5714
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16304 5092 16356 5098
rect 16304 5034 16356 5040
rect 16408 4690 16436 5306
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 15842 3159 15898 3168
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 15672 2774 15884 2802
rect 14832 1896 14884 1902
rect 14832 1838 14884 1844
rect 15476 1896 15528 1902
rect 15476 1838 15528 1844
rect 15476 1760 15528 1766
rect 15476 1702 15528 1708
rect 14568 1414 14780 1442
rect 14372 1284 14424 1290
rect 14372 1226 14424 1232
rect 14384 480 14412 1226
rect 14752 480 14780 1414
rect 15108 1420 15160 1426
rect 15108 1362 15160 1368
rect 15120 480 15148 1362
rect 15488 480 15516 1702
rect 15856 480 15884 2774
rect 16224 480 16252 4422
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16408 3602 16436 4082
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16408 3058 16436 3538
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16302 2680 16358 2689
rect 16302 2615 16304 2624
rect 16356 2615 16358 2624
rect 16304 2586 16356 2592
rect 16500 2446 16528 9386
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16592 4826 16620 8978
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16592 3670 16620 4558
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 16684 2650 16712 8774
rect 16776 2990 16804 10911
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16868 10062 16896 10610
rect 16960 10606 16988 11036
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16960 10169 16988 10542
rect 16946 10160 17002 10169
rect 16946 10095 17002 10104
rect 16856 10056 16908 10062
rect 16948 10056 17000 10062
rect 16856 9998 16908 10004
rect 16946 10024 16948 10033
rect 17000 10024 17002 10033
rect 16946 9959 17002 9968
rect 17052 9908 17080 12566
rect 17406 12543 17462 12552
rect 17224 12368 17276 12374
rect 17224 12310 17276 12316
rect 17132 11552 17184 11558
rect 17236 11540 17264 12310
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17184 11512 17264 11540
rect 17132 11494 17184 11500
rect 17144 11150 17172 11494
rect 17224 11212 17276 11218
rect 17224 11154 17276 11160
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17144 10674 17172 11086
rect 17236 10810 17264 11154
rect 17328 11082 17356 11698
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17144 10526 17356 10554
rect 17144 9926 17172 10526
rect 17328 10470 17356 10526
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 16868 9880 17080 9908
rect 17132 9920 17184 9926
rect 16868 6905 16896 9880
rect 17132 9862 17184 9868
rect 17132 9648 17184 9654
rect 17130 9616 17132 9625
rect 17184 9616 17186 9625
rect 17130 9551 17186 9560
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16960 8537 16988 8978
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 16946 8528 17002 8537
rect 16946 8463 17002 8472
rect 16946 8392 17002 8401
rect 17052 8362 17080 8910
rect 17144 8430 17172 9551
rect 17236 8566 17264 10406
rect 17420 10282 17448 12543
rect 17328 10254 17448 10282
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 16946 8327 17002 8336
rect 17040 8356 17092 8362
rect 16854 6896 16910 6905
rect 16854 6831 16910 6840
rect 16960 6633 16988 8327
rect 17040 8298 17092 8304
rect 17038 8256 17094 8265
rect 17038 8191 17094 8200
rect 17052 7954 17080 8191
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17038 7712 17094 7721
rect 17038 7647 17094 7656
rect 17052 6798 17080 7647
rect 17236 6905 17264 7890
rect 17222 6896 17278 6905
rect 17222 6831 17278 6840
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 16946 6624 17002 6633
rect 16946 6559 17002 6568
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16868 3534 16896 4218
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16868 2990 16896 3470
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16856 2984 16908 2990
rect 16856 2926 16908 2932
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16776 1358 16804 2926
rect 16764 1352 16816 1358
rect 16764 1294 16816 1300
rect 16580 1148 16632 1154
rect 16580 1090 16632 1096
rect 16592 480 16620 1090
rect 16960 480 16988 5238
rect 17236 5166 17264 6831
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 17144 4214 17172 4626
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 17052 2009 17080 4150
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17144 3194 17172 3878
rect 17328 3602 17356 10254
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17420 9178 17448 10066
rect 17512 9518 17540 12650
rect 17604 12442 17632 13670
rect 17696 13530 17724 15506
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17682 13288 17738 13297
rect 17682 13223 17738 13232
rect 17696 12918 17724 13223
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17604 10554 17632 12378
rect 17696 10849 17724 12650
rect 17788 11830 17816 16594
rect 18064 16561 18092 16662
rect 18050 16552 18106 16561
rect 18050 16487 18106 16496
rect 18616 16454 18644 17546
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18892 17377 18920 17478
rect 18878 17368 18934 17377
rect 18878 17303 18934 17312
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18788 16516 18840 16522
rect 18788 16458 18840 16464
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18510 16144 18566 16153
rect 18800 16114 18828 16458
rect 18510 16079 18566 16088
rect 18788 16108 18840 16114
rect 17960 15972 18012 15978
rect 18012 15932 18092 15960
rect 17960 15914 18012 15920
rect 18064 15638 18092 15932
rect 18524 15910 18552 16079
rect 18788 16050 18840 16056
rect 18144 15904 18196 15910
rect 18142 15872 18144 15881
rect 18512 15904 18564 15910
rect 18196 15872 18198 15881
rect 18512 15846 18564 15852
rect 18142 15807 18198 15816
rect 18326 15736 18382 15745
rect 18236 15700 18288 15706
rect 18800 15706 18828 16050
rect 18326 15671 18328 15680
rect 18236 15642 18288 15648
rect 18380 15671 18382 15680
rect 18788 15700 18840 15706
rect 18328 15642 18380 15648
rect 18788 15642 18840 15648
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 18052 15632 18104 15638
rect 18052 15574 18104 15580
rect 17868 15496 17920 15502
rect 17972 15473 18000 15574
rect 17868 15438 17920 15444
rect 17958 15464 18014 15473
rect 17880 15162 17908 15438
rect 17958 15399 18014 15408
rect 18248 15416 18276 15642
rect 18696 15632 18748 15638
rect 18696 15574 18748 15580
rect 18328 15564 18380 15570
rect 18380 15524 18644 15552
rect 18328 15506 18380 15512
rect 18248 15388 18552 15416
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17880 14550 17908 15098
rect 17972 14958 18000 15302
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18328 15088 18380 15094
rect 18050 15056 18106 15065
rect 18328 15030 18380 15036
rect 18050 14991 18106 15000
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17868 14544 17920 14550
rect 17868 14486 17920 14492
rect 17972 13954 18000 14758
rect 18064 14414 18092 14991
rect 18340 14521 18368 15030
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18432 14618 18460 14962
rect 18524 14958 18552 15388
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18616 14618 18644 15524
rect 18708 14872 18736 15574
rect 18708 14844 18828 14872
rect 18694 14784 18750 14793
rect 18694 14719 18750 14728
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18142 14512 18198 14521
rect 18142 14447 18198 14456
rect 18326 14512 18382 14521
rect 18326 14447 18382 14456
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18156 14346 18184 14447
rect 18432 14362 18460 14554
rect 18708 14482 18736 14719
rect 18800 14550 18828 14844
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18694 14376 18750 14385
rect 18144 14340 18196 14346
rect 18432 14334 18552 14362
rect 18144 14282 18196 14288
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18524 13954 18552 14334
rect 18694 14311 18750 14320
rect 18788 14340 18840 14346
rect 18708 14074 18736 14311
rect 18788 14282 18840 14288
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 17880 13926 18000 13954
rect 18340 13926 18552 13954
rect 17880 12594 17908 13926
rect 18340 13870 18368 13926
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 17972 12866 18000 13806
rect 18800 13802 18828 14282
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 18892 13705 18920 17138
rect 18984 16726 19012 18566
rect 19246 18527 19302 18536
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 19168 17338 19196 17682
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 19076 17218 19104 17274
rect 19076 17190 19196 17218
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18984 14657 19012 16390
rect 18970 14648 19026 14657
rect 18970 14583 19026 14592
rect 18878 13696 18934 13705
rect 18878 13631 18934 13640
rect 18050 13560 18106 13569
rect 18050 13495 18106 13504
rect 18064 13462 18092 13495
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 18144 13456 18196 13462
rect 18144 13398 18196 13404
rect 18604 13456 18656 13462
rect 18604 13398 18656 13404
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18156 13172 18184 13398
rect 18420 13252 18472 13258
rect 18472 13212 18552 13240
rect 18420 13194 18472 13200
rect 18053 13144 18184 13172
rect 18524 13161 18552 13212
rect 18510 13152 18566 13161
rect 18053 12968 18081 13144
rect 18116 13084 18412 13104
rect 18510 13087 18566 13096
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18053 12940 18184 12968
rect 17972 12838 18092 12866
rect 17880 12566 18000 12594
rect 17866 12472 17922 12481
rect 17866 12407 17922 12416
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 17788 11286 17816 11630
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17682 10840 17738 10849
rect 17682 10775 17738 10784
rect 17604 10526 17816 10554
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17604 10130 17632 10406
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17590 9888 17646 9897
rect 17590 9823 17646 9832
rect 17604 9722 17632 9823
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17592 9444 17644 9450
rect 17592 9386 17644 9392
rect 17604 9353 17632 9386
rect 17590 9344 17646 9353
rect 17590 9279 17646 9288
rect 17696 9194 17724 10202
rect 17788 9994 17816 10526
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17788 9704 17816 9930
rect 17880 9897 17908 12407
rect 17972 11694 18000 12566
rect 18064 12306 18092 12838
rect 18156 12646 18184 12940
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 18432 12084 18460 12582
rect 18524 12374 18552 12718
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18510 12200 18566 12209
rect 18510 12135 18566 12144
rect 18053 12056 18460 12084
rect 18053 11880 18081 12056
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18053 11852 18092 11880
rect 17960 11688 18012 11694
rect 18064 11665 18092 11852
rect 17960 11630 18012 11636
rect 18050 11656 18106 11665
rect 18050 11591 18106 11600
rect 18418 11520 18474 11529
rect 18418 11455 18474 11464
rect 18432 11354 18460 11455
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17866 9888 17922 9897
rect 17866 9823 17922 9832
rect 17972 9722 18000 11018
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18052 10532 18104 10538
rect 18052 10474 18104 10480
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 18064 10033 18092 10474
rect 18142 10432 18198 10441
rect 18142 10367 18198 10376
rect 18156 10266 18184 10367
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18142 10160 18198 10169
rect 18142 10095 18144 10104
rect 18196 10095 18198 10104
rect 18144 10066 18196 10072
rect 18050 10024 18106 10033
rect 18050 9959 18106 9968
rect 18248 9908 18276 10474
rect 18053 9880 18276 9908
rect 17960 9716 18012 9722
rect 17788 9676 17908 9704
rect 17880 9586 17908 9676
rect 18053 9704 18081 9880
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18053 9676 18092 9704
rect 17960 9658 18012 9664
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17512 9166 17724 9194
rect 17512 7732 17540 9166
rect 17788 9042 17816 9522
rect 18064 9042 18092 9676
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 17420 7704 17540 7732
rect 17420 6769 17448 7704
rect 17498 7576 17554 7585
rect 17498 7511 17554 7520
rect 17512 7342 17540 7511
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 17500 6792 17552 6798
rect 17406 6760 17462 6769
rect 17500 6734 17552 6740
rect 17406 6695 17462 6704
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 6322 17448 6598
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17512 5778 17540 6734
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17512 5370 17540 5714
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17498 5264 17554 5273
rect 17498 5199 17554 5208
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17420 4593 17448 5102
rect 17406 4584 17462 4593
rect 17406 4519 17462 4528
rect 17408 4004 17460 4010
rect 17408 3946 17460 3952
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17420 3398 17448 3946
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17406 3224 17462 3233
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17224 3188 17276 3194
rect 17406 3159 17462 3168
rect 17224 3130 17276 3136
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17144 2650 17172 2994
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17236 2496 17264 3130
rect 17420 2990 17448 3159
rect 17512 3058 17540 5199
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17498 2816 17554 2825
rect 17498 2751 17554 2760
rect 17512 2650 17540 2751
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17604 2553 17632 8978
rect 17960 8968 18012 8974
rect 17880 8928 17960 8956
rect 17880 8498 17908 8928
rect 17960 8910 18012 8916
rect 18064 8820 18092 8978
rect 18524 8922 18552 12135
rect 18616 11898 18644 13398
rect 18800 13297 18828 13398
rect 18972 13320 19024 13326
rect 18786 13288 18842 13297
rect 18972 13262 19024 13268
rect 18786 13223 18842 13232
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18708 13025 18736 13126
rect 18694 13016 18750 13025
rect 18694 12951 18750 12960
rect 18788 12980 18840 12986
rect 18984 12968 19012 13262
rect 18788 12922 18840 12928
rect 18892 12940 19012 12968
rect 18800 12753 18828 12922
rect 18892 12782 18920 12940
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18880 12776 18932 12782
rect 18786 12744 18842 12753
rect 18880 12718 18932 12724
rect 18786 12679 18842 12688
rect 18694 12608 18750 12617
rect 18694 12543 18750 12552
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18708 11200 18736 12543
rect 18788 12368 18840 12374
rect 18788 12310 18840 12316
rect 18616 11172 18736 11200
rect 18616 9353 18644 11172
rect 18800 11150 18828 12310
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18708 10538 18736 11018
rect 18786 10704 18842 10713
rect 18786 10639 18842 10648
rect 18800 10538 18828 10639
rect 18892 10606 18920 12038
rect 18984 11762 19012 12786
rect 19076 12617 19104 17070
rect 19168 17066 19196 17190
rect 19156 17060 19208 17066
rect 19156 17002 19208 17008
rect 19154 16960 19210 16969
rect 19154 16895 19210 16904
rect 19168 16726 19196 16895
rect 19156 16720 19208 16726
rect 19156 16662 19208 16668
rect 19260 16590 19288 17614
rect 19352 17270 19380 18158
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19340 17128 19392 17134
rect 19444 17105 19472 19110
rect 19536 17270 19564 19178
rect 19720 18834 19748 19751
rect 19904 19394 19932 22320
rect 20364 19922 20392 22320
rect 20626 21856 20682 21865
rect 20626 21791 20682 21800
rect 20640 19990 20668 21791
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 19812 19366 19932 19394
rect 19812 19310 19840 19366
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19616 18216 19668 18222
rect 19616 18158 19668 18164
rect 19524 17264 19576 17270
rect 19524 17206 19576 17212
rect 19340 17070 19392 17076
rect 19430 17096 19486 17105
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19260 16425 19288 16526
rect 19246 16416 19302 16425
rect 19246 16351 19302 16360
rect 19352 16266 19380 17070
rect 19430 17031 19486 17040
rect 19432 16992 19484 16998
rect 19628 16946 19656 18158
rect 19720 18154 19748 18770
rect 19708 18148 19760 18154
rect 19708 18090 19760 18096
rect 19800 18148 19852 18154
rect 19800 18090 19852 18096
rect 19708 17264 19760 17270
rect 19708 17206 19760 17212
rect 19432 16934 19484 16940
rect 19168 16238 19380 16266
rect 19168 13682 19196 16238
rect 19248 16176 19300 16182
rect 19246 16144 19248 16153
rect 19300 16144 19302 16153
rect 19246 16079 19302 16088
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19248 16040 19300 16046
rect 19352 16017 19380 16050
rect 19248 15982 19300 15988
rect 19338 16008 19394 16017
rect 19260 15502 19288 15982
rect 19338 15943 19394 15952
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19352 15706 19380 15846
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19246 15328 19302 15337
rect 19246 15263 19302 15272
rect 19260 14550 19288 15263
rect 19444 15042 19472 16934
rect 19352 15014 19472 15042
rect 19536 16918 19656 16946
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 19168 13654 19288 13682
rect 19154 13560 19210 13569
rect 19154 13495 19210 13504
rect 19168 12918 19196 13495
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19156 12640 19208 12646
rect 19062 12608 19118 12617
rect 19156 12582 19208 12588
rect 19062 12543 19118 12552
rect 19064 12368 19116 12374
rect 19064 12310 19116 12316
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 18984 11558 19012 11698
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 18696 10532 18748 10538
rect 18696 10474 18748 10480
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18708 10282 18736 10474
rect 18984 10452 19012 10542
rect 18892 10424 19012 10452
rect 18708 10254 18828 10282
rect 18800 10198 18828 10254
rect 18696 10192 18748 10198
rect 18696 10134 18748 10140
rect 18788 10192 18840 10198
rect 18788 10134 18840 10140
rect 18602 9344 18658 9353
rect 18602 9279 18658 9288
rect 18602 9072 18658 9081
rect 18602 9007 18604 9016
rect 18656 9007 18658 9016
rect 18604 8978 18656 8984
rect 18524 8894 18644 8922
rect 17958 8800 18014 8809
rect 17958 8735 18014 8744
rect 18053 8792 18092 8820
rect 18510 8800 18566 8809
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17696 7410 17724 7890
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17774 6896 17830 6905
rect 17774 6831 17830 6840
rect 17684 6724 17736 6730
rect 17684 6666 17736 6672
rect 17696 6497 17724 6666
rect 17682 6488 17738 6497
rect 17682 6423 17738 6432
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17696 5574 17724 6258
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 17696 4758 17724 5510
rect 17684 4752 17736 4758
rect 17684 4694 17736 4700
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17696 3942 17724 4082
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17788 3754 17816 6831
rect 17880 6662 17908 8026
rect 17972 8022 18000 8735
rect 18053 8616 18081 8792
rect 18116 8732 18412 8752
rect 18510 8735 18566 8744
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18524 8634 18552 8735
rect 18512 8628 18564 8634
rect 18053 8588 18092 8616
rect 18064 8090 18092 8588
rect 18512 8570 18564 8576
rect 18328 8560 18380 8566
rect 18328 8502 18380 8508
rect 18234 8120 18290 8129
rect 18052 8084 18104 8090
rect 18340 8090 18368 8502
rect 18234 8055 18290 8064
rect 18328 8084 18380 8090
rect 18052 8026 18104 8032
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 18248 7732 18276 8055
rect 18328 8026 18380 8032
rect 18616 7834 18644 8894
rect 18708 8265 18736 10134
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18694 8256 18750 8265
rect 18694 8191 18750 8200
rect 17972 7704 18276 7732
rect 18524 7806 18644 7834
rect 18696 7812 18748 7818
rect 17972 7546 18000 7704
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 18524 7342 18552 7806
rect 18696 7754 18748 7760
rect 18604 7744 18656 7750
rect 18708 7721 18736 7754
rect 18604 7686 18656 7692
rect 18694 7712 18750 7721
rect 18616 7585 18644 7686
rect 18694 7647 18750 7656
rect 18602 7576 18658 7585
rect 18602 7511 18658 7520
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 18064 7002 18092 7142
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 17868 6656 17920 6662
rect 17920 6616 18000 6644
rect 17868 6598 17920 6604
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17880 5642 17908 6054
rect 17972 5914 18000 6616
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18418 6352 18474 6361
rect 18418 6287 18420 6296
rect 18472 6287 18474 6296
rect 18420 6258 18472 6264
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 18064 5914 18092 6054
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 17960 5704 18012 5710
rect 17958 5672 17960 5681
rect 18012 5672 18014 5681
rect 17868 5636 17920 5642
rect 17958 5607 18014 5616
rect 17868 5578 17920 5584
rect 18156 5556 18184 5714
rect 17972 5528 18184 5556
rect 17972 5409 18000 5528
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 17958 5400 18014 5409
rect 18116 5392 18412 5412
rect 17958 5335 18014 5344
rect 17958 5264 18014 5273
rect 17958 5199 18014 5208
rect 17972 4826 18000 5199
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 18524 4758 18552 7278
rect 18616 6905 18644 7511
rect 18694 7440 18750 7449
rect 18694 7375 18750 7384
rect 18602 6896 18658 6905
rect 18602 6831 18658 6840
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18616 6322 18644 6734
rect 18708 6633 18736 7375
rect 18694 6624 18750 6633
rect 18694 6559 18750 6568
rect 18800 6458 18828 9998
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18694 5808 18750 5817
rect 18694 5743 18750 5752
rect 18708 5574 18736 5743
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18800 5234 18828 6258
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18512 4752 18564 4758
rect 18512 4694 18564 4700
rect 18892 4434 18920 10424
rect 19076 10169 19104 12310
rect 19168 11937 19196 12582
rect 19260 12374 19288 13654
rect 19352 12753 19380 15014
rect 19432 14952 19484 14958
rect 19536 14929 19564 16918
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19432 14894 19484 14900
rect 19522 14920 19578 14929
rect 19444 13841 19472 14894
rect 19522 14855 19578 14864
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19430 13832 19486 13841
rect 19430 13767 19486 13776
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19338 12744 19394 12753
rect 19338 12679 19394 12688
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19154 11928 19210 11937
rect 19154 11863 19210 11872
rect 19248 11824 19300 11830
rect 19248 11766 19300 11772
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19168 11354 19196 11494
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19260 11286 19288 11766
rect 19248 11280 19300 11286
rect 19154 11248 19210 11257
rect 19248 11222 19300 11228
rect 19154 11183 19210 11192
rect 19168 10810 19196 11183
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19062 10160 19118 10169
rect 19352 10130 19380 12378
rect 19444 11801 19472 12786
rect 19430 11792 19486 11801
rect 19430 11727 19432 11736
rect 19484 11727 19486 11736
rect 19432 11698 19484 11704
rect 19444 11667 19472 11698
rect 19432 11552 19484 11558
rect 19430 11520 19432 11529
rect 19484 11520 19486 11529
rect 19430 11455 19486 11464
rect 19062 10095 19118 10104
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18984 8634 19012 9862
rect 19064 9648 19116 9654
rect 19168 9636 19196 10066
rect 19248 9648 19300 9654
rect 19168 9608 19248 9636
rect 19064 9590 19116 9596
rect 19248 9590 19300 9596
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18984 6225 19012 8366
rect 18970 6216 19026 6225
rect 18970 6151 19026 6160
rect 18970 5944 19026 5953
rect 18970 5879 19026 5888
rect 18984 5370 19012 5879
rect 18972 5364 19024 5370
rect 18972 5306 19024 5312
rect 18800 4406 18920 4434
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 17696 3726 17816 3754
rect 17960 3732 18012 3738
rect 17696 2650 17724 3726
rect 17960 3674 18012 3680
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17144 2468 17264 2496
rect 17590 2544 17646 2553
rect 17590 2479 17646 2488
rect 17038 2000 17094 2009
rect 17038 1935 17094 1944
rect 17144 1154 17172 2468
rect 17222 2408 17278 2417
rect 17222 2343 17278 2352
rect 17236 2310 17264 2343
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17328 1834 17356 2246
rect 17408 1896 17460 1902
rect 17408 1838 17460 1844
rect 17316 1828 17368 1834
rect 17316 1770 17368 1776
rect 17132 1148 17184 1154
rect 17132 1090 17184 1096
rect 17420 480 17448 1838
rect 17788 480 17816 3062
rect 17880 2972 17908 3334
rect 17972 3108 18000 3674
rect 18616 3618 18644 3674
rect 18524 3590 18644 3618
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18524 3194 18552 3590
rect 18708 3534 18736 3946
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18800 3380 18828 4406
rect 18878 4040 18934 4049
rect 18878 3975 18934 3984
rect 18616 3352 18828 3380
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 17972 3080 18276 3108
rect 17880 2944 18000 2972
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 17880 2446 17908 2586
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 17972 1442 18000 2944
rect 18248 2650 18276 3080
rect 18616 2922 18644 3352
rect 18694 3224 18750 3233
rect 18694 3159 18750 3168
rect 18328 2916 18380 2922
rect 18328 2858 18380 2864
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 18236 2644 18288 2650
rect 18236 2586 18288 2592
rect 18340 2378 18368 2858
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18432 2394 18460 2790
rect 18328 2372 18380 2378
rect 18432 2366 18552 2394
rect 18328 2314 18380 2320
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1414 18184 1442
rect 17960 1352 18012 1358
rect 17960 1294 18012 1300
rect 17972 513 18000 1294
rect 17958 504 18014 513
rect 3422 232 3478 241
rect 3422 167 3478 176
rect 3514 0 3570 480
rect 3882 0 3938 480
rect 4250 0 4306 480
rect 4618 0 4674 480
rect 4986 0 5042 480
rect 5354 0 5410 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7286 0 7342 480
rect 7654 0 7710 480
rect 8022 0 8078 480
rect 8390 0 8446 480
rect 8758 0 8814 480
rect 9126 0 9182 480
rect 9494 0 9550 480
rect 9862 0 9918 480
rect 10230 0 10286 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12530 0 12586 480
rect 12898 0 12954 480
rect 13266 0 13322 480
rect 13634 0 13690 480
rect 14002 0 14058 480
rect 14370 0 14426 480
rect 14738 0 14794 480
rect 15106 0 15162 480
rect 15474 0 15530 480
rect 15842 0 15898 480
rect 16210 0 16266 480
rect 16578 0 16634 480
rect 16946 0 17002 480
rect 17406 0 17462 480
rect 17774 0 17830 480
rect 18156 480 18184 1414
rect 18524 480 18552 2366
rect 18616 2145 18644 2858
rect 18708 2854 18736 3159
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18602 2136 18658 2145
rect 18602 2071 18658 2080
rect 18708 1329 18736 2790
rect 18786 2544 18842 2553
rect 18786 2479 18842 2488
rect 18694 1320 18750 1329
rect 18694 1255 18750 1264
rect 17958 439 18014 448
rect 18142 0 18198 480
rect 18510 0 18566 480
rect 18800 241 18828 2479
rect 18892 480 18920 3975
rect 18984 3058 19012 4422
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18984 2825 19012 2994
rect 18970 2816 19026 2825
rect 18970 2751 19026 2760
rect 18984 2446 19012 2751
rect 19076 2582 19104 9590
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 19168 7546 19196 9454
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 19260 9178 19288 9386
rect 19352 9178 19380 10066
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19260 7721 19288 8570
rect 19352 8498 19380 8910
rect 19444 8906 19472 9318
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 19430 8528 19486 8537
rect 19340 8492 19392 8498
rect 19430 8463 19486 8472
rect 19340 8434 19392 8440
rect 19352 8129 19380 8434
rect 19444 8294 19472 8463
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19338 8120 19394 8129
rect 19338 8055 19394 8064
rect 19536 8072 19564 14758
rect 19628 14550 19656 16730
rect 19720 15609 19748 17206
rect 19812 15638 19840 18090
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19800 15632 19852 15638
rect 19706 15600 19762 15609
rect 19800 15574 19852 15580
rect 19706 15535 19762 15544
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19616 14544 19668 14550
rect 19616 14486 19668 14492
rect 19720 14414 19748 14962
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19614 14240 19670 14249
rect 19614 14175 19670 14184
rect 19628 14074 19656 14175
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19720 13954 19748 14350
rect 19812 14113 19840 15574
rect 19798 14104 19854 14113
rect 19798 14039 19854 14048
rect 19628 13926 19748 13954
rect 19628 12442 19656 13926
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19720 12782 19748 13126
rect 19798 12880 19854 12889
rect 19798 12815 19854 12824
rect 19812 12782 19840 12815
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19904 12594 19932 17614
rect 19996 16046 20024 18906
rect 20076 18080 20128 18086
rect 20076 18022 20128 18028
rect 20088 16794 20116 18022
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 20076 16652 20128 16658
rect 20076 16594 20128 16600
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19982 15600 20038 15609
rect 19982 15535 20038 15544
rect 19996 14929 20024 15535
rect 19982 14920 20038 14929
rect 19982 14855 20038 14864
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19720 12566 19932 12594
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 19614 11928 19670 11937
rect 19614 11863 19670 11872
rect 19628 11626 19656 11863
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19720 9704 19748 12566
rect 19890 12472 19946 12481
rect 19890 12407 19892 12416
rect 19944 12407 19946 12416
rect 19892 12378 19944 12384
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 19890 12200 19946 12209
rect 19812 11014 19840 12174
rect 19890 12135 19946 12144
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19800 10464 19852 10470
rect 19800 10406 19852 10412
rect 19628 9676 19748 9704
rect 19628 9586 19656 9676
rect 19616 9580 19668 9586
rect 19616 9522 19668 9528
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19720 9466 19748 9522
rect 19812 9518 19840 10406
rect 19628 9450 19748 9466
rect 19800 9512 19852 9518
rect 19800 9454 19852 9460
rect 19616 9444 19748 9450
rect 19668 9438 19748 9444
rect 19616 9386 19668 9392
rect 19708 9376 19760 9382
rect 19706 9344 19708 9353
rect 19800 9376 19852 9382
rect 19760 9344 19762 9353
rect 19800 9318 19852 9324
rect 19706 9279 19762 9288
rect 19706 9072 19762 9081
rect 19706 9007 19762 9016
rect 19616 8900 19668 8906
rect 19616 8842 19668 8848
rect 19628 8294 19656 8842
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19536 8044 19656 8072
rect 19340 8016 19392 8022
rect 19338 7984 19340 7993
rect 19392 7984 19394 7993
rect 19338 7919 19394 7928
rect 19246 7712 19302 7721
rect 19246 7647 19302 7656
rect 19628 7546 19656 8044
rect 19720 7698 19748 9007
rect 19812 8838 19840 9318
rect 19904 8974 19932 12135
rect 19996 9042 20024 14758
rect 20088 13938 20116 16594
rect 20180 14793 20208 19110
rect 20364 18698 20392 19858
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20260 17808 20312 17814
rect 20260 17750 20312 17756
rect 20350 17776 20406 17785
rect 20166 14784 20222 14793
rect 20166 14719 20222 14728
rect 20166 14648 20222 14657
rect 20166 14583 20222 14592
rect 20180 14074 20208 14583
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 20074 13016 20130 13025
rect 20074 12951 20130 12960
rect 20088 12442 20116 12951
rect 20180 12918 20208 13262
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 20180 11694 20208 12582
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20166 11112 20222 11121
rect 20166 11047 20222 11056
rect 20180 10674 20208 11047
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20088 10266 20116 10406
rect 20272 10282 20300 17750
rect 20350 17711 20406 17720
rect 20364 16114 20392 17711
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20456 17202 20484 17614
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20364 11286 20392 14962
rect 20548 14906 20576 17070
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20640 16454 20668 16934
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 20732 15745 20760 22320
rect 20824 19310 20852 22607
rect 21086 22320 21142 22800
rect 21454 22320 21510 22800
rect 21822 22320 21878 22800
rect 22190 22320 22246 22800
rect 22558 22320 22614 22800
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20916 18290 20944 18566
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20916 17678 20944 18226
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20916 17202 20944 17614
rect 21100 17354 21128 22320
rect 21468 19786 21496 22320
rect 21836 20058 21864 22320
rect 21824 20052 21876 20058
rect 21824 19994 21876 20000
rect 22204 19854 22232 22320
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 21456 19780 21508 19786
rect 21456 19722 21508 19728
rect 22572 18766 22600 22320
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 21456 17876 21508 17882
rect 21456 17818 21508 17824
rect 21100 17326 21404 17354
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20902 17096 20958 17105
rect 20902 17031 20958 17040
rect 20718 15736 20774 15745
rect 20718 15671 20774 15680
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20456 14878 20576 14906
rect 20456 12986 20484 14878
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20548 14618 20576 14758
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20444 12980 20496 12986
rect 20496 12940 20576 12968
rect 20444 12922 20496 12928
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20180 10254 20300 10282
rect 20364 10266 20392 11222
rect 20352 10260 20404 10266
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19812 8362 19840 8774
rect 19996 8634 20024 8774
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19800 8356 19852 8362
rect 19800 8298 19852 8304
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19720 7670 19840 7698
rect 19706 7576 19762 7585
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19616 7540 19668 7546
rect 19706 7511 19762 7520
rect 19616 7482 19668 7488
rect 19168 7177 19196 7482
rect 19522 7440 19578 7449
rect 19444 7410 19522 7426
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19432 7404 19522 7410
rect 19484 7398 19522 7404
rect 19522 7375 19578 7384
rect 19432 7346 19484 7352
rect 19352 7290 19380 7346
rect 19522 7304 19578 7313
rect 19352 7262 19522 7290
rect 19522 7239 19578 7248
rect 19248 7200 19300 7206
rect 19154 7168 19210 7177
rect 19616 7200 19668 7206
rect 19300 7160 19564 7188
rect 19248 7142 19300 7148
rect 19154 7103 19210 7112
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19168 6322 19196 6734
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19260 5794 19288 6802
rect 19352 5914 19380 6938
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19444 6662 19472 6802
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19536 6458 19564 7160
rect 19616 7142 19668 7148
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19444 5914 19472 6122
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19260 5766 19380 5794
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19154 4176 19210 4185
rect 19154 4111 19210 4120
rect 19168 4078 19196 4111
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 19260 2990 19288 4966
rect 19352 4826 19380 5766
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19352 3738 19380 4558
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19338 3224 19394 3233
rect 19444 3194 19472 4626
rect 19628 4282 19656 7142
rect 19720 5642 19748 7511
rect 19812 7410 19840 7670
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19800 7268 19852 7274
rect 19800 7210 19852 7216
rect 19708 5636 19760 5642
rect 19708 5578 19760 5584
rect 19812 5234 19840 7210
rect 19904 5409 19932 8026
rect 19996 7954 20024 8434
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19982 7848 20038 7857
rect 19982 7783 20038 7792
rect 19996 7313 20024 7783
rect 19982 7304 20038 7313
rect 19982 7239 20038 7248
rect 19982 7168 20038 7177
rect 19982 7103 20038 7112
rect 19996 5710 20024 7103
rect 20088 6905 20116 10202
rect 20180 8566 20208 10254
rect 20352 10202 20404 10208
rect 20260 10192 20312 10198
rect 20260 10134 20312 10140
rect 20168 8560 20220 8566
rect 20168 8502 20220 8508
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20074 6896 20130 6905
rect 20074 6831 20130 6840
rect 20180 6769 20208 8026
rect 20166 6760 20222 6769
rect 20166 6695 20168 6704
rect 20220 6695 20222 6704
rect 20168 6666 20220 6672
rect 20168 6180 20220 6186
rect 20168 6122 20220 6128
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 19890 5400 19946 5409
rect 19890 5335 19946 5344
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19800 5228 19852 5234
rect 19800 5170 19852 5176
rect 19892 5092 19944 5098
rect 19892 5034 19944 5040
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19536 3738 19564 4014
rect 19708 4004 19760 4010
rect 19628 3964 19708 3992
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19628 3346 19656 3964
rect 19708 3946 19760 3952
rect 19812 3738 19840 4762
rect 19904 4622 19932 5034
rect 19996 4690 20024 5306
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19892 4616 19944 4622
rect 20088 4570 20116 5510
rect 20180 5370 20208 6122
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 19892 4558 19944 4564
rect 19904 3942 19932 4558
rect 19996 4542 20116 4570
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 19536 3318 19656 3346
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19338 3159 19394 3168
rect 19432 3188 19484 3194
rect 19352 2990 19380 3159
rect 19432 3130 19484 3136
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19248 2848 19300 2854
rect 19154 2816 19210 2825
rect 19300 2808 19380 2836
rect 19248 2790 19300 2796
rect 19154 2751 19210 2760
rect 19168 2650 19196 2751
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 19064 2576 19116 2582
rect 19064 2518 19116 2524
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 18970 2272 19026 2281
rect 18970 2207 19026 2216
rect 18984 2038 19012 2207
rect 18972 2032 19024 2038
rect 19260 2009 19288 2518
rect 18972 1974 19024 1980
rect 19246 2000 19302 2009
rect 19246 1935 19302 1944
rect 19352 1850 19380 2808
rect 19536 2650 19564 3318
rect 19616 3188 19668 3194
rect 19616 3130 19668 3136
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 19260 1822 19380 1850
rect 19260 480 19288 1822
rect 19628 480 19656 3130
rect 19720 2650 19748 3334
rect 19812 3058 19840 3470
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 19904 2446 19932 3878
rect 19996 2972 20024 4542
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 20088 4078 20116 4422
rect 20180 4214 20208 5306
rect 20168 4208 20220 4214
rect 20168 4150 20220 4156
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 20088 3126 20116 3334
rect 20076 3120 20128 3126
rect 20076 3062 20128 3068
rect 19996 2944 20116 2972
rect 20088 2514 20116 2944
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 19892 2440 19944 2446
rect 20180 2394 20208 3674
rect 19892 2382 19944 2388
rect 19996 2366 20208 2394
rect 19996 480 20024 2366
rect 20272 1970 20300 10134
rect 20350 10024 20406 10033
rect 20350 9959 20406 9968
rect 20364 8022 20392 9959
rect 20456 8430 20484 12242
rect 20548 10606 20576 12940
rect 20640 11218 20668 15438
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20732 13530 20760 14350
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20718 13424 20774 13433
rect 20718 13359 20774 13368
rect 20732 12918 20760 13359
rect 20720 12912 20772 12918
rect 20720 12854 20772 12860
rect 20824 12730 20852 14894
rect 20916 14074 20944 17031
rect 20994 16280 21050 16289
rect 20994 16215 21050 16224
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20824 12702 20944 12730
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20548 8634 20576 9318
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20640 8498 20668 10610
rect 20732 10198 20760 11494
rect 20720 10192 20772 10198
rect 20720 10134 20772 10140
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20732 9178 20760 9658
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20352 8016 20404 8022
rect 20352 7958 20404 7964
rect 20536 7948 20588 7954
rect 20536 7890 20588 7896
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20364 7478 20392 7822
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20456 6458 20484 6598
rect 20548 6497 20576 7890
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 20732 6633 20760 7754
rect 20824 7449 20852 12582
rect 20916 10606 20944 12702
rect 21008 11898 21036 16215
rect 21178 15872 21234 15881
rect 21178 15807 21234 15816
rect 21086 13968 21142 13977
rect 21086 13903 21142 13912
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21100 11830 21128 13903
rect 21088 11824 21140 11830
rect 21088 11766 21140 11772
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 21086 11656 21142 11665
rect 20904 10600 20956 10606
rect 20904 10542 20956 10548
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20916 9450 20944 9998
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 20810 7440 20866 7449
rect 20810 7375 20866 7384
rect 21008 7041 21036 11630
rect 21086 11591 21142 11600
rect 21100 8673 21128 11591
rect 21192 10810 21220 15807
rect 21270 11248 21326 11257
rect 21270 11183 21326 11192
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 21284 8838 21312 11183
rect 21376 8945 21404 17326
rect 21468 12442 21496 17818
rect 21732 17604 21784 17610
rect 21732 17546 21784 17552
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21456 12436 21508 12442
rect 21456 12378 21508 12384
rect 21362 8936 21418 8945
rect 21362 8871 21418 8880
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21086 8664 21142 8673
rect 21086 8599 21142 8608
rect 21088 8016 21140 8022
rect 21088 7958 21140 7964
rect 21100 7342 21128 7958
rect 21088 7336 21140 7342
rect 21088 7278 21140 7284
rect 21652 7206 21680 17002
rect 21640 7200 21692 7206
rect 21640 7142 21692 7148
rect 20994 7032 21050 7041
rect 21744 7018 21772 17546
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 20994 6967 21050 6976
rect 21100 6990 21772 7018
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20718 6624 20774 6633
rect 20718 6559 20774 6568
rect 20534 6488 20590 6497
rect 20444 6452 20496 6458
rect 20534 6423 20590 6432
rect 20444 6394 20496 6400
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20260 1964 20312 1970
rect 20260 1906 20312 1912
rect 20364 480 20392 4558
rect 20456 4282 20484 5102
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20456 3194 20484 3878
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20444 2984 20496 2990
rect 20442 2952 20444 2961
rect 20496 2952 20498 2961
rect 20548 2922 20576 4558
rect 20732 3777 20760 6559
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20824 4078 20852 4626
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20718 3768 20774 3777
rect 20718 3703 20774 3712
rect 20718 3496 20774 3505
rect 20718 3431 20774 3440
rect 20732 3194 20760 3431
rect 20810 3224 20866 3233
rect 20720 3188 20772 3194
rect 20810 3159 20866 3168
rect 20720 3130 20772 3136
rect 20442 2887 20498 2896
rect 20536 2916 20588 2922
rect 20536 2858 20588 2864
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20640 2582 20668 2858
rect 20628 2576 20680 2582
rect 20628 2518 20680 2524
rect 20824 2258 20852 3159
rect 20732 2230 20852 2258
rect 20732 480 20760 2230
rect 20916 2106 20944 6734
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 21008 2553 21036 5714
rect 20994 2544 21050 2553
rect 20994 2479 21050 2488
rect 20904 2100 20956 2106
rect 20904 2042 20956 2048
rect 21100 480 21128 6990
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21180 4752 21232 4758
rect 21180 4694 21232 4700
rect 21192 1737 21220 4694
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 21178 1728 21234 1737
rect 21178 1663 21234 1672
rect 21468 480 21496 2314
rect 21836 480 21864 6054
rect 21928 3369 21956 10406
rect 21914 3360 21970 3369
rect 21914 3295 21970 3304
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 22204 480 22232 2858
rect 22572 480 22600 2926
rect 18786 232 18842 241
rect 18786 167 18842 176
rect 18878 0 18934 480
rect 19246 0 19302 480
rect 19614 0 19670 480
rect 19982 0 20038 480
rect 20350 0 20406 480
rect 20718 0 20774 480
rect 21086 0 21142 480
rect 21454 0 21510 480
rect 21822 0 21878 480
rect 22190 0 22246 480
rect 22558 0 22614 480
<< via2 >>
rect 20810 22616 20866 22672
rect 1950 20984 2006 21040
rect 1858 20576 1914 20632
rect 1950 19352 2006 19408
rect 2318 19916 2374 19952
rect 2318 19896 2320 19916
rect 2320 19896 2372 19916
rect 2372 19896 2374 19916
rect 2778 19796 2780 19816
rect 2780 19796 2832 19816
rect 2832 19796 2834 19816
rect 2778 19760 2834 19796
rect 1950 18672 2006 18728
rect 1674 17992 1730 18048
rect 1490 17856 1546 17912
rect 1858 17720 1914 17776
rect 1766 17584 1822 17640
rect 1582 17040 1638 17096
rect 1582 14320 1638 14376
rect 1674 13504 1730 13560
rect 1490 12824 1546 12880
rect 1582 11192 1638 11248
rect 1950 12688 2006 12744
rect 1858 10512 1914 10568
rect 1858 9288 1914 9344
rect 1674 7384 1730 7440
rect 2410 16088 2466 16144
rect 3238 18264 3294 18320
rect 3146 18128 3202 18184
rect 2778 17448 2834 17504
rect 3330 18128 3386 18184
rect 3882 22208 3938 22264
rect 3698 21800 3754 21856
rect 3882 20168 3938 20224
rect 3882 18808 3938 18864
rect 3606 17992 3662 18048
rect 2778 17040 2834 17096
rect 2594 15544 2650 15600
rect 2778 16224 2834 16280
rect 2686 14320 2742 14376
rect 2042 9152 2098 9208
rect 3422 17176 3478 17232
rect 4066 21392 4122 21448
rect 4710 19760 4766 19816
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4066 19352 4122 19408
rect 4434 19216 4490 19272
rect 4342 19080 4398 19136
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4434 18300 4436 18320
rect 4436 18300 4488 18320
rect 4488 18300 4490 18320
rect 4434 18264 4490 18300
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 3974 16904 4030 16960
rect 3238 15680 3294 15736
rect 2870 13776 2926 13832
rect 2870 13096 2926 13152
rect 3054 12280 3110 12336
rect 3330 14864 3386 14920
rect 3514 15952 3570 16008
rect 4342 16668 4344 16688
rect 4344 16668 4396 16688
rect 4396 16668 4398 16688
rect 4342 16632 4398 16668
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4066 15816 4122 15872
rect 3974 15408 4030 15464
rect 3790 14728 3846 14784
rect 3238 12008 3294 12064
rect 3146 11872 3202 11928
rect 3054 9152 3110 9208
rect 2226 6840 2282 6896
rect 2410 3848 2466 3904
rect 2410 3304 2466 3360
rect 2042 2488 2098 2544
rect 2870 3440 2926 3496
rect 2778 2624 2834 2680
rect 2778 1672 2834 1728
rect 3606 11600 3662 11656
rect 3146 8472 3202 8528
rect 3698 11464 3754 11520
rect 3698 10784 3754 10840
rect 3882 12552 3938 12608
rect 4066 15136 4122 15192
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4250 13912 4306 13968
rect 3974 12144 4030 12200
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 3422 7792 3478 7848
rect 3330 6160 3386 6216
rect 3146 4120 3202 4176
rect 4066 10376 4122 10432
rect 5170 18944 5226 19000
rect 5538 19352 5594 19408
rect 5262 17720 5318 17776
rect 5262 15952 5318 16008
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4710 9424 4766 9480
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4066 7692 4068 7712
rect 4068 7692 4120 7712
rect 4120 7692 4122 7712
rect 4710 8356 4766 8392
rect 4710 8336 4712 8356
rect 4712 8336 4764 8356
rect 4764 8336 4766 8356
rect 4066 7656 4122 7692
rect 3606 6704 3662 6760
rect 3238 2896 3294 2952
rect 3054 448 3110 504
rect 3330 856 3386 912
rect 3606 2624 3662 2680
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4618 6316 4674 6352
rect 4618 6296 4620 6316
rect 4620 6296 4672 6316
rect 4672 6296 4674 6316
rect 4066 5616 4122 5672
rect 3974 4936 4030 4992
rect 3882 2896 3938 2952
rect 3698 2080 3754 2136
rect 4066 3984 4122 4040
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4894 12960 4950 13016
rect 4894 10784 4950 10840
rect 4894 6332 4896 6352
rect 4896 6332 4948 6352
rect 4948 6332 4950 6352
rect 4894 6296 4950 6332
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4434 3984 4490 4040
rect 4250 3732 4306 3768
rect 4250 3712 4252 3732
rect 4252 3712 4304 3732
rect 4304 3712 4306 3732
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 3974 1264 4030 1320
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 5170 12552 5226 12608
rect 5170 12280 5226 12336
rect 5078 11056 5134 11112
rect 5630 15544 5686 15600
rect 5446 14592 5502 14648
rect 5630 14320 5686 14376
rect 5262 10920 5318 10976
rect 5630 13524 5686 13560
rect 5630 13504 5632 13524
rect 5632 13504 5684 13524
rect 5684 13504 5686 13524
rect 5722 13368 5778 13424
rect 6090 19760 6146 19816
rect 6458 18536 6514 18592
rect 6090 17604 6146 17640
rect 6090 17584 6092 17604
rect 6092 17584 6144 17604
rect 6144 17584 6146 17604
rect 6090 17040 6146 17096
rect 6090 14592 6146 14648
rect 6090 14320 6146 14376
rect 5998 13504 6054 13560
rect 5906 11736 5962 11792
rect 5722 9968 5778 10024
rect 5170 9016 5226 9072
rect 5078 8880 5134 8936
rect 5170 8336 5226 8392
rect 5354 8472 5410 8528
rect 5262 6024 5318 6080
rect 5262 4120 5318 4176
rect 5630 8744 5686 8800
rect 5906 10512 5962 10568
rect 5906 9424 5962 9480
rect 5538 6976 5594 7032
rect 5538 4800 5594 4856
rect 5538 4120 5594 4176
rect 5538 3596 5594 3632
rect 5538 3576 5540 3596
rect 5540 3576 5592 3596
rect 5592 3576 5594 3596
rect 5814 7248 5870 7304
rect 5722 2760 5778 2816
rect 6090 12824 6146 12880
rect 6550 16632 6606 16688
rect 6458 15000 6514 15056
rect 6642 15408 6698 15464
rect 6734 15272 6790 15328
rect 6734 13776 6790 13832
rect 6734 12824 6790 12880
rect 7378 18944 7434 19000
rect 7194 18400 7250 18456
rect 7194 17992 7250 18048
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7562 18944 7618 19000
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 8390 19352 8446 19408
rect 8574 19080 8630 19136
rect 8390 18400 8446 18456
rect 8390 17992 8446 18048
rect 7286 15544 7342 15600
rect 7102 13504 7158 13560
rect 6182 10240 6238 10296
rect 6182 8472 6238 8528
rect 6182 8336 6238 8392
rect 6366 9596 6368 9616
rect 6368 9596 6420 9616
rect 6420 9596 6422 9616
rect 6366 9560 6422 9596
rect 6366 9424 6422 9480
rect 6366 8200 6422 8256
rect 6182 6976 6238 7032
rect 7102 12416 7158 12472
rect 6642 10920 6698 10976
rect 6826 10648 6882 10704
rect 6642 8744 6698 8800
rect 6918 10104 6974 10160
rect 6826 9424 6882 9480
rect 6826 9036 6882 9072
rect 6826 9016 6828 9036
rect 6828 9016 6880 9036
rect 6880 9016 6882 9036
rect 6458 7520 6514 7576
rect 6182 5344 6238 5400
rect 6734 8472 6790 8528
rect 6826 8200 6882 8256
rect 6550 7248 6606 7304
rect 6734 6976 6790 7032
rect 6458 6568 6514 6624
rect 6366 6432 6422 6488
rect 6274 4392 6330 4448
rect 6918 5752 6974 5808
rect 6458 2760 6514 2816
rect 6734 5208 6790 5264
rect 6642 3984 6698 4040
rect 6826 3304 6882 3360
rect 6826 3032 6882 3088
rect 7562 15680 7618 15736
rect 7470 15136 7526 15192
rect 7654 15408 7710 15464
rect 7470 13932 7526 13968
rect 7470 13912 7472 13932
rect 7472 13912 7524 13932
rect 7524 13912 7526 13932
rect 7378 13268 7380 13288
rect 7380 13268 7432 13288
rect 7432 13268 7434 13288
rect 7378 13232 7434 13268
rect 7286 12008 7342 12064
rect 8022 17196 8078 17232
rect 8022 17176 8024 17196
rect 8024 17176 8076 17196
rect 8076 17176 8078 17196
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 8114 15020 8170 15056
rect 8114 15000 8116 15020
rect 8116 15000 8168 15020
rect 8168 15000 8170 15020
rect 8298 15000 8354 15056
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7470 12144 7526 12200
rect 7562 12008 7618 12064
rect 8206 13232 8262 13288
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 8114 12280 8170 12336
rect 7470 11600 7526 11656
rect 7194 10648 7250 10704
rect 7194 9016 7250 9072
rect 7378 8744 7434 8800
rect 8298 12280 8354 12336
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 8114 10124 8170 10160
rect 8114 10104 8116 10124
rect 8116 10104 8168 10124
rect 8168 10104 8170 10124
rect 7470 7384 7526 7440
rect 7102 6024 7158 6080
rect 7286 6568 7342 6624
rect 7286 5888 7342 5944
rect 7102 5208 7158 5264
rect 7286 4528 7342 4584
rect 7194 2352 7250 2408
rect 7654 7692 7656 7712
rect 7656 7692 7708 7712
rect 7708 7692 7710 7712
rect 7654 7656 7710 7692
rect 8206 9832 8262 9888
rect 8758 19896 8814 19952
rect 8666 18264 8722 18320
rect 8482 15544 8538 15600
rect 9034 17992 9090 18048
rect 8942 16632 8998 16688
rect 8850 15952 8906 16008
rect 8758 12416 8814 12472
rect 8574 12008 8630 12064
rect 8574 11872 8630 11928
rect 8666 11056 8722 11112
rect 8482 10784 8538 10840
rect 8298 9288 8354 9344
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 8206 9172 8262 9208
rect 8206 9152 8208 9172
rect 8208 9152 8260 9172
rect 8260 9152 8262 9172
rect 8022 8744 8078 8800
rect 8298 8880 8354 8936
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7654 7112 7710 7168
rect 7562 6976 7618 7032
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 8022 6840 8078 6896
rect 8022 6568 8078 6624
rect 7470 5636 7526 5672
rect 7470 5616 7472 5636
rect 7472 5616 7524 5636
rect 7524 5616 7526 5636
rect 8482 7928 8538 7984
rect 8666 9696 8722 9752
rect 8942 12960 8998 13016
rect 9770 18164 9772 18184
rect 9772 18164 9824 18184
rect 9824 18164 9826 18184
rect 9770 18128 9826 18164
rect 9126 15000 9182 15056
rect 9034 11600 9090 11656
rect 9034 10920 9090 10976
rect 9034 9968 9090 10024
rect 8666 8064 8722 8120
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7562 4936 7618 4992
rect 7562 3848 7618 3904
rect 8298 6024 8354 6080
rect 8666 6568 8722 6624
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 8022 4256 8078 4312
rect 9034 8200 9090 8256
rect 9218 12280 9274 12336
rect 9586 15136 9642 15192
rect 9586 12280 9642 12336
rect 10046 18944 10102 19000
rect 9862 15544 9918 15600
rect 9402 11872 9458 11928
rect 9586 11600 9642 11656
rect 9862 13776 9918 13832
rect 9310 10684 9312 10704
rect 9312 10684 9364 10704
rect 9364 10684 9366 10704
rect 9310 10648 9366 10684
rect 9218 10104 9274 10160
rect 9218 9560 9274 9616
rect 9218 8880 9274 8936
rect 8758 5888 8814 5944
rect 8482 4800 8538 4856
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 8114 3440 8170 3496
rect 7746 3168 7802 3224
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 8022 2488 8078 2544
rect 8482 3032 8538 3088
rect 8666 3848 8722 3904
rect 8482 2896 8538 2952
rect 9494 9016 9550 9072
rect 9954 11328 10010 11384
rect 9954 10512 10010 10568
rect 9862 9832 9918 9888
rect 9862 9424 9918 9480
rect 10690 18128 10746 18184
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 10966 16904 11022 16960
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 10414 15680 10470 15736
rect 10598 15408 10654 15464
rect 10598 13368 10654 13424
rect 10230 12960 10286 13016
rect 10138 12824 10194 12880
rect 10138 12552 10194 12608
rect 10046 9424 10102 9480
rect 10598 12416 10654 12472
rect 10414 12144 10470 12200
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11334 14476 11390 14512
rect 11334 14456 11336 14476
rect 11336 14456 11388 14476
rect 11388 14456 11390 14476
rect 11426 14356 11428 14376
rect 11428 14356 11480 14376
rect 11480 14356 11482 14376
rect 11426 14320 11482 14356
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11150 13912 11206 13968
rect 11518 13676 11520 13696
rect 11520 13676 11572 13696
rect 11572 13676 11574 13696
rect 11518 13640 11574 13676
rect 11058 13096 11114 13152
rect 10414 11600 10470 11656
rect 10322 9968 10378 10024
rect 9862 9016 9918 9072
rect 9310 7112 9366 7168
rect 9218 6996 9274 7032
rect 9218 6976 9220 6996
rect 9220 6976 9272 6996
rect 9272 6976 9274 6996
rect 9126 6432 9182 6488
rect 8942 5772 8998 5808
rect 8942 5752 8944 5772
rect 8944 5752 8996 5772
rect 8996 5752 8998 5772
rect 8942 3576 8998 3632
rect 8942 3440 8998 3496
rect 10046 8744 10102 8800
rect 9862 8064 9918 8120
rect 9862 6432 9918 6488
rect 9402 5752 9458 5808
rect 9770 6160 9826 6216
rect 9218 4800 9274 4856
rect 9126 4256 9182 4312
rect 9310 3848 9366 3904
rect 9034 3032 9090 3088
rect 9494 4800 9550 4856
rect 9126 2624 9182 2680
rect 8942 2488 8998 2544
rect 8758 2216 8814 2272
rect 8942 2080 8998 2136
rect 10414 8880 10470 8936
rect 10322 8608 10378 8664
rect 10414 8356 10470 8392
rect 10414 8336 10416 8356
rect 10416 8336 10468 8356
rect 10468 8336 10470 8356
rect 10874 11328 10930 11384
rect 10782 9696 10838 9752
rect 10506 8064 10562 8120
rect 10322 7792 10378 7848
rect 10598 7792 10654 7848
rect 10138 5072 10194 5128
rect 10046 4528 10102 4584
rect 10322 5072 10378 5128
rect 10322 4528 10378 4584
rect 10138 3476 10140 3496
rect 10140 3476 10192 3496
rect 10192 3476 10194 3496
rect 10138 3440 10194 3476
rect 10138 3032 10194 3088
rect 10690 7520 10746 7576
rect 10690 6976 10746 7032
rect 10690 6568 10746 6624
rect 10690 6024 10746 6080
rect 10690 5480 10746 5536
rect 10690 4256 10746 4312
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11518 12824 11574 12880
rect 11794 17076 11796 17096
rect 11796 17076 11848 17096
rect 11848 17076 11850 17096
rect 11794 17040 11850 17076
rect 12070 16768 12126 16824
rect 11978 16088 12034 16144
rect 11518 12280 11574 12336
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11150 10512 11206 10568
rect 11978 13096 12034 13152
rect 11886 12552 11942 12608
rect 11518 10376 11574 10432
rect 11058 8608 11114 8664
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11334 9424 11390 9480
rect 11702 9832 11758 9888
rect 11794 9696 11850 9752
rect 11702 9444 11758 9480
rect 12254 19080 12310 19136
rect 12530 18028 12532 18048
rect 12532 18028 12584 18048
rect 12584 18028 12586 18048
rect 12530 17992 12586 18028
rect 12714 17060 12770 17096
rect 13266 18944 13322 19000
rect 12714 17040 12716 17060
rect 12716 17040 12768 17060
rect 12768 17040 12770 17060
rect 13082 16904 13138 16960
rect 13450 18536 13506 18592
rect 13910 18944 13966 19000
rect 13726 18264 13782 18320
rect 13542 17720 13598 17776
rect 13358 16768 13414 16824
rect 12714 14864 12770 14920
rect 12438 14184 12494 14240
rect 12162 12436 12218 12472
rect 12162 12416 12164 12436
rect 12164 12416 12216 12436
rect 12216 12416 12218 12436
rect 12162 11600 12218 11656
rect 12162 11464 12218 11520
rect 12162 10784 12218 10840
rect 11702 9424 11704 9444
rect 11704 9424 11756 9444
rect 11756 9424 11758 9444
rect 12070 10240 12126 10296
rect 12070 9968 12126 10024
rect 12898 14320 12954 14376
rect 12438 10260 12494 10296
rect 12438 10240 12440 10260
rect 12440 10240 12492 10260
rect 12492 10240 12494 10260
rect 12622 10240 12678 10296
rect 11334 8880 11390 8936
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11242 8064 11298 8120
rect 11426 8336 11482 8392
rect 11058 7656 11114 7712
rect 10874 5344 10930 5400
rect 10506 3304 10562 3360
rect 10966 3032 11022 3088
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11150 7112 11206 7168
rect 11242 6996 11298 7032
rect 11242 6976 11244 6996
rect 11244 6976 11296 6996
rect 11296 6976 11298 6996
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11518 4800 11574 4856
rect 11702 5480 11758 5536
rect 11886 7792 11942 7848
rect 11886 6568 11942 6624
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 12530 8608 12586 8664
rect 12438 8472 12494 8528
rect 12530 7112 12586 7168
rect 13082 13504 13138 13560
rect 12990 12960 13046 13016
rect 13542 16224 13598 16280
rect 13358 12280 13414 12336
rect 13082 11872 13138 11928
rect 13358 11872 13414 11928
rect 13266 11192 13322 11248
rect 12898 9696 12954 9752
rect 12530 6432 12586 6488
rect 12438 5344 12494 5400
rect 12254 5108 12256 5128
rect 12256 5108 12308 5128
rect 12308 5108 12310 5128
rect 12254 5072 12310 5108
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11150 2488 11206 2544
rect 11334 2508 11390 2544
rect 11334 2488 11336 2508
rect 11336 2488 11388 2508
rect 11388 2488 11390 2508
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 11978 3984 12034 4040
rect 12530 4256 12586 4312
rect 12530 3884 12532 3904
rect 12532 3884 12584 3904
rect 12584 3884 12586 3904
rect 12530 3848 12586 3884
rect 12346 2896 12402 2952
rect 12990 8744 13046 8800
rect 13082 8064 13138 8120
rect 12898 7520 12954 7576
rect 12806 6432 12862 6488
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 14370 18128 14426 18184
rect 14278 17856 14334 17912
rect 14186 15952 14242 16008
rect 14094 14356 14096 14376
rect 14096 14356 14148 14376
rect 14148 14356 14150 14376
rect 14094 14320 14150 14356
rect 13726 11872 13782 11928
rect 13726 11212 13782 11248
rect 13726 11192 13728 11212
rect 13728 11192 13780 11212
rect 13780 11192 13782 11212
rect 13726 11056 13782 11112
rect 14094 12280 14150 12336
rect 14002 11736 14058 11792
rect 14094 11328 14150 11384
rect 13818 10648 13874 10704
rect 13634 10240 13690 10296
rect 13542 9696 13598 9752
rect 13358 8744 13414 8800
rect 13634 9016 13690 9072
rect 12898 4972 12900 4992
rect 12900 4972 12952 4992
rect 12952 4972 12954 4992
rect 12898 4936 12954 4972
rect 13174 6024 13230 6080
rect 13082 3052 13138 3088
rect 13082 3032 13084 3052
rect 13084 3032 13136 3052
rect 13136 3032 13138 3052
rect 13358 7520 13414 7576
rect 13358 4664 13414 4720
rect 14186 10376 14242 10432
rect 14370 16904 14426 16960
rect 14370 16652 14426 16688
rect 14370 16632 14372 16652
rect 14372 16632 14424 16652
rect 14424 16632 14426 16652
rect 14370 15000 14426 15056
rect 14922 19352 14978 19408
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14554 18128 14610 18184
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14646 17584 14702 17640
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14370 12824 14426 12880
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 15290 17584 15346 17640
rect 15934 19488 15990 19544
rect 15842 18400 15898 18456
rect 15750 16496 15806 16552
rect 15382 15272 15438 15328
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14922 12960 14978 13016
rect 14462 12552 14518 12608
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14554 11600 14610 11656
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 15198 13776 15254 13832
rect 15290 12960 15346 13016
rect 15106 11872 15162 11928
rect 14370 11056 14426 11112
rect 15106 11192 15162 11248
rect 15014 10920 15070 10976
rect 14370 10104 14426 10160
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14646 10104 14702 10160
rect 13818 8200 13874 8256
rect 13818 7656 13874 7712
rect 13726 7112 13782 7168
rect 14094 7520 14150 7576
rect 14278 8608 14334 8664
rect 14094 6976 14150 7032
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 15750 14320 15806 14376
rect 15750 14184 15806 14240
rect 15658 13504 15714 13560
rect 15658 13232 15714 13288
rect 15750 12960 15806 13016
rect 15566 11464 15622 11520
rect 15474 11328 15530 11384
rect 15014 8608 15070 8664
rect 14462 7112 14518 7168
rect 14370 5888 14426 5944
rect 13726 5616 13782 5672
rect 13634 4120 13690 4176
rect 13542 3440 13598 3496
rect 13910 3848 13966 3904
rect 14002 3576 14058 3632
rect 13910 3440 13966 3496
rect 14002 2760 14058 2816
rect 14462 5752 14518 5808
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 15106 7112 15162 7168
rect 14646 5616 14702 5672
rect 14554 5072 14610 5128
rect 14370 4800 14426 4856
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 15014 4664 15070 4720
rect 14278 3712 14334 3768
rect 16026 17448 16082 17504
rect 16486 19488 16542 19544
rect 16302 18264 16358 18320
rect 16394 17176 16450 17232
rect 16302 16360 16358 16416
rect 15842 11872 15898 11928
rect 15842 11600 15898 11656
rect 15842 11348 15898 11384
rect 15842 11328 15844 11348
rect 15844 11328 15896 11348
rect 15896 11328 15898 11348
rect 15842 9832 15898 9888
rect 15566 8608 15622 8664
rect 15566 8472 15622 8528
rect 15474 7792 15530 7848
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14462 3304 14518 3360
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15382 4664 15438 4720
rect 15658 8200 15714 8256
rect 15658 7928 15714 7984
rect 15750 7656 15806 7712
rect 16026 12416 16082 12472
rect 16026 11328 16082 11384
rect 15934 9560 15990 9616
rect 15934 9152 15990 9208
rect 15934 8880 15990 8936
rect 16026 8336 16082 8392
rect 16026 7520 16082 7576
rect 15750 7112 15806 7168
rect 15934 6976 15990 7032
rect 15842 5480 15898 5536
rect 15842 4800 15898 4856
rect 16026 4664 16082 4720
rect 15842 3168 15898 3224
rect 16210 15852 16212 15872
rect 16212 15852 16264 15872
rect 16264 15852 16266 15872
rect 16210 15816 16266 15852
rect 16210 13776 16266 13832
rect 16578 17076 16580 17096
rect 16580 17076 16632 17096
rect 16632 17076 16634 17096
rect 16578 17040 16634 17076
rect 16486 15816 16542 15872
rect 16394 15680 16450 15736
rect 16302 12960 16358 13016
rect 16486 15136 16542 15192
rect 17222 19080 17278 19136
rect 17038 18536 17094 18592
rect 16854 16088 16910 16144
rect 16670 13096 16726 13152
rect 16946 13912 17002 13968
rect 16670 12552 16726 12608
rect 16486 12280 16542 12336
rect 16302 10512 16358 10568
rect 16762 12144 16818 12200
rect 16854 11872 16910 11928
rect 17222 18536 17278 18592
rect 17130 16088 17186 16144
rect 17038 13232 17094 13288
rect 17130 12960 17186 13016
rect 17038 12708 17094 12744
rect 17038 12688 17040 12708
rect 17040 12688 17092 12708
rect 17092 12688 17094 12708
rect 17498 16632 17554 16688
rect 18602 21392 18658 21448
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18142 19352 18198 19408
rect 17774 18128 17830 18184
rect 18694 20984 18750 21040
rect 19246 22208 19302 22264
rect 19154 20576 19210 20632
rect 18142 18844 18144 18864
rect 18144 18844 18196 18864
rect 18196 18844 18198 18864
rect 18142 18808 18198 18844
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 17958 18264 18014 18320
rect 18418 18028 18420 18048
rect 18420 18028 18472 18048
rect 18472 18028 18474 18048
rect 18418 17992 18474 18028
rect 19154 19352 19210 19408
rect 18970 19216 19026 19272
rect 19338 20168 19394 20224
rect 19706 19760 19762 19816
rect 18970 18672 19026 18728
rect 18878 17856 18934 17912
rect 18510 17448 18566 17504
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18326 16904 18382 16960
rect 18418 16768 18474 16824
rect 17958 16632 18014 16688
rect 17682 16360 17738 16416
rect 17498 14864 17554 14920
rect 17406 14320 17462 14376
rect 16762 10920 16818 10976
rect 16394 9036 16450 9072
rect 16394 9016 16396 9036
rect 16396 9016 16448 9036
rect 16448 9016 16450 9036
rect 16210 8336 16266 8392
rect 16302 2644 16358 2680
rect 16302 2624 16304 2644
rect 16304 2624 16356 2644
rect 16356 2624 16358 2644
rect 16946 10104 17002 10160
rect 16946 10004 16948 10024
rect 16948 10004 17000 10024
rect 17000 10004 17002 10024
rect 16946 9968 17002 10004
rect 17406 12552 17462 12608
rect 17130 9596 17132 9616
rect 17132 9596 17184 9616
rect 17184 9596 17186 9616
rect 17130 9560 17186 9596
rect 16946 8472 17002 8528
rect 16946 8336 17002 8392
rect 16854 6840 16910 6896
rect 17038 8200 17094 8256
rect 17038 7656 17094 7712
rect 17222 6840 17278 6896
rect 16946 6568 17002 6624
rect 17682 13232 17738 13288
rect 18050 16496 18106 16552
rect 18878 17312 18934 17368
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18510 16088 18566 16144
rect 18142 15852 18144 15872
rect 18144 15852 18196 15872
rect 18196 15852 18198 15872
rect 18142 15816 18198 15852
rect 18326 15700 18382 15736
rect 18326 15680 18328 15700
rect 18328 15680 18380 15700
rect 18380 15680 18382 15700
rect 17958 15408 18014 15464
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18050 15000 18106 15056
rect 18694 14728 18750 14784
rect 18142 14456 18198 14512
rect 18326 14456 18382 14512
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18694 14320 18750 14376
rect 19246 18536 19302 18592
rect 18970 14592 19026 14648
rect 18878 13640 18934 13696
rect 18050 13504 18106 13560
rect 18510 13096 18566 13152
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 17866 12416 17922 12472
rect 17682 10784 17738 10840
rect 17590 9832 17646 9888
rect 17590 9288 17646 9344
rect 18510 12144 18566 12200
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18050 11600 18106 11656
rect 18418 11464 18474 11520
rect 17866 9832 17922 9888
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18142 10376 18198 10432
rect 18142 10124 18198 10160
rect 18142 10104 18144 10124
rect 18144 10104 18196 10124
rect 18196 10104 18198 10124
rect 18050 9968 18106 10024
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 17498 7520 17554 7576
rect 17406 6704 17462 6760
rect 17498 5208 17554 5264
rect 17406 4528 17462 4584
rect 17406 3168 17462 3224
rect 17498 2760 17554 2816
rect 18786 13232 18842 13288
rect 18694 12960 18750 13016
rect 18786 12688 18842 12744
rect 18694 12552 18750 12608
rect 18786 10648 18842 10704
rect 19154 16904 19210 16960
rect 20626 21800 20682 21856
rect 19246 16360 19302 16416
rect 19430 17040 19486 17096
rect 19246 16124 19248 16144
rect 19248 16124 19300 16144
rect 19300 16124 19302 16144
rect 19246 16088 19302 16124
rect 19338 15952 19394 16008
rect 19246 15272 19302 15328
rect 19154 13504 19210 13560
rect 19062 12552 19118 12608
rect 18602 9288 18658 9344
rect 18602 9036 18658 9072
rect 18602 9016 18604 9036
rect 18604 9016 18656 9036
rect 18656 9016 18658 9036
rect 17958 8744 18014 8800
rect 17774 6840 17830 6896
rect 17682 6432 17738 6488
rect 18510 8744 18566 8800
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18234 8064 18290 8120
rect 18694 8200 18750 8256
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18694 7656 18750 7712
rect 18602 7520 18658 7576
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18418 6316 18474 6352
rect 18418 6296 18420 6316
rect 18420 6296 18472 6316
rect 18472 6296 18474 6316
rect 17958 5652 17960 5672
rect 17960 5652 18012 5672
rect 18012 5652 18014 5672
rect 17958 5616 18014 5652
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 17958 5344 18014 5400
rect 17958 5208 18014 5264
rect 18694 7384 18750 7440
rect 18602 6840 18658 6896
rect 18694 6568 18750 6624
rect 18694 5752 18750 5808
rect 19522 14864 19578 14920
rect 19430 13776 19486 13832
rect 19338 12688 19394 12744
rect 19154 11872 19210 11928
rect 19154 11192 19210 11248
rect 19062 10104 19118 10160
rect 19430 11756 19486 11792
rect 19430 11736 19432 11756
rect 19432 11736 19484 11756
rect 19484 11736 19486 11756
rect 19430 11500 19432 11520
rect 19432 11500 19484 11520
rect 19484 11500 19486 11520
rect 19430 11464 19486 11500
rect 18970 6160 19026 6216
rect 18970 5888 19026 5944
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 17590 2488 17646 2544
rect 17038 1944 17094 2000
rect 17222 2352 17278 2408
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18878 3984 18934 4040
rect 18694 3168 18750 3224
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 3422 176 3478 232
rect 17958 448 18014 504
rect 18602 2080 18658 2136
rect 18786 2488 18842 2544
rect 18694 1264 18750 1320
rect 18970 2760 19026 2816
rect 19430 8472 19486 8528
rect 19338 8064 19394 8120
rect 19706 15544 19762 15600
rect 19614 14184 19670 14240
rect 19798 14048 19854 14104
rect 19798 12824 19854 12880
rect 19982 15544 20038 15600
rect 19982 14864 20038 14920
rect 19614 11872 19670 11928
rect 19890 12436 19946 12472
rect 19890 12416 19892 12436
rect 19892 12416 19944 12436
rect 19944 12416 19946 12436
rect 19890 12144 19946 12200
rect 19706 9324 19708 9344
rect 19708 9324 19760 9344
rect 19760 9324 19762 9344
rect 19706 9288 19762 9324
rect 19706 9016 19762 9072
rect 19338 7964 19340 7984
rect 19340 7964 19392 7984
rect 19392 7964 19394 7984
rect 19338 7928 19394 7964
rect 19246 7656 19302 7712
rect 20166 14728 20222 14784
rect 20166 14592 20222 14648
rect 20074 12960 20130 13016
rect 20166 11056 20222 11112
rect 20350 17720 20406 17776
rect 20902 17040 20958 17096
rect 20718 15680 20774 15736
rect 19706 7520 19762 7576
rect 19522 7384 19578 7440
rect 19522 7248 19578 7304
rect 19154 7112 19210 7168
rect 19154 4120 19210 4176
rect 19338 3168 19394 3224
rect 19982 7792 20038 7848
rect 19982 7248 20038 7304
rect 19982 7112 20038 7168
rect 20074 6840 20130 6896
rect 20166 6724 20222 6760
rect 20166 6704 20168 6724
rect 20168 6704 20220 6724
rect 20220 6704 20222 6724
rect 19890 5344 19946 5400
rect 19154 2760 19210 2816
rect 18970 2216 19026 2272
rect 19246 1944 19302 2000
rect 20350 9968 20406 10024
rect 20718 13368 20774 13424
rect 20994 16224 21050 16280
rect 21178 15816 21234 15872
rect 21086 13912 21142 13968
rect 20810 7384 20866 7440
rect 21086 11600 21142 11656
rect 21270 11192 21326 11248
rect 21362 8880 21418 8936
rect 21086 8608 21142 8664
rect 20994 6976 21050 7032
rect 20718 6568 20774 6624
rect 20534 6432 20590 6488
rect 20442 2932 20444 2952
rect 20444 2932 20496 2952
rect 20496 2932 20498 2952
rect 20442 2896 20498 2932
rect 20718 3712 20774 3768
rect 20718 3440 20774 3496
rect 20810 3168 20866 3224
rect 20994 2488 21050 2544
rect 21178 1672 21234 1728
rect 21914 3304 21970 3360
rect 18786 176 18842 232
<< metal3 >>
rect 0 22674 480 22704
rect 3550 22674 3556 22676
rect 0 22614 3556 22674
rect 0 22584 480 22614
rect 3550 22612 3556 22614
rect 3620 22612 3626 22676
rect 20805 22674 20871 22677
rect 22320 22674 22800 22704
rect 20805 22672 22800 22674
rect 20805 22616 20810 22672
rect 20866 22616 22800 22672
rect 20805 22614 22800 22616
rect 20805 22611 20871 22614
rect 22320 22584 22800 22614
rect 0 22266 480 22296
rect 3877 22266 3943 22269
rect 0 22264 3943 22266
rect 0 22208 3882 22264
rect 3938 22208 3943 22264
rect 0 22206 3943 22208
rect 0 22176 480 22206
rect 3877 22203 3943 22206
rect 19241 22266 19307 22269
rect 22320 22266 22800 22296
rect 19241 22264 22800 22266
rect 19241 22208 19246 22264
rect 19302 22208 22800 22264
rect 19241 22206 22800 22208
rect 19241 22203 19307 22206
rect 22320 22176 22800 22206
rect 0 21858 480 21888
rect 3693 21858 3759 21861
rect 0 21856 3759 21858
rect 0 21800 3698 21856
rect 3754 21800 3759 21856
rect 0 21798 3759 21800
rect 0 21768 480 21798
rect 3693 21795 3759 21798
rect 20621 21858 20687 21861
rect 22320 21858 22800 21888
rect 20621 21856 22800 21858
rect 20621 21800 20626 21856
rect 20682 21800 22800 21856
rect 20621 21798 22800 21800
rect 20621 21795 20687 21798
rect 22320 21768 22800 21798
rect 0 21450 480 21480
rect 4061 21450 4127 21453
rect 0 21448 4127 21450
rect 0 21392 4066 21448
rect 4122 21392 4127 21448
rect 0 21390 4127 21392
rect 0 21360 480 21390
rect 4061 21387 4127 21390
rect 18597 21450 18663 21453
rect 22320 21450 22800 21480
rect 18597 21448 22800 21450
rect 18597 21392 18602 21448
rect 18658 21392 22800 21448
rect 18597 21390 22800 21392
rect 18597 21387 18663 21390
rect 22320 21360 22800 21390
rect 0 21042 480 21072
rect 1945 21042 2011 21045
rect 0 21040 2011 21042
rect 0 20984 1950 21040
rect 2006 20984 2011 21040
rect 0 20982 2011 20984
rect 0 20952 480 20982
rect 1945 20979 2011 20982
rect 18689 21042 18755 21045
rect 22320 21042 22800 21072
rect 18689 21040 22800 21042
rect 18689 20984 18694 21040
rect 18750 20984 22800 21040
rect 18689 20982 22800 20984
rect 18689 20979 18755 20982
rect 22320 20952 22800 20982
rect 0 20634 480 20664
rect 1853 20634 1919 20637
rect 0 20632 1919 20634
rect 0 20576 1858 20632
rect 1914 20576 1919 20632
rect 0 20574 1919 20576
rect 0 20544 480 20574
rect 1853 20571 1919 20574
rect 19149 20634 19215 20637
rect 22320 20634 22800 20664
rect 19149 20632 22800 20634
rect 19149 20576 19154 20632
rect 19210 20576 22800 20632
rect 19149 20574 22800 20576
rect 19149 20571 19215 20574
rect 22320 20544 22800 20574
rect 0 20226 480 20256
rect 3877 20226 3943 20229
rect 0 20224 3943 20226
rect 0 20168 3882 20224
rect 3938 20168 3943 20224
rect 0 20166 3943 20168
rect 0 20136 480 20166
rect 3877 20163 3943 20166
rect 19333 20226 19399 20229
rect 22320 20226 22800 20256
rect 19333 20224 22800 20226
rect 19333 20168 19338 20224
rect 19394 20168 22800 20224
rect 19333 20166 22800 20168
rect 19333 20163 19399 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 2313 19954 2379 19957
rect 8753 19954 8819 19957
rect 2313 19952 8819 19954
rect 2313 19896 2318 19952
rect 2374 19896 8758 19952
rect 8814 19896 8819 19952
rect 2313 19894 8819 19896
rect 2313 19891 2379 19894
rect 0 19818 480 19848
rect 2773 19818 2839 19821
rect 0 19816 2839 19818
rect 0 19760 2778 19816
rect 2834 19760 2839 19816
rect 0 19758 2839 19760
rect 0 19728 480 19758
rect 2773 19755 2839 19758
rect 4705 19818 4771 19821
rect 6085 19818 6151 19821
rect 4705 19816 6151 19818
rect 4705 19760 4710 19816
rect 4766 19760 6090 19816
rect 6146 19760 6151 19816
rect 4705 19758 6151 19760
rect 4705 19755 4771 19758
rect 6085 19755 6151 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 0 19410 480 19440
rect 8342 19413 8402 19894
rect 8753 19891 8819 19894
rect 19701 19818 19767 19821
rect 22320 19818 22800 19848
rect 19701 19816 22800 19818
rect 19701 19760 19706 19816
rect 19762 19760 22800 19816
rect 19701 19758 22800 19760
rect 19701 19755 19767 19758
rect 22320 19728 22800 19758
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 15929 19546 15995 19549
rect 16481 19546 16547 19549
rect 15929 19544 16547 19546
rect 15929 19488 15934 19544
rect 15990 19488 16486 19544
rect 16542 19488 16547 19544
rect 15929 19486 16547 19488
rect 15929 19483 15995 19486
rect 16481 19483 16547 19486
rect 1945 19410 2011 19413
rect 0 19408 2011 19410
rect 0 19352 1950 19408
rect 2006 19352 2011 19408
rect 0 19350 2011 19352
rect 0 19320 480 19350
rect 1945 19347 2011 19350
rect 4061 19410 4127 19413
rect 5533 19410 5599 19413
rect 4061 19408 5599 19410
rect 4061 19352 4066 19408
rect 4122 19352 5538 19408
rect 5594 19352 5599 19408
rect 4061 19350 5599 19352
rect 8342 19408 8451 19413
rect 8342 19352 8390 19408
rect 8446 19352 8451 19408
rect 8342 19350 8451 19352
rect 4061 19347 4127 19350
rect 5533 19347 5599 19350
rect 8385 19347 8451 19350
rect 14917 19410 14983 19413
rect 18137 19410 18203 19413
rect 14917 19408 18203 19410
rect 14917 19352 14922 19408
rect 14978 19352 18142 19408
rect 18198 19352 18203 19408
rect 14917 19350 18203 19352
rect 14917 19347 14983 19350
rect 18137 19347 18203 19350
rect 19149 19410 19215 19413
rect 22320 19410 22800 19440
rect 19149 19408 22800 19410
rect 19149 19352 19154 19408
rect 19210 19352 22800 19408
rect 19149 19350 22800 19352
rect 19149 19347 19215 19350
rect 22320 19320 22800 19350
rect 4429 19274 4495 19277
rect 11830 19274 11836 19276
rect 4429 19272 11836 19274
rect 4429 19216 4434 19272
rect 4490 19216 11836 19272
rect 4429 19214 11836 19216
rect 4429 19211 4495 19214
rect 11830 19212 11836 19214
rect 11900 19212 11906 19276
rect 12014 19212 12020 19276
rect 12084 19274 12090 19276
rect 18965 19274 19031 19277
rect 12084 19272 19031 19274
rect 12084 19216 18970 19272
rect 19026 19216 19031 19272
rect 12084 19214 19031 19216
rect 12084 19212 12090 19214
rect 18965 19211 19031 19214
rect 0 19138 480 19168
rect 4337 19138 4403 19141
rect 4838 19138 4844 19140
rect 0 19078 2146 19138
rect 0 19048 480 19078
rect 0 18730 480 18760
rect 1945 18730 2011 18733
rect 0 18728 2011 18730
rect 0 18672 1950 18728
rect 2006 18672 2011 18728
rect 0 18670 2011 18672
rect 2086 18730 2146 19078
rect 4337 19136 4844 19138
rect 4337 19080 4342 19136
rect 4398 19080 4844 19136
rect 4337 19078 4844 19080
rect 4337 19075 4403 19078
rect 4838 19076 4844 19078
rect 4908 19076 4914 19140
rect 8569 19138 8635 19141
rect 9806 19138 9812 19140
rect 8569 19136 9812 19138
rect 8569 19080 8574 19136
rect 8630 19080 9812 19136
rect 8569 19078 9812 19080
rect 8569 19075 8635 19078
rect 9806 19076 9812 19078
rect 9876 19138 9882 19140
rect 12249 19138 12315 19141
rect 9876 19136 12315 19138
rect 9876 19080 12254 19136
rect 12310 19080 12315 19136
rect 9876 19078 12315 19080
rect 9876 19076 9882 19078
rect 12249 19075 12315 19078
rect 17217 19138 17283 19141
rect 17718 19138 17724 19140
rect 17217 19136 17724 19138
rect 17217 19080 17222 19136
rect 17278 19080 17724 19136
rect 17217 19078 17724 19080
rect 17217 19075 17283 19078
rect 17718 19076 17724 19078
rect 17788 19138 17794 19140
rect 22320 19138 22800 19168
rect 17788 19078 22800 19138
rect 17788 19076 17794 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 22320 19048 22800 19078
rect 14672 19007 14992 19008
rect 5165 19002 5231 19005
rect 5390 19002 5396 19004
rect 5165 19000 5396 19002
rect 5165 18944 5170 19000
rect 5226 18944 5396 19000
rect 5165 18942 5396 18944
rect 5165 18939 5231 18942
rect 5390 18940 5396 18942
rect 5460 18940 5466 19004
rect 7373 19002 7439 19005
rect 7557 19002 7623 19005
rect 7373 19000 7623 19002
rect 7373 18944 7378 19000
rect 7434 18944 7562 19000
rect 7618 18944 7623 19000
rect 7373 18942 7623 18944
rect 7373 18939 7439 18942
rect 7557 18939 7623 18942
rect 10041 19002 10107 19005
rect 13261 19002 13327 19005
rect 10041 19000 13327 19002
rect 10041 18944 10046 19000
rect 10102 18944 13266 19000
rect 13322 18944 13327 19000
rect 10041 18942 13327 18944
rect 10041 18939 10107 18942
rect 13261 18939 13327 18942
rect 13905 19002 13971 19005
rect 14038 19002 14044 19004
rect 13905 19000 14044 19002
rect 13905 18944 13910 19000
rect 13966 18944 14044 19000
rect 13905 18942 14044 18944
rect 13905 18939 13971 18942
rect 14038 18940 14044 18942
rect 14108 18940 14114 19004
rect 3877 18866 3943 18869
rect 18137 18866 18203 18869
rect 3877 18864 18203 18866
rect 3877 18808 3882 18864
rect 3938 18808 18142 18864
rect 18198 18808 18203 18864
rect 3877 18806 18203 18808
rect 3877 18803 3943 18806
rect 18137 18803 18203 18806
rect 18965 18730 19031 18733
rect 22320 18730 22800 18760
rect 2086 18670 18568 18730
rect 0 18640 480 18670
rect 1945 18667 2011 18670
rect 4838 18532 4844 18596
rect 4908 18594 4914 18596
rect 6453 18594 6519 18597
rect 4908 18592 6519 18594
rect 4908 18536 6458 18592
rect 6514 18536 6519 18592
rect 4908 18534 6519 18536
rect 4908 18532 4914 18534
rect 6453 18531 6519 18534
rect 13445 18594 13511 18597
rect 17033 18594 17099 18597
rect 17217 18594 17283 18597
rect 13445 18592 17283 18594
rect 13445 18536 13450 18592
rect 13506 18536 17038 18592
rect 17094 18536 17222 18592
rect 17278 18536 17283 18592
rect 13445 18534 17283 18536
rect 18508 18594 18568 18670
rect 18965 18728 22800 18730
rect 18965 18672 18970 18728
rect 19026 18672 22800 18728
rect 18965 18670 22800 18672
rect 18965 18667 19031 18670
rect 22320 18640 22800 18670
rect 19241 18594 19307 18597
rect 18508 18592 19307 18594
rect 18508 18536 19246 18592
rect 19302 18536 19307 18592
rect 18508 18534 19307 18536
rect 13445 18531 13511 18534
rect 17033 18531 17099 18534
rect 17217 18531 17283 18534
rect 19241 18531 19307 18534
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 7189 18458 7255 18461
rect 8385 18458 8451 18461
rect 10174 18458 10180 18460
rect 7189 18456 8451 18458
rect 7189 18400 7194 18456
rect 7250 18400 8390 18456
rect 8446 18400 8451 18456
rect 7189 18398 8451 18400
rect 7189 18395 7255 18398
rect 8385 18395 8451 18398
rect 8526 18398 10180 18458
rect 0 18322 480 18352
rect 3233 18322 3299 18325
rect 3918 18322 3924 18324
rect 0 18262 1410 18322
rect 0 18232 480 18262
rect 1350 18186 1410 18262
rect 3233 18320 3924 18322
rect 3233 18264 3238 18320
rect 3294 18264 3924 18320
rect 3233 18262 3924 18264
rect 3233 18259 3299 18262
rect 3918 18260 3924 18262
rect 3988 18260 3994 18324
rect 4429 18322 4495 18325
rect 8526 18322 8586 18398
rect 10174 18396 10180 18398
rect 10244 18396 10250 18460
rect 12750 18396 12756 18460
rect 12820 18458 12826 18460
rect 15837 18458 15903 18461
rect 12820 18456 15903 18458
rect 12820 18400 15842 18456
rect 15898 18400 15903 18456
rect 12820 18398 15903 18400
rect 12820 18396 12826 18398
rect 15837 18395 15903 18398
rect 4429 18320 8586 18322
rect 4429 18264 4434 18320
rect 4490 18264 8586 18320
rect 4429 18262 8586 18264
rect 8661 18322 8727 18325
rect 9438 18322 9444 18324
rect 8661 18320 9444 18322
rect 8661 18264 8666 18320
rect 8722 18264 9444 18320
rect 8661 18262 9444 18264
rect 4429 18259 4495 18262
rect 8661 18259 8727 18262
rect 9438 18260 9444 18262
rect 9508 18322 9514 18324
rect 13721 18322 13787 18325
rect 9508 18320 13787 18322
rect 9508 18264 13726 18320
rect 13782 18264 13787 18320
rect 9508 18262 13787 18264
rect 9508 18260 9514 18262
rect 13721 18259 13787 18262
rect 15142 18260 15148 18324
rect 15212 18322 15218 18324
rect 16297 18322 16363 18325
rect 15212 18320 16363 18322
rect 15212 18264 16302 18320
rect 16358 18264 16363 18320
rect 15212 18262 16363 18264
rect 15212 18260 15218 18262
rect 16297 18259 16363 18262
rect 17953 18322 18019 18325
rect 22320 18322 22800 18352
rect 17953 18320 22800 18322
rect 17953 18264 17958 18320
rect 18014 18264 22800 18320
rect 17953 18262 22800 18264
rect 17953 18259 18019 18262
rect 22320 18232 22800 18262
rect 3141 18186 3207 18189
rect 1350 18184 3207 18186
rect 1350 18128 3146 18184
rect 3202 18128 3207 18184
rect 1350 18126 3207 18128
rect 3141 18123 3207 18126
rect 3325 18186 3391 18189
rect 9765 18186 9831 18189
rect 3325 18184 9831 18186
rect 3325 18128 3330 18184
rect 3386 18128 9770 18184
rect 9826 18128 9831 18184
rect 3325 18126 9831 18128
rect 3325 18123 3391 18126
rect 9765 18123 9831 18126
rect 10685 18186 10751 18189
rect 11646 18186 11652 18188
rect 10685 18184 11652 18186
rect 10685 18128 10690 18184
rect 10746 18128 11652 18184
rect 10685 18126 11652 18128
rect 10685 18123 10751 18126
rect 11646 18124 11652 18126
rect 11716 18124 11722 18188
rect 14365 18186 14431 18189
rect 14549 18186 14615 18189
rect 17769 18186 17835 18189
rect 14365 18184 14474 18186
rect 14365 18128 14370 18184
rect 14426 18128 14474 18184
rect 14365 18123 14474 18128
rect 14549 18184 17835 18186
rect 14549 18128 14554 18184
rect 14610 18128 17774 18184
rect 17830 18128 17835 18184
rect 14549 18126 17835 18128
rect 14549 18123 14615 18126
rect 17769 18123 17835 18126
rect 1669 18050 1735 18053
rect 3601 18050 3667 18053
rect 3734 18050 3740 18052
rect 1669 18048 3434 18050
rect 1669 17992 1674 18048
rect 1730 17992 3434 18048
rect 1669 17990 3434 17992
rect 1669 17987 1735 17990
rect 0 17914 480 17944
rect 1485 17914 1551 17917
rect 0 17912 1551 17914
rect 0 17856 1490 17912
rect 1546 17856 1551 17912
rect 0 17854 1551 17856
rect 3374 17914 3434 17990
rect 3601 18048 3740 18050
rect 3601 17992 3606 18048
rect 3662 17992 3740 18048
rect 3601 17990 3740 17992
rect 3601 17987 3667 17990
rect 3734 17988 3740 17990
rect 3804 17988 3810 18052
rect 7189 18050 7255 18053
rect 3926 18048 7255 18050
rect 3926 17992 7194 18048
rect 7250 17992 7255 18048
rect 3926 17990 7255 17992
rect 3926 17914 3986 17990
rect 7189 17987 7255 17990
rect 8385 18050 8451 18053
rect 9029 18050 9095 18053
rect 12525 18050 12591 18053
rect 8385 18048 12591 18050
rect 8385 17992 8390 18048
rect 8446 17992 9034 18048
rect 9090 17992 12530 18048
rect 12586 17992 12591 18048
rect 8385 17990 12591 17992
rect 8385 17987 8451 17990
rect 9029 17987 9095 17990
rect 12525 17987 12591 17990
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 3374 17854 3986 17914
rect 14273 17914 14339 17917
rect 14414 17914 14474 18123
rect 18413 18050 18479 18053
rect 18638 18050 18644 18052
rect 18413 18048 18644 18050
rect 18413 17992 18418 18048
rect 18474 17992 18644 18048
rect 18413 17990 18644 17992
rect 18413 17987 18479 17990
rect 18638 17988 18644 17990
rect 18708 17988 18714 18052
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 14273 17912 14474 17914
rect 14273 17856 14278 17912
rect 14334 17856 14474 17912
rect 14273 17854 14474 17856
rect 18873 17914 18939 17917
rect 22320 17914 22800 17944
rect 18873 17912 22800 17914
rect 18873 17856 18878 17912
rect 18934 17856 22800 17912
rect 18873 17854 22800 17856
rect 0 17824 480 17854
rect 1485 17851 1551 17854
rect 14273 17851 14339 17854
rect 18873 17851 18939 17854
rect 22320 17824 22800 17854
rect 1853 17778 1919 17781
rect 5257 17778 5323 17781
rect 1853 17776 5323 17778
rect 1853 17720 1858 17776
rect 1914 17720 5262 17776
rect 5318 17720 5323 17776
rect 1853 17718 5323 17720
rect 1853 17715 1919 17718
rect 5257 17715 5323 17718
rect 13537 17778 13603 17781
rect 20345 17778 20411 17781
rect 13537 17776 20411 17778
rect 13537 17720 13542 17776
rect 13598 17720 20350 17776
rect 20406 17720 20411 17776
rect 13537 17718 20411 17720
rect 13537 17715 13603 17718
rect 20345 17715 20411 17718
rect 1761 17642 1827 17645
rect 6085 17642 6151 17645
rect 1761 17640 6151 17642
rect 1761 17584 1766 17640
rect 1822 17584 6090 17640
rect 6146 17584 6151 17640
rect 1761 17582 6151 17584
rect 1761 17579 1827 17582
rect 6085 17579 6151 17582
rect 14641 17642 14707 17645
rect 15285 17644 15351 17645
rect 15285 17642 15332 17644
rect 14641 17640 15332 17642
rect 14641 17584 14646 17640
rect 14702 17584 15290 17640
rect 14641 17582 15332 17584
rect 14641 17579 14707 17582
rect 15285 17580 15332 17582
rect 15396 17580 15402 17644
rect 15285 17579 15351 17580
rect 0 17506 480 17536
rect 2773 17506 2839 17509
rect 0 17504 2839 17506
rect 0 17448 2778 17504
rect 2834 17448 2839 17504
rect 0 17446 2839 17448
rect 0 17416 480 17446
rect 2773 17443 2839 17446
rect 14406 17444 14412 17508
rect 14476 17506 14482 17508
rect 16021 17506 16087 17509
rect 14476 17504 16087 17506
rect 14476 17448 16026 17504
rect 16082 17448 16087 17504
rect 14476 17446 16087 17448
rect 14476 17444 14482 17446
rect 16021 17443 16087 17446
rect 18505 17506 18571 17509
rect 22320 17506 22800 17536
rect 18505 17504 22800 17506
rect 18505 17448 18510 17504
rect 18566 17448 22800 17504
rect 18505 17446 22800 17448
rect 18505 17443 18571 17446
rect 4376 17440 4696 17441
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 22320 17416 22800 17446
rect 18104 17375 18424 17376
rect 18873 17370 18939 17373
rect 19006 17370 19012 17372
rect 18873 17368 19012 17370
rect 18873 17312 18878 17368
rect 18934 17312 19012 17368
rect 18873 17310 19012 17312
rect 18873 17307 18939 17310
rect 19006 17308 19012 17310
rect 19076 17308 19082 17372
rect 3417 17234 3483 17237
rect 7414 17234 7420 17236
rect 3417 17232 7420 17234
rect 3417 17176 3422 17232
rect 3478 17176 7420 17232
rect 3417 17174 7420 17176
rect 3417 17171 3483 17174
rect 7414 17172 7420 17174
rect 7484 17234 7490 17236
rect 8017 17234 8083 17237
rect 7484 17232 8083 17234
rect 7484 17176 8022 17232
rect 8078 17176 8083 17232
rect 7484 17174 8083 17176
rect 7484 17172 7490 17174
rect 8017 17171 8083 17174
rect 10542 17172 10548 17236
rect 10612 17234 10618 17236
rect 16389 17234 16455 17237
rect 10612 17232 16455 17234
rect 10612 17176 16394 17232
rect 16450 17176 16455 17232
rect 10612 17174 16455 17176
rect 10612 17172 10618 17174
rect 16389 17171 16455 17174
rect 0 17098 480 17128
rect 1577 17098 1643 17101
rect 0 17096 1643 17098
rect 0 17040 1582 17096
rect 1638 17040 1643 17096
rect 0 17038 1643 17040
rect 0 17008 480 17038
rect 1577 17035 1643 17038
rect 2773 17098 2839 17101
rect 6085 17098 6151 17101
rect 11789 17098 11855 17101
rect 2773 17096 11855 17098
rect 2773 17040 2778 17096
rect 2834 17040 6090 17096
rect 6146 17040 11794 17096
rect 11850 17040 11855 17096
rect 2773 17038 11855 17040
rect 2773 17035 2839 17038
rect 6085 17035 6151 17038
rect 11789 17035 11855 17038
rect 12709 17098 12775 17101
rect 12934 17098 12940 17100
rect 12709 17096 12940 17098
rect 12709 17040 12714 17096
rect 12770 17040 12940 17096
rect 12709 17038 12940 17040
rect 12709 17035 12775 17038
rect 12934 17036 12940 17038
rect 13004 17098 13010 17100
rect 16573 17098 16639 17101
rect 13004 17096 16639 17098
rect 13004 17040 16578 17096
rect 16634 17040 16639 17096
rect 13004 17038 16639 17040
rect 13004 17036 13010 17038
rect 16573 17035 16639 17038
rect 18822 17036 18828 17100
rect 18892 17098 18898 17100
rect 19425 17098 19491 17101
rect 18892 17096 19491 17098
rect 18892 17040 19430 17096
rect 19486 17040 19491 17096
rect 18892 17038 19491 17040
rect 18892 17036 18898 17038
rect 19425 17035 19491 17038
rect 20897 17098 20963 17101
rect 22320 17098 22800 17128
rect 20897 17096 22800 17098
rect 20897 17040 20902 17096
rect 20958 17040 22800 17096
rect 20897 17038 22800 17040
rect 20897 17035 20963 17038
rect 22320 17008 22800 17038
rect 3969 16962 4035 16965
rect 4838 16962 4844 16964
rect 3969 16960 4844 16962
rect 3969 16904 3974 16960
rect 4030 16904 4844 16960
rect 3969 16902 4844 16904
rect 3969 16899 4035 16902
rect 4838 16900 4844 16902
rect 4908 16900 4914 16964
rect 10961 16962 11027 16965
rect 13077 16962 13143 16965
rect 10961 16960 13143 16962
rect 10961 16904 10966 16960
rect 11022 16904 13082 16960
rect 13138 16904 13143 16960
rect 10961 16902 13143 16904
rect 10961 16899 11027 16902
rect 13077 16899 13143 16902
rect 14222 16900 14228 16964
rect 14292 16962 14298 16964
rect 14365 16962 14431 16965
rect 14292 16960 14431 16962
rect 14292 16904 14370 16960
rect 14426 16904 14431 16960
rect 14292 16902 14431 16904
rect 14292 16900 14298 16902
rect 14365 16899 14431 16902
rect 18321 16962 18387 16965
rect 19149 16962 19215 16965
rect 18321 16960 19215 16962
rect 18321 16904 18326 16960
rect 18382 16904 19154 16960
rect 19210 16904 19215 16960
rect 18321 16902 19215 16904
rect 18321 16899 18387 16902
rect 19149 16899 19215 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 9990 16764 9996 16828
rect 10060 16826 10066 16828
rect 12065 16826 12131 16829
rect 13353 16826 13419 16829
rect 10060 16824 13419 16826
rect 10060 16768 12070 16824
rect 12126 16768 13358 16824
rect 13414 16768 13419 16824
rect 10060 16766 13419 16768
rect 10060 16764 10066 16766
rect 12065 16763 12131 16766
rect 13353 16763 13419 16766
rect 17902 16764 17908 16828
rect 17972 16826 17978 16828
rect 18413 16826 18479 16829
rect 17972 16824 18479 16826
rect 17972 16768 18418 16824
rect 18474 16768 18479 16824
rect 17972 16766 18479 16768
rect 17972 16764 17978 16766
rect 18413 16763 18479 16766
rect 0 16690 480 16720
rect 4337 16690 4403 16693
rect 0 16688 4403 16690
rect 0 16632 4342 16688
rect 4398 16632 4403 16688
rect 0 16630 4403 16632
rect 0 16600 480 16630
rect 4337 16627 4403 16630
rect 6545 16690 6611 16693
rect 8937 16690 9003 16693
rect 6545 16688 9003 16690
rect 6545 16632 6550 16688
rect 6606 16632 8942 16688
rect 8998 16632 9003 16688
rect 6545 16630 9003 16632
rect 6545 16627 6611 16630
rect 8937 16627 9003 16630
rect 14365 16690 14431 16693
rect 17493 16690 17559 16693
rect 14365 16688 17559 16690
rect 14365 16632 14370 16688
rect 14426 16632 17498 16688
rect 17554 16632 17559 16688
rect 14365 16630 17559 16632
rect 14365 16627 14431 16630
rect 17493 16627 17559 16630
rect 17953 16690 18019 16693
rect 22320 16690 22800 16720
rect 17953 16688 22800 16690
rect 17953 16632 17958 16688
rect 18014 16632 22800 16688
rect 17953 16630 22800 16632
rect 17953 16627 18019 16630
rect 22320 16600 22800 16630
rect 10174 16492 10180 16556
rect 10244 16554 10250 16556
rect 15745 16554 15811 16557
rect 10244 16552 15811 16554
rect 10244 16496 15750 16552
rect 15806 16496 15811 16552
rect 10244 16494 15811 16496
rect 10244 16492 10250 16494
rect 15745 16491 15811 16494
rect 17350 16492 17356 16556
rect 17420 16554 17426 16556
rect 18045 16554 18111 16557
rect 17420 16552 18111 16554
rect 17420 16496 18050 16552
rect 18106 16496 18111 16552
rect 17420 16494 18111 16496
rect 17420 16492 17426 16494
rect 18045 16491 18111 16494
rect 16297 16418 16363 16421
rect 17677 16418 17743 16421
rect 16297 16416 17743 16418
rect 16297 16360 16302 16416
rect 16358 16360 17682 16416
rect 17738 16360 17743 16416
rect 16297 16358 17743 16360
rect 16297 16355 16363 16358
rect 17677 16355 17743 16358
rect 19241 16418 19307 16421
rect 19558 16418 19564 16420
rect 19241 16416 19564 16418
rect 19241 16360 19246 16416
rect 19302 16360 19564 16416
rect 19241 16358 19564 16360
rect 19241 16355 19307 16358
rect 19558 16356 19564 16358
rect 19628 16356 19634 16420
rect 4376 16352 4696 16353
rect 0 16282 480 16312
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 2773 16282 2839 16285
rect 0 16280 2839 16282
rect 0 16224 2778 16280
rect 2834 16224 2839 16280
rect 0 16222 2839 16224
rect 0 16192 480 16222
rect 2773 16219 2839 16222
rect 5206 16220 5212 16284
rect 5276 16220 5282 16284
rect 11830 16220 11836 16284
rect 11900 16282 11906 16284
rect 13537 16282 13603 16285
rect 11900 16280 13603 16282
rect 11900 16224 13542 16280
rect 13598 16224 13603 16280
rect 11900 16222 13603 16224
rect 11900 16220 11906 16222
rect 2405 16146 2471 16149
rect 5214 16146 5274 16220
rect 13537 16219 13603 16222
rect 20989 16282 21055 16285
rect 22320 16282 22800 16312
rect 20989 16280 22800 16282
rect 20989 16224 20994 16280
rect 21050 16224 22800 16280
rect 20989 16222 22800 16224
rect 20989 16219 21055 16222
rect 22320 16192 22800 16222
rect 11973 16146 12039 16149
rect 2405 16144 12039 16146
rect 2405 16088 2410 16144
rect 2466 16088 11978 16144
rect 12034 16088 12039 16144
rect 2405 16086 12039 16088
rect 2405 16083 2471 16086
rect 11973 16083 12039 16086
rect 16430 16084 16436 16148
rect 16500 16146 16506 16148
rect 16849 16146 16915 16149
rect 16500 16144 16915 16146
rect 16500 16088 16854 16144
rect 16910 16088 16915 16144
rect 16500 16086 16915 16088
rect 16500 16084 16506 16086
rect 16849 16083 16915 16086
rect 17125 16146 17191 16149
rect 18505 16146 18571 16149
rect 19241 16146 19307 16149
rect 17125 16144 18571 16146
rect 17125 16088 17130 16144
rect 17186 16088 18510 16144
rect 18566 16088 18571 16144
rect 17125 16086 18571 16088
rect 17125 16083 17191 16086
rect 18505 16083 18571 16086
rect 18646 16144 19307 16146
rect 18646 16088 19246 16144
rect 19302 16088 19307 16144
rect 18646 16086 19307 16088
rect 3509 16010 3575 16013
rect 5257 16010 5323 16013
rect 8845 16010 8911 16013
rect 3509 16008 8911 16010
rect 3509 15952 3514 16008
rect 3570 15952 5262 16008
rect 5318 15952 8850 16008
rect 8906 15952 8911 16008
rect 3509 15950 8911 15952
rect 3509 15947 3575 15950
rect 5257 15947 5323 15950
rect 8845 15947 8911 15950
rect 14181 16010 14247 16013
rect 18646 16010 18706 16086
rect 19241 16083 19307 16086
rect 19333 16012 19399 16013
rect 19333 16010 19380 16012
rect 14181 16008 18706 16010
rect 14181 15952 14186 16008
rect 14242 15952 18706 16008
rect 14181 15950 18706 15952
rect 19288 16008 19380 16010
rect 19288 15952 19338 16008
rect 19288 15950 19380 15952
rect 14181 15947 14247 15950
rect 19333 15948 19380 15950
rect 19444 15948 19450 16012
rect 19333 15947 19399 15948
rect 0 15874 480 15904
rect 4061 15874 4127 15877
rect 16205 15876 16271 15877
rect 16205 15874 16252 15876
rect 0 15872 4127 15874
rect 0 15816 4066 15872
rect 4122 15816 4127 15872
rect 0 15814 4127 15816
rect 16160 15872 16252 15874
rect 16160 15816 16210 15872
rect 16160 15814 16252 15816
rect 0 15784 480 15814
rect 4061 15811 4127 15814
rect 16205 15812 16252 15814
rect 16316 15812 16322 15876
rect 16481 15874 16547 15877
rect 18137 15874 18203 15877
rect 16481 15872 18203 15874
rect 16481 15816 16486 15872
rect 16542 15816 18142 15872
rect 18198 15816 18203 15872
rect 16481 15814 18203 15816
rect 16205 15811 16271 15812
rect 16481 15811 16547 15814
rect 18137 15811 18203 15814
rect 21173 15874 21239 15877
rect 22320 15874 22800 15904
rect 21173 15872 22800 15874
rect 21173 15816 21178 15872
rect 21234 15816 22800 15872
rect 21173 15814 22800 15816
rect 21173 15811 21239 15814
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 22320 15784 22800 15814
rect 14672 15743 14992 15744
rect 3233 15738 3299 15741
rect 3366 15738 3372 15740
rect 3233 15736 3372 15738
rect 3233 15680 3238 15736
rect 3294 15680 3372 15736
rect 3233 15678 3372 15680
rect 3233 15675 3299 15678
rect 3366 15676 3372 15678
rect 3436 15676 3442 15740
rect 7557 15738 7623 15741
rect 10409 15740 10475 15741
rect 10358 15738 10364 15740
rect 7422 15736 7623 15738
rect 7422 15680 7562 15736
rect 7618 15680 7623 15736
rect 7422 15678 7623 15680
rect 10318 15678 10364 15738
rect 10428 15736 10475 15740
rect 10470 15680 10475 15736
rect 2589 15602 2655 15605
rect 5625 15602 5691 15605
rect 2589 15600 5691 15602
rect 2589 15544 2594 15600
rect 2650 15544 5630 15600
rect 5686 15544 5691 15600
rect 2589 15542 5691 15544
rect 2589 15539 2655 15542
rect 5625 15539 5691 15542
rect 7281 15602 7347 15605
rect 7422 15602 7482 15678
rect 7557 15675 7623 15678
rect 10358 15676 10364 15678
rect 10428 15676 10475 15680
rect 10409 15675 10475 15676
rect 16389 15738 16455 15741
rect 18321 15738 18387 15741
rect 20713 15738 20779 15741
rect 16389 15736 18387 15738
rect 16389 15680 16394 15736
rect 16450 15680 18326 15736
rect 18382 15680 18387 15736
rect 16389 15678 18387 15680
rect 16389 15675 16455 15678
rect 18321 15675 18387 15678
rect 18600 15736 20779 15738
rect 18600 15680 20718 15736
rect 20774 15680 20779 15736
rect 18600 15678 20779 15680
rect 7281 15600 7482 15602
rect 7281 15544 7286 15600
rect 7342 15544 7482 15600
rect 7281 15542 7482 15544
rect 8477 15602 8543 15605
rect 8702 15602 8708 15604
rect 8477 15600 8708 15602
rect 8477 15544 8482 15600
rect 8538 15544 8708 15600
rect 8477 15542 8708 15544
rect 7281 15539 7347 15542
rect 8477 15539 8543 15542
rect 8702 15540 8708 15542
rect 8772 15540 8778 15604
rect 9857 15602 9923 15605
rect 18600 15602 18660 15678
rect 20713 15675 20779 15678
rect 9857 15600 18660 15602
rect 9857 15544 9862 15600
rect 9918 15544 18660 15600
rect 9857 15542 18660 15544
rect 19701 15602 19767 15605
rect 19977 15602 20043 15605
rect 19701 15600 20043 15602
rect 19701 15544 19706 15600
rect 19762 15544 19982 15600
rect 20038 15544 20043 15600
rect 19701 15542 20043 15544
rect 9857 15539 9923 15542
rect 19701 15539 19767 15542
rect 19977 15539 20043 15542
rect 0 15466 480 15496
rect 3969 15466 4035 15469
rect 0 15464 4035 15466
rect 0 15408 3974 15464
rect 4030 15408 4035 15464
rect 0 15406 4035 15408
rect 0 15376 480 15406
rect 3969 15403 4035 15406
rect 6637 15466 6703 15469
rect 7649 15466 7715 15469
rect 6637 15464 7715 15466
rect 6637 15408 6642 15464
rect 6698 15408 7654 15464
rect 7710 15408 7715 15464
rect 6637 15406 7715 15408
rect 6637 15403 6703 15406
rect 7649 15403 7715 15406
rect 10593 15466 10659 15469
rect 16246 15466 16252 15468
rect 10593 15464 16252 15466
rect 10593 15408 10598 15464
rect 10654 15408 16252 15464
rect 10593 15406 16252 15408
rect 10593 15403 10659 15406
rect 16246 15404 16252 15406
rect 16316 15404 16322 15468
rect 17953 15466 18019 15469
rect 22320 15466 22800 15496
rect 17953 15464 22800 15466
rect 17953 15408 17958 15464
rect 18014 15408 22800 15464
rect 17953 15406 22800 15408
rect 17953 15403 18019 15406
rect 22320 15376 22800 15406
rect 6729 15330 6795 15333
rect 8886 15330 8892 15332
rect 6729 15328 8892 15330
rect 6729 15272 6734 15328
rect 6790 15272 8892 15328
rect 6729 15270 8892 15272
rect 6729 15267 6795 15270
rect 8886 15268 8892 15270
rect 8956 15268 8962 15332
rect 12566 15268 12572 15332
rect 12636 15330 12642 15332
rect 15377 15330 15443 15333
rect 12636 15328 15443 15330
rect 12636 15272 15382 15328
rect 15438 15272 15443 15328
rect 12636 15270 15443 15272
rect 12636 15268 12642 15270
rect 15377 15267 15443 15270
rect 19006 15268 19012 15332
rect 19076 15330 19082 15332
rect 19241 15330 19307 15333
rect 19076 15328 19307 15330
rect 19076 15272 19246 15328
rect 19302 15272 19307 15328
rect 19076 15270 19307 15272
rect 19076 15268 19082 15270
rect 19241 15267 19307 15270
rect 4376 15264 4696 15265
rect 0 15194 480 15224
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 4061 15194 4127 15197
rect 0 15192 4127 15194
rect 0 15136 4066 15192
rect 4122 15136 4127 15192
rect 0 15134 4127 15136
rect 0 15104 480 15134
rect 4061 15131 4127 15134
rect 7465 15194 7531 15197
rect 9581 15194 9647 15197
rect 10910 15194 10916 15196
rect 7465 15192 10916 15194
rect 7465 15136 7470 15192
rect 7526 15136 9586 15192
rect 9642 15136 10916 15192
rect 7465 15134 10916 15136
rect 7465 15131 7531 15134
rect 9581 15131 9647 15134
rect 10910 15132 10916 15134
rect 10980 15132 10986 15196
rect 13486 15132 13492 15196
rect 13556 15194 13562 15196
rect 16481 15194 16547 15197
rect 22320 15194 22800 15224
rect 13556 15192 16547 15194
rect 13556 15136 16486 15192
rect 16542 15136 16547 15192
rect 13556 15134 16547 15136
rect 13556 15132 13562 15134
rect 16481 15131 16547 15134
rect 18876 15134 22800 15194
rect 6453 15058 6519 15061
rect 8109 15058 8175 15061
rect 6453 15056 8175 15058
rect 6453 15000 6458 15056
rect 6514 15000 8114 15056
rect 8170 15000 8175 15056
rect 6453 14998 8175 15000
rect 6453 14995 6519 14998
rect 8109 14995 8175 14998
rect 8293 15058 8359 15061
rect 9121 15058 9187 15061
rect 14365 15058 14431 15061
rect 18045 15058 18111 15061
rect 8293 15056 9187 15058
rect 8293 15000 8298 15056
rect 8354 15000 9126 15056
rect 9182 15000 9187 15056
rect 8293 14998 9187 15000
rect 8293 14995 8359 14998
rect 9121 14995 9187 14998
rect 12712 14998 14290 15058
rect 12712 14925 12772 14998
rect 3325 14922 3391 14925
rect 12709 14922 12775 14925
rect 3325 14920 12775 14922
rect 3325 14864 3330 14920
rect 3386 14864 12714 14920
rect 12770 14864 12775 14920
rect 3325 14862 12775 14864
rect 14230 14922 14290 14998
rect 14365 15056 18111 15058
rect 14365 15000 14370 15056
rect 14426 15000 18050 15056
rect 18106 15000 18111 15056
rect 14365 14998 18111 15000
rect 14365 14995 14431 14998
rect 18045 14995 18111 14998
rect 17493 14922 17559 14925
rect 18876 14922 18936 15134
rect 22320 15104 22800 15134
rect 14230 14862 17418 14922
rect 3325 14859 3391 14862
rect 12709 14859 12775 14862
rect 0 14786 480 14816
rect 3785 14786 3851 14789
rect 0 14784 3851 14786
rect 0 14728 3790 14784
rect 3846 14728 3851 14784
rect 0 14726 3851 14728
rect 17358 14786 17418 14862
rect 17493 14920 18936 14922
rect 17493 14864 17498 14920
rect 17554 14864 18936 14920
rect 17493 14862 18936 14864
rect 17493 14859 17559 14862
rect 19006 14860 19012 14924
rect 19076 14922 19082 14924
rect 19517 14922 19583 14925
rect 19977 14922 20043 14925
rect 19076 14920 19583 14922
rect 19076 14864 19522 14920
rect 19578 14864 19583 14920
rect 19076 14862 19583 14864
rect 19076 14860 19082 14862
rect 19517 14859 19583 14862
rect 19934 14920 20043 14922
rect 19934 14864 19982 14920
rect 20038 14864 20043 14920
rect 19934 14859 20043 14864
rect 18689 14786 18755 14789
rect 18822 14786 18828 14788
rect 17358 14784 18828 14786
rect 17358 14728 18694 14784
rect 18750 14728 18828 14784
rect 17358 14726 18828 14728
rect 0 14696 480 14726
rect 3785 14723 3851 14726
rect 18689 14723 18755 14726
rect 18822 14724 18828 14726
rect 18892 14724 18898 14788
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 5441 14650 5507 14653
rect 6085 14650 6151 14653
rect 5441 14648 6151 14650
rect 5441 14592 5446 14648
rect 5502 14592 6090 14648
rect 6146 14592 6151 14648
rect 5441 14590 6151 14592
rect 5441 14587 5507 14590
rect 6085 14587 6151 14590
rect 18822 14588 18828 14652
rect 18892 14650 18898 14652
rect 18965 14650 19031 14653
rect 18892 14648 19031 14650
rect 18892 14592 18970 14648
rect 19026 14592 19031 14648
rect 18892 14590 19031 14592
rect 19934 14650 19994 14859
rect 20161 14786 20227 14789
rect 22320 14786 22800 14816
rect 20161 14784 22800 14786
rect 20161 14728 20166 14784
rect 20222 14728 22800 14784
rect 20161 14726 22800 14728
rect 20161 14723 20227 14726
rect 22320 14696 22800 14726
rect 20161 14650 20227 14653
rect 19934 14648 20227 14650
rect 19934 14592 20166 14648
rect 20222 14592 20227 14648
rect 19934 14590 20227 14592
rect 18892 14588 18898 14590
rect 18965 14587 19031 14590
rect 20161 14587 20227 14590
rect 11329 14514 11395 14517
rect 14038 14514 14044 14516
rect 11329 14512 14044 14514
rect 11329 14456 11334 14512
rect 11390 14456 14044 14512
rect 11329 14454 14044 14456
rect 11329 14451 11395 14454
rect 14038 14452 14044 14454
rect 14108 14514 14114 14516
rect 18137 14514 18203 14517
rect 14108 14512 18203 14514
rect 14108 14456 18142 14512
rect 18198 14456 18203 14512
rect 14108 14454 18203 14456
rect 14108 14452 14114 14454
rect 18137 14451 18203 14454
rect 18321 14514 18387 14517
rect 19926 14514 19932 14516
rect 18321 14512 19932 14514
rect 18321 14456 18326 14512
rect 18382 14456 19932 14512
rect 18321 14454 19932 14456
rect 18321 14451 18387 14454
rect 19926 14452 19932 14454
rect 19996 14452 20002 14516
rect 0 14378 480 14408
rect 1577 14378 1643 14381
rect 0 14376 1643 14378
rect 0 14320 1582 14376
rect 1638 14320 1643 14376
rect 0 14318 1643 14320
rect 0 14288 480 14318
rect 1577 14315 1643 14318
rect 2681 14378 2747 14381
rect 5625 14378 5691 14381
rect 2681 14376 5691 14378
rect 2681 14320 2686 14376
rect 2742 14320 5630 14376
rect 5686 14320 5691 14376
rect 2681 14318 5691 14320
rect 2681 14315 2747 14318
rect 5625 14315 5691 14318
rect 6085 14378 6151 14381
rect 11421 14378 11487 14381
rect 12893 14378 12959 14381
rect 6085 14376 12959 14378
rect 6085 14320 6090 14376
rect 6146 14320 11426 14376
rect 11482 14320 12898 14376
rect 12954 14320 12959 14376
rect 6085 14318 12959 14320
rect 6085 14315 6151 14318
rect 11421 14315 11487 14318
rect 12893 14315 12959 14318
rect 13670 14316 13676 14380
rect 13740 14378 13746 14380
rect 14089 14378 14155 14381
rect 13740 14376 14155 14378
rect 13740 14320 14094 14376
rect 14150 14320 14155 14376
rect 13740 14318 14155 14320
rect 13740 14316 13746 14318
rect 14089 14315 14155 14318
rect 15745 14378 15811 14381
rect 15878 14378 15884 14380
rect 15745 14376 15884 14378
rect 15745 14320 15750 14376
rect 15806 14320 15884 14376
rect 15745 14318 15884 14320
rect 15745 14315 15811 14318
rect 15878 14316 15884 14318
rect 15948 14316 15954 14380
rect 16614 14316 16620 14380
rect 16684 14378 16690 14380
rect 17401 14378 17467 14381
rect 18689 14378 18755 14381
rect 22320 14378 22800 14408
rect 16684 14376 18568 14378
rect 16684 14320 17406 14376
rect 17462 14320 18568 14376
rect 16684 14318 18568 14320
rect 16684 14316 16690 14318
rect 17401 14315 17467 14318
rect 12433 14242 12499 14245
rect 15745 14242 15811 14245
rect 12433 14240 15811 14242
rect 12433 14184 12438 14240
rect 12494 14184 15750 14240
rect 15806 14184 15811 14240
rect 12433 14182 15811 14184
rect 18508 14242 18568 14318
rect 18689 14376 22800 14378
rect 18689 14320 18694 14376
rect 18750 14320 22800 14376
rect 18689 14318 22800 14320
rect 18689 14315 18755 14318
rect 22320 14288 22800 14318
rect 19374 14242 19380 14244
rect 18508 14182 19380 14242
rect 12433 14179 12499 14182
rect 15745 14179 15811 14182
rect 19374 14180 19380 14182
rect 19444 14242 19450 14244
rect 19609 14242 19675 14245
rect 19444 14240 19675 14242
rect 19444 14184 19614 14240
rect 19670 14184 19675 14240
rect 19444 14182 19675 14184
rect 19444 14180 19450 14182
rect 19609 14179 19675 14182
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 19793 14108 19859 14109
rect 19742 14044 19748 14108
rect 19812 14106 19859 14108
rect 19812 14104 19904 14106
rect 19854 14048 19904 14104
rect 19812 14046 19904 14048
rect 19812 14044 19859 14046
rect 19793 14043 19859 14044
rect 0 13970 480 14000
rect 4245 13970 4311 13973
rect 7465 13972 7531 13973
rect 11145 13972 11211 13973
rect 0 13968 4311 13970
rect 0 13912 4250 13968
rect 4306 13912 4311 13968
rect 0 13910 4311 13912
rect 0 13880 480 13910
rect 4245 13907 4311 13910
rect 7414 13908 7420 13972
rect 7484 13970 7531 13972
rect 11094 13970 11100 13972
rect 7484 13968 7576 13970
rect 7526 13912 7576 13968
rect 7484 13910 7576 13912
rect 11018 13910 11100 13970
rect 11164 13970 11211 13972
rect 16941 13970 17007 13973
rect 11164 13968 17007 13970
rect 11206 13912 16946 13968
rect 17002 13912 17007 13968
rect 7484 13908 7531 13910
rect 11094 13908 11100 13910
rect 11164 13910 17007 13912
rect 11164 13908 11211 13910
rect 7465 13907 7531 13908
rect 11145 13907 11211 13908
rect 16941 13907 17007 13910
rect 21081 13970 21147 13973
rect 22320 13970 22800 14000
rect 21081 13968 22800 13970
rect 21081 13912 21086 13968
rect 21142 13912 22800 13968
rect 21081 13910 22800 13912
rect 21081 13907 21147 13910
rect 22320 13880 22800 13910
rect 2865 13836 2931 13837
rect 2814 13834 2820 13836
rect 2774 13774 2820 13834
rect 2884 13832 2931 13836
rect 2926 13776 2931 13832
rect 2814 13772 2820 13774
rect 2884 13772 2931 13776
rect 2865 13771 2931 13772
rect 6729 13834 6795 13837
rect 9857 13834 9923 13837
rect 6729 13832 9923 13834
rect 6729 13776 6734 13832
rect 6790 13776 9862 13832
rect 9918 13776 9923 13832
rect 6729 13774 9923 13776
rect 6729 13771 6795 13774
rect 9857 13771 9923 13774
rect 10910 13772 10916 13836
rect 10980 13834 10986 13836
rect 15193 13834 15259 13837
rect 10980 13832 15259 13834
rect 10980 13776 15198 13832
rect 15254 13776 15259 13832
rect 10980 13774 15259 13776
rect 10980 13772 10986 13774
rect 15193 13771 15259 13774
rect 16205 13834 16271 13837
rect 16982 13834 16988 13836
rect 16205 13832 16988 13834
rect 16205 13776 16210 13832
rect 16266 13776 16988 13832
rect 16205 13774 16988 13776
rect 16205 13771 16271 13774
rect 16982 13772 16988 13774
rect 17052 13772 17058 13836
rect 19425 13834 19491 13837
rect 19558 13834 19564 13836
rect 19425 13832 19564 13834
rect 19425 13776 19430 13832
rect 19486 13776 19564 13832
rect 19425 13774 19564 13776
rect 19425 13771 19491 13774
rect 19558 13772 19564 13774
rect 19628 13772 19634 13836
rect 11513 13698 11579 13701
rect 13854 13698 13860 13700
rect 11513 13696 13860 13698
rect 11513 13640 11518 13696
rect 11574 13640 13860 13696
rect 11513 13638 13860 13640
rect 11513 13635 11579 13638
rect 13854 13636 13860 13638
rect 13924 13636 13930 13700
rect 17534 13636 17540 13700
rect 17604 13698 17610 13700
rect 18873 13698 18939 13701
rect 17604 13696 18939 13698
rect 17604 13640 18878 13696
rect 18934 13640 18939 13696
rect 17604 13638 18939 13640
rect 17604 13636 17610 13638
rect 18873 13635 18939 13638
rect 7808 13632 8128 13633
rect 0 13562 480 13592
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 1669 13562 1735 13565
rect 0 13560 1735 13562
rect 0 13504 1674 13560
rect 1730 13504 1735 13560
rect 0 13502 1735 13504
rect 0 13472 480 13502
rect 1669 13499 1735 13502
rect 5625 13562 5691 13565
rect 5993 13562 6059 13565
rect 7097 13562 7163 13565
rect 5625 13560 7163 13562
rect 5625 13504 5630 13560
rect 5686 13504 5998 13560
rect 6054 13504 7102 13560
rect 7158 13504 7163 13560
rect 5625 13502 7163 13504
rect 5625 13499 5691 13502
rect 5993 13499 6059 13502
rect 7097 13499 7163 13502
rect 8334 13500 8340 13564
rect 8404 13562 8410 13564
rect 13077 13562 13143 13565
rect 8404 13560 13143 13562
rect 8404 13504 13082 13560
rect 13138 13504 13143 13560
rect 8404 13502 13143 13504
rect 8404 13500 8410 13502
rect 13077 13499 13143 13502
rect 15653 13564 15719 13565
rect 15653 13560 15700 13564
rect 15764 13562 15770 13564
rect 15653 13504 15658 13560
rect 15653 13500 15700 13504
rect 15764 13502 15810 13562
rect 15764 13500 15770 13502
rect 16798 13500 16804 13564
rect 16868 13562 16874 13564
rect 18045 13562 18111 13565
rect 19006 13562 19012 13564
rect 16868 13560 19012 13562
rect 16868 13504 18050 13560
rect 18106 13504 19012 13560
rect 16868 13502 19012 13504
rect 16868 13500 16874 13502
rect 15653 13499 15719 13500
rect 18045 13499 18111 13502
rect 19006 13500 19012 13502
rect 19076 13500 19082 13564
rect 19149 13562 19215 13565
rect 22320 13562 22800 13592
rect 19149 13560 22800 13562
rect 19149 13504 19154 13560
rect 19210 13504 22800 13560
rect 19149 13502 22800 13504
rect 19149 13499 19215 13502
rect 22320 13472 22800 13502
rect 5717 13426 5783 13429
rect 10593 13426 10659 13429
rect 20713 13426 20779 13429
rect 5717 13424 6378 13426
rect 5717 13368 5722 13424
rect 5778 13368 6378 13424
rect 5717 13366 6378 13368
rect 5717 13363 5783 13366
rect 6318 13292 6378 13366
rect 10593 13424 20779 13426
rect 10593 13368 10598 13424
rect 10654 13368 20718 13424
rect 20774 13368 20779 13424
rect 10593 13366 20779 13368
rect 10593 13363 10659 13366
rect 20713 13363 20779 13366
rect 6310 13228 6316 13292
rect 6380 13290 6386 13292
rect 7373 13290 7439 13293
rect 6380 13288 7439 13290
rect 6380 13232 7378 13288
rect 7434 13232 7439 13288
rect 6380 13230 7439 13232
rect 6380 13228 6386 13230
rect 7373 13227 7439 13230
rect 8201 13290 8267 13293
rect 8518 13290 8524 13292
rect 8201 13288 8524 13290
rect 8201 13232 8206 13288
rect 8262 13232 8524 13288
rect 8201 13230 8524 13232
rect 8201 13227 8267 13230
rect 8518 13228 8524 13230
rect 8588 13228 8594 13292
rect 8886 13228 8892 13292
rect 8956 13290 8962 13292
rect 15653 13290 15719 13293
rect 8956 13288 15719 13290
rect 8956 13232 15658 13288
rect 15714 13232 15719 13288
rect 8956 13230 15719 13232
rect 8956 13228 8962 13230
rect 15653 13227 15719 13230
rect 16062 13228 16068 13292
rect 16132 13290 16138 13292
rect 17033 13290 17099 13293
rect 16132 13288 17099 13290
rect 16132 13232 17038 13288
rect 17094 13232 17099 13288
rect 16132 13230 17099 13232
rect 16132 13228 16138 13230
rect 17033 13227 17099 13230
rect 17677 13290 17743 13293
rect 18781 13290 18847 13293
rect 17677 13288 18847 13290
rect 17677 13232 17682 13288
rect 17738 13232 18786 13288
rect 18842 13232 18847 13288
rect 17677 13230 18847 13232
rect 17677 13227 17743 13230
rect 18781 13227 18847 13230
rect 0 13154 480 13184
rect 2865 13154 2931 13157
rect 0 13152 2931 13154
rect 0 13096 2870 13152
rect 2926 13096 2931 13152
rect 0 13094 2931 13096
rect 0 13064 480 13094
rect 2865 13091 2931 13094
rect 10910 13092 10916 13156
rect 10980 13154 10986 13156
rect 11053 13154 11119 13157
rect 10980 13152 11119 13154
rect 10980 13096 11058 13152
rect 11114 13096 11119 13152
rect 10980 13094 11119 13096
rect 10980 13092 10986 13094
rect 11053 13091 11119 13094
rect 11973 13154 12039 13157
rect 16665 13154 16731 13157
rect 11973 13152 16731 13154
rect 11973 13096 11978 13152
rect 12034 13096 16670 13152
rect 16726 13096 16731 13152
rect 11973 13094 16731 13096
rect 11973 13091 12039 13094
rect 16665 13091 16731 13094
rect 18505 13154 18571 13157
rect 22320 13154 22800 13184
rect 18505 13152 22800 13154
rect 18505 13096 18510 13152
rect 18566 13096 22800 13152
rect 18505 13094 22800 13096
rect 18505 13091 18571 13094
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 22320 13064 22800 13094
rect 18104 13023 18424 13024
rect 4889 13018 4955 13021
rect 8937 13018 9003 13021
rect 10225 13020 10291 13021
rect 12985 13020 13051 13021
rect 9070 13018 9076 13020
rect 4889 13016 8816 13018
rect 4889 12960 4894 13016
rect 4950 12960 8816 13016
rect 4889 12958 8816 12960
rect 4889 12955 4955 12958
rect 1485 12882 1551 12885
rect 6085 12882 6151 12885
rect 1485 12880 6151 12882
rect 1485 12824 1490 12880
rect 1546 12824 6090 12880
rect 6146 12824 6151 12880
rect 1485 12822 6151 12824
rect 1485 12819 1551 12822
rect 6085 12819 6151 12822
rect 6729 12882 6795 12885
rect 7230 12882 7236 12884
rect 6729 12880 7236 12882
rect 6729 12824 6734 12880
rect 6790 12824 7236 12880
rect 6729 12822 7236 12824
rect 6729 12819 6795 12822
rect 7230 12820 7236 12822
rect 7300 12820 7306 12884
rect 8756 12882 8816 12958
rect 8937 13016 9076 13018
rect 8937 12960 8942 13016
rect 8998 12960 9076 13016
rect 8937 12958 9076 12960
rect 8937 12955 9003 12958
rect 9070 12956 9076 12958
rect 9140 12956 9146 13020
rect 10174 12956 10180 13020
rect 10244 13018 10291 13020
rect 10244 13016 10336 13018
rect 10286 12960 10336 13016
rect 10244 12958 10336 12960
rect 10244 12956 10291 12958
rect 12934 12956 12940 13020
rect 13004 13018 13051 13020
rect 14917 13018 14983 13021
rect 13004 13016 13096 13018
rect 13046 12960 13096 13016
rect 13004 12958 13096 12960
rect 14230 13016 14983 13018
rect 14230 12960 14922 13016
rect 14978 12960 14983 13016
rect 14230 12958 14983 12960
rect 13004 12956 13051 12958
rect 10225 12955 10291 12956
rect 12985 12955 13051 12956
rect 10133 12882 10199 12885
rect 8756 12880 10199 12882
rect 8756 12824 10138 12880
rect 10194 12824 10199 12880
rect 8756 12822 10199 12824
rect 10133 12819 10199 12822
rect 11513 12882 11579 12885
rect 14230 12882 14290 12958
rect 14917 12955 14983 12958
rect 15285 13020 15351 13021
rect 15285 13016 15332 13020
rect 15396 13018 15402 13020
rect 15745 13018 15811 13021
rect 16297 13018 16363 13021
rect 15285 12960 15290 13016
rect 15285 12956 15332 12960
rect 15396 12958 15442 13018
rect 15745 13016 16363 13018
rect 15745 12960 15750 13016
rect 15806 12960 16302 13016
rect 16358 12960 16363 13016
rect 15745 12958 16363 12960
rect 15396 12956 15402 12958
rect 15285 12955 15351 12956
rect 15745 12955 15811 12958
rect 16297 12955 16363 12958
rect 17125 13020 17191 13021
rect 17125 13016 17172 13020
rect 17236 13018 17242 13020
rect 18689 13018 18755 13021
rect 20069 13018 20135 13021
rect 17125 12960 17130 13016
rect 17125 12956 17172 12960
rect 17236 12958 17282 13018
rect 18689 13016 20135 13018
rect 18689 12960 18694 13016
rect 18750 12960 20074 13016
rect 20130 12960 20135 13016
rect 18689 12958 20135 12960
rect 17236 12956 17242 12958
rect 17125 12955 17191 12956
rect 18689 12955 18755 12958
rect 20069 12955 20135 12958
rect 11513 12880 14290 12882
rect 11513 12824 11518 12880
rect 11574 12824 14290 12880
rect 11513 12822 14290 12824
rect 14365 12882 14431 12885
rect 15326 12882 15332 12884
rect 14365 12880 15332 12882
rect 14365 12824 14370 12880
rect 14426 12824 15332 12880
rect 14365 12822 15332 12824
rect 11513 12819 11579 12822
rect 14365 12819 14431 12822
rect 15326 12820 15332 12822
rect 15396 12820 15402 12884
rect 19793 12882 19859 12885
rect 15472 12880 19859 12882
rect 15472 12824 19798 12880
rect 19854 12824 19859 12880
rect 15472 12822 19859 12824
rect 0 12746 480 12776
rect 1945 12746 2011 12749
rect 15472 12746 15532 12822
rect 19793 12819 19859 12822
rect 0 12686 1410 12746
rect 0 12656 480 12686
rect 1350 12610 1410 12686
rect 1945 12744 15532 12746
rect 1945 12688 1950 12744
rect 2006 12688 15532 12744
rect 1945 12686 15532 12688
rect 17033 12746 17099 12749
rect 18781 12746 18847 12749
rect 17033 12744 18847 12746
rect 17033 12688 17038 12744
rect 17094 12688 18786 12744
rect 18842 12688 18847 12744
rect 17033 12686 18847 12688
rect 1945 12683 2011 12686
rect 17033 12683 17099 12686
rect 18781 12683 18847 12686
rect 19190 12684 19196 12748
rect 19260 12746 19266 12748
rect 19333 12746 19399 12749
rect 22320 12746 22800 12776
rect 19260 12744 19399 12746
rect 19260 12688 19338 12744
rect 19394 12688 19399 12744
rect 19260 12686 19399 12688
rect 19260 12684 19266 12686
rect 19333 12683 19399 12686
rect 19750 12686 22800 12746
rect 3877 12610 3943 12613
rect 1350 12608 3943 12610
rect 1350 12552 3882 12608
rect 3938 12552 3943 12608
rect 1350 12550 3943 12552
rect 3877 12547 3943 12550
rect 5165 12610 5231 12613
rect 6678 12610 6684 12612
rect 5165 12608 6684 12610
rect 5165 12552 5170 12608
rect 5226 12552 6684 12608
rect 5165 12550 6684 12552
rect 5165 12547 5231 12550
rect 6678 12548 6684 12550
rect 6748 12548 6754 12612
rect 9806 12548 9812 12612
rect 9876 12610 9882 12612
rect 10133 12610 10199 12613
rect 9876 12608 10199 12610
rect 9876 12552 10138 12608
rect 10194 12552 10199 12608
rect 9876 12550 10199 12552
rect 9876 12548 9882 12550
rect 10133 12547 10199 12550
rect 11881 12610 11947 12613
rect 14457 12610 14523 12613
rect 11881 12608 14523 12610
rect 11881 12552 11886 12608
rect 11942 12552 14462 12608
rect 14518 12552 14523 12608
rect 11881 12550 14523 12552
rect 11881 12547 11947 12550
rect 14457 12547 14523 12550
rect 16665 12610 16731 12613
rect 17401 12610 17467 12613
rect 16665 12608 17467 12610
rect 16665 12552 16670 12608
rect 16726 12552 17406 12608
rect 17462 12552 17467 12608
rect 16665 12550 17467 12552
rect 16665 12547 16731 12550
rect 17401 12547 17467 12550
rect 17718 12548 17724 12612
rect 17788 12610 17794 12612
rect 18689 12610 18755 12613
rect 19057 12612 19123 12613
rect 19006 12610 19012 12612
rect 17788 12608 18755 12610
rect 17788 12552 18694 12608
rect 18750 12552 18755 12608
rect 17788 12550 18755 12552
rect 18966 12550 19012 12610
rect 19076 12608 19123 12612
rect 19118 12552 19123 12608
rect 17788 12548 17794 12550
rect 18689 12547 18755 12550
rect 19006 12548 19012 12550
rect 19076 12548 19123 12552
rect 19057 12547 19123 12548
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 6862 12412 6868 12476
rect 6932 12474 6938 12476
rect 7097 12474 7163 12477
rect 6932 12472 7163 12474
rect 6932 12416 7102 12472
rect 7158 12416 7163 12472
rect 6932 12414 7163 12416
rect 6932 12412 6938 12414
rect 7097 12411 7163 12414
rect 8753 12474 8819 12477
rect 8753 12472 10104 12474
rect 8753 12416 8758 12472
rect 8814 12416 10104 12472
rect 8753 12414 10104 12416
rect 8753 12411 8819 12414
rect 0 12338 480 12368
rect 3049 12338 3115 12341
rect 0 12336 3115 12338
rect 0 12280 3054 12336
rect 3110 12280 3115 12336
rect 0 12278 3115 12280
rect 0 12248 480 12278
rect 3049 12275 3115 12278
rect 5165 12338 5231 12341
rect 6678 12338 6684 12340
rect 5165 12336 6684 12338
rect 5165 12280 5170 12336
rect 5226 12280 6684 12336
rect 5165 12278 6684 12280
rect 5165 12275 5231 12278
rect 6678 12276 6684 12278
rect 6748 12276 6754 12340
rect 8109 12338 8175 12341
rect 7008 12336 8175 12338
rect 7008 12280 8114 12336
rect 8170 12280 8175 12336
rect 7008 12278 8175 12280
rect 3969 12202 4035 12205
rect 7008 12202 7068 12278
rect 8109 12275 8175 12278
rect 8293 12338 8359 12341
rect 8702 12338 8708 12340
rect 8293 12336 8708 12338
rect 8293 12280 8298 12336
rect 8354 12280 8708 12336
rect 8293 12278 8708 12280
rect 8293 12275 8359 12278
rect 8702 12276 8708 12278
rect 8772 12276 8778 12340
rect 9213 12338 9279 12341
rect 8894 12336 9279 12338
rect 8894 12280 9218 12336
rect 9274 12280 9279 12336
rect 8894 12278 9279 12280
rect 7465 12204 7531 12205
rect 7414 12202 7420 12204
rect 3969 12200 7068 12202
rect 3969 12144 3974 12200
rect 4030 12144 7068 12200
rect 3969 12142 7068 12144
rect 7374 12142 7420 12202
rect 7484 12200 7531 12204
rect 7526 12144 7531 12200
rect 3969 12139 4035 12142
rect 7414 12140 7420 12142
rect 7484 12140 7531 12144
rect 8702 12140 8708 12204
rect 8772 12202 8778 12204
rect 8894 12202 8954 12278
rect 9213 12275 9279 12278
rect 9581 12338 9647 12341
rect 9806 12338 9812 12340
rect 9581 12336 9812 12338
rect 9581 12280 9586 12336
rect 9642 12280 9812 12336
rect 9581 12278 9812 12280
rect 9581 12275 9647 12278
rect 9806 12276 9812 12278
rect 9876 12276 9882 12340
rect 10044 12338 10104 12414
rect 10174 12412 10180 12476
rect 10244 12474 10250 12476
rect 10593 12474 10659 12477
rect 10244 12472 10659 12474
rect 10244 12416 10598 12472
rect 10654 12416 10659 12472
rect 10244 12414 10659 12416
rect 10244 12412 10250 12414
rect 10593 12411 10659 12414
rect 11830 12412 11836 12476
rect 11900 12474 11906 12476
rect 12157 12474 12223 12477
rect 11900 12472 12223 12474
rect 11900 12416 12162 12472
rect 12218 12416 12223 12472
rect 11900 12414 12223 12416
rect 11900 12412 11906 12414
rect 12157 12411 12223 12414
rect 16021 12474 16087 12477
rect 16614 12474 16620 12476
rect 16021 12472 16620 12474
rect 16021 12416 16026 12472
rect 16082 12416 16620 12472
rect 16021 12414 16620 12416
rect 16021 12411 16087 12414
rect 16614 12412 16620 12414
rect 16684 12412 16690 12476
rect 17861 12474 17927 12477
rect 19750 12474 19810 12686
rect 22320 12656 22800 12686
rect 17861 12472 19810 12474
rect 17861 12416 17866 12472
rect 17922 12416 19810 12472
rect 17861 12414 19810 12416
rect 19885 12476 19951 12477
rect 19885 12472 19932 12476
rect 19996 12474 20002 12476
rect 19885 12416 19890 12472
rect 17861 12411 17927 12414
rect 19885 12412 19932 12416
rect 19996 12414 20042 12474
rect 19996 12412 20002 12414
rect 19885 12411 19951 12412
rect 11513 12338 11579 12341
rect 10044 12336 11579 12338
rect 10044 12280 11518 12336
rect 11574 12280 11579 12336
rect 10044 12278 11579 12280
rect 11513 12275 11579 12278
rect 13353 12338 13419 12341
rect 13670 12338 13676 12340
rect 13353 12336 13676 12338
rect 13353 12280 13358 12336
rect 13414 12280 13676 12336
rect 13353 12278 13676 12280
rect 13353 12275 13419 12278
rect 13670 12276 13676 12278
rect 13740 12276 13746 12340
rect 14089 12338 14155 12341
rect 16062 12338 16068 12340
rect 14089 12336 16068 12338
rect 14089 12280 14094 12336
rect 14150 12280 16068 12336
rect 14089 12278 16068 12280
rect 14089 12275 14155 12278
rect 16062 12276 16068 12278
rect 16132 12276 16138 12340
rect 16481 12338 16547 12341
rect 22320 12338 22800 12368
rect 16481 12336 22800 12338
rect 16481 12280 16486 12336
rect 16542 12280 22800 12336
rect 16481 12278 22800 12280
rect 16481 12275 16547 12278
rect 22320 12248 22800 12278
rect 8772 12142 8954 12202
rect 8772 12140 8778 12142
rect 9254 12140 9260 12204
rect 9324 12202 9330 12204
rect 10409 12202 10475 12205
rect 16757 12202 16823 12205
rect 9324 12200 16823 12202
rect 9324 12144 10414 12200
rect 10470 12144 16762 12200
rect 16818 12144 16823 12200
rect 9324 12142 16823 12144
rect 9324 12140 9330 12142
rect 7465 12139 7531 12140
rect 10409 12139 10475 12142
rect 16757 12139 16823 12142
rect 18505 12202 18571 12205
rect 18822 12202 18828 12204
rect 18505 12200 18828 12202
rect 18505 12144 18510 12200
rect 18566 12144 18828 12200
rect 18505 12142 18828 12144
rect 18505 12139 18571 12142
rect 18822 12140 18828 12142
rect 18892 12140 18898 12204
rect 19190 12140 19196 12204
rect 19260 12202 19266 12204
rect 19885 12202 19951 12205
rect 19260 12200 19951 12202
rect 19260 12144 19890 12200
rect 19946 12144 19951 12200
rect 19260 12142 19951 12144
rect 19260 12140 19266 12142
rect 19885 12139 19951 12142
rect 3233 12068 3299 12069
rect 3182 12004 3188 12068
rect 3252 12066 3299 12068
rect 3252 12064 3344 12066
rect 3294 12008 3344 12064
rect 3252 12006 3344 12008
rect 3252 12004 3299 12006
rect 7046 12004 7052 12068
rect 7116 12066 7122 12068
rect 7281 12066 7347 12069
rect 7116 12064 7347 12066
rect 7116 12008 7286 12064
rect 7342 12008 7347 12064
rect 7116 12006 7347 12008
rect 7116 12004 7122 12006
rect 3233 12003 3299 12004
rect 7281 12003 7347 12006
rect 7557 12066 7623 12069
rect 8569 12066 8635 12069
rect 17350 12066 17356 12068
rect 7557 12064 8635 12066
rect 7557 12008 7562 12064
rect 7618 12008 8574 12064
rect 8630 12008 8635 12064
rect 7557 12006 8635 12008
rect 7557 12003 7623 12006
rect 8569 12003 8635 12006
rect 12252 12006 17356 12066
rect 4376 12000 4696 12001
rect 0 11930 480 11960
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 3141 11930 3207 11933
rect 0 11928 3207 11930
rect 0 11872 3146 11928
rect 3202 11872 3207 11928
rect 0 11870 3207 11872
rect 0 11840 480 11870
rect 3141 11867 3207 11870
rect 8569 11930 8635 11933
rect 9397 11930 9463 11933
rect 8569 11928 9463 11930
rect 8569 11872 8574 11928
rect 8630 11872 9402 11928
rect 9458 11872 9463 11928
rect 8569 11870 9463 11872
rect 8569 11867 8635 11870
rect 9397 11867 9463 11870
rect 5901 11794 5967 11797
rect 12252 11794 12312 12006
rect 17350 12004 17356 12006
rect 17420 12004 17426 12068
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 13077 11930 13143 11933
rect 13353 11930 13419 11933
rect 13721 11930 13787 11933
rect 15101 11930 15167 11933
rect 13077 11928 13419 11930
rect 13077 11872 13082 11928
rect 13138 11872 13358 11928
rect 13414 11872 13419 11928
rect 13077 11870 13419 11872
rect 13077 11867 13143 11870
rect 13353 11867 13419 11870
rect 13494 11928 15167 11930
rect 13494 11872 13726 11928
rect 13782 11872 15106 11928
rect 15162 11872 15167 11928
rect 13494 11870 15167 11872
rect 5901 11792 12312 11794
rect 5901 11736 5906 11792
rect 5962 11736 12312 11792
rect 5901 11734 12312 11736
rect 5901 11731 5967 11734
rect 12382 11732 12388 11796
rect 12452 11794 12458 11796
rect 13494 11794 13554 11870
rect 13721 11867 13787 11870
rect 15101 11867 15167 11870
rect 15837 11930 15903 11933
rect 16849 11930 16915 11933
rect 15837 11928 16915 11930
rect 15837 11872 15842 11928
rect 15898 11872 16854 11928
rect 16910 11872 16915 11928
rect 15837 11870 16915 11872
rect 15837 11867 15903 11870
rect 16849 11867 16915 11870
rect 19149 11930 19215 11933
rect 19374 11930 19380 11932
rect 19149 11928 19380 11930
rect 19149 11872 19154 11928
rect 19210 11872 19380 11928
rect 19149 11870 19380 11872
rect 19149 11867 19215 11870
rect 19374 11868 19380 11870
rect 19444 11868 19450 11932
rect 19609 11930 19675 11933
rect 22320 11930 22800 11960
rect 19609 11928 22800 11930
rect 19609 11872 19614 11928
rect 19670 11872 22800 11928
rect 19609 11870 22800 11872
rect 19609 11867 19675 11870
rect 22320 11840 22800 11870
rect 12452 11734 13554 11794
rect 13997 11794 14063 11797
rect 19425 11794 19491 11797
rect 13997 11792 19491 11794
rect 13997 11736 14002 11792
rect 14058 11736 19430 11792
rect 19486 11736 19491 11792
rect 13997 11734 19491 11736
rect 12452 11732 12458 11734
rect 13997 11731 14063 11734
rect 19425 11731 19491 11734
rect 0 11658 480 11688
rect 3601 11658 3667 11661
rect 0 11656 3667 11658
rect 0 11600 3606 11656
rect 3662 11600 3667 11656
rect 0 11598 3667 11600
rect 0 11568 480 11598
rect 3601 11595 3667 11598
rect 7230 11596 7236 11660
rect 7300 11658 7306 11660
rect 7465 11658 7531 11661
rect 9029 11658 9095 11661
rect 9581 11658 9647 11661
rect 10409 11658 10475 11661
rect 12014 11658 12020 11660
rect 7300 11656 7531 11658
rect 7300 11600 7470 11656
rect 7526 11600 7531 11656
rect 7300 11598 7531 11600
rect 7300 11596 7306 11598
rect 7465 11595 7531 11598
rect 7652 11656 9095 11658
rect 7652 11600 9034 11656
rect 9090 11600 9095 11656
rect 7652 11598 9095 11600
rect 9540 11656 9828 11658
rect 9540 11600 9586 11656
rect 9642 11600 9828 11656
rect 9540 11598 9828 11600
rect 3693 11522 3759 11525
rect 7652 11522 7712 11598
rect 9029 11595 9095 11598
rect 9581 11595 9647 11598
rect 3693 11520 7712 11522
rect 3693 11464 3698 11520
rect 3754 11464 7712 11520
rect 3693 11462 7712 11464
rect 3693 11459 3759 11462
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 9622 11324 9628 11388
rect 9692 11386 9698 11388
rect 9768 11386 9828 11598
rect 10409 11656 12020 11658
rect 10409 11600 10414 11656
rect 10470 11600 12020 11656
rect 10409 11598 12020 11600
rect 10409 11595 10475 11598
rect 12014 11596 12020 11598
rect 12084 11596 12090 11660
rect 12157 11658 12223 11661
rect 14549 11658 14615 11661
rect 12157 11656 14615 11658
rect 12157 11600 12162 11656
rect 12218 11600 14554 11656
rect 14610 11600 14615 11656
rect 12157 11598 14615 11600
rect 12157 11595 12223 11598
rect 14549 11595 14615 11598
rect 15837 11658 15903 11661
rect 18045 11658 18111 11661
rect 15837 11656 18111 11658
rect 15837 11600 15842 11656
rect 15898 11600 18050 11656
rect 18106 11600 18111 11656
rect 15837 11598 18111 11600
rect 15837 11595 15903 11598
rect 18045 11595 18111 11598
rect 21081 11658 21147 11661
rect 22320 11658 22800 11688
rect 21081 11656 22800 11658
rect 21081 11600 21086 11656
rect 21142 11600 22800 11656
rect 21081 11598 22800 11600
rect 21081 11595 21147 11598
rect 22320 11568 22800 11598
rect 12157 11522 12223 11525
rect 13486 11522 13492 11524
rect 12157 11520 13492 11522
rect 12157 11464 12162 11520
rect 12218 11464 13492 11520
rect 12157 11462 13492 11464
rect 12157 11459 12223 11462
rect 13486 11460 13492 11462
rect 13556 11460 13562 11524
rect 15561 11522 15627 11525
rect 18413 11522 18479 11525
rect 19425 11522 19491 11525
rect 15561 11520 18479 11522
rect 15561 11464 15566 11520
rect 15622 11464 18418 11520
rect 18474 11464 18479 11520
rect 15561 11462 18479 11464
rect 15561 11459 15627 11462
rect 18413 11459 18479 11462
rect 18646 11520 19491 11522
rect 18646 11464 19430 11520
rect 19486 11464 19491 11520
rect 18646 11462 19491 11464
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 9692 11326 9828 11386
rect 9949 11388 10015 11389
rect 9949 11384 9996 11388
rect 10060 11386 10066 11388
rect 10869 11386 10935 11389
rect 14089 11386 14155 11389
rect 9949 11328 9954 11384
rect 9692 11324 9698 11326
rect 9949 11324 9996 11328
rect 10060 11326 10106 11386
rect 10869 11384 14155 11386
rect 10869 11328 10874 11384
rect 10930 11328 14094 11384
rect 14150 11328 14155 11384
rect 10869 11326 14155 11328
rect 10060 11324 10066 11326
rect 9949 11323 10015 11324
rect 10869 11323 10935 11326
rect 14089 11323 14155 11326
rect 15469 11386 15535 11389
rect 15694 11386 15700 11388
rect 15469 11384 15700 11386
rect 15469 11328 15474 11384
rect 15530 11328 15700 11384
rect 15469 11326 15700 11328
rect 15469 11323 15535 11326
rect 15694 11324 15700 11326
rect 15764 11386 15770 11388
rect 15837 11386 15903 11389
rect 15764 11384 15903 11386
rect 15764 11328 15842 11384
rect 15898 11328 15903 11384
rect 15764 11326 15903 11328
rect 15764 11324 15770 11326
rect 15837 11323 15903 11326
rect 16021 11386 16087 11389
rect 18646 11386 18706 11462
rect 19425 11459 19491 11462
rect 16021 11384 18706 11386
rect 16021 11328 16026 11384
rect 16082 11328 18706 11384
rect 16021 11326 18706 11328
rect 16021 11323 16087 11326
rect 0 11250 480 11280
rect 1577 11250 1643 11253
rect 13261 11250 13327 11253
rect 0 11248 1643 11250
rect 0 11192 1582 11248
rect 1638 11192 1643 11248
rect 0 11190 1643 11192
rect 0 11160 480 11190
rect 1577 11187 1643 11190
rect 10872 11248 13327 11250
rect 10872 11192 13266 11248
rect 13322 11192 13327 11248
rect 10872 11190 13327 11192
rect 4838 11052 4844 11116
rect 4908 11114 4914 11116
rect 5073 11114 5139 11117
rect 4908 11112 5139 11114
rect 4908 11056 5078 11112
rect 5134 11056 5139 11112
rect 4908 11054 5139 11056
rect 4908 11052 4914 11054
rect 5073 11051 5139 11054
rect 8661 11114 8727 11117
rect 9438 11114 9444 11116
rect 8661 11112 9444 11114
rect 8661 11056 8666 11112
rect 8722 11056 9444 11112
rect 8661 11054 9444 11056
rect 8661 11051 8727 11054
rect 9438 11052 9444 11054
rect 9508 11114 9514 11116
rect 10872 11114 10932 11190
rect 13261 11187 13327 11190
rect 13721 11250 13787 11253
rect 15101 11250 15167 11253
rect 18822 11250 18828 11252
rect 13721 11248 14428 11250
rect 13721 11192 13726 11248
rect 13782 11192 14428 11248
rect 13721 11190 14428 11192
rect 13721 11187 13787 11190
rect 14368 11117 14428 11190
rect 15101 11248 18828 11250
rect 15101 11192 15106 11248
rect 15162 11192 18828 11248
rect 15101 11190 18828 11192
rect 15101 11187 15167 11190
rect 18822 11188 18828 11190
rect 18892 11188 18898 11252
rect 19006 11188 19012 11252
rect 19076 11250 19082 11252
rect 19149 11250 19215 11253
rect 19076 11248 19215 11250
rect 19076 11192 19154 11248
rect 19210 11192 19215 11248
rect 19076 11190 19215 11192
rect 19076 11188 19082 11190
rect 19149 11187 19215 11190
rect 21265 11250 21331 11253
rect 22320 11250 22800 11280
rect 21265 11248 22800 11250
rect 21265 11192 21270 11248
rect 21326 11192 22800 11248
rect 21265 11190 22800 11192
rect 21265 11187 21331 11190
rect 22320 11160 22800 11190
rect 12750 11114 12756 11116
rect 9508 11054 10932 11114
rect 11102 11054 12756 11114
rect 9508 11052 9514 11054
rect 4838 10916 4844 10980
rect 4908 10978 4914 10980
rect 5257 10978 5323 10981
rect 4908 10976 5323 10978
rect 4908 10920 5262 10976
rect 5318 10920 5323 10976
rect 4908 10918 5323 10920
rect 4908 10916 4914 10918
rect 5257 10915 5323 10918
rect 5390 10916 5396 10980
rect 5460 10978 5466 10980
rect 6637 10978 6703 10981
rect 5460 10976 6703 10978
rect 5460 10920 6642 10976
rect 6698 10920 6703 10976
rect 5460 10918 6703 10920
rect 5460 10916 5466 10918
rect 6637 10915 6703 10918
rect 9029 10978 9095 10981
rect 11102 10978 11162 11054
rect 12750 11052 12756 11054
rect 12820 11052 12826 11116
rect 13721 11114 13787 11117
rect 14365 11114 14431 11117
rect 20161 11114 20227 11117
rect 13721 11112 14290 11114
rect 13721 11056 13726 11112
rect 13782 11056 14290 11112
rect 13721 11054 14290 11056
rect 13721 11051 13787 11054
rect 9029 10976 11162 10978
rect 9029 10920 9034 10976
rect 9090 10920 11162 10976
rect 9029 10918 11162 10920
rect 9029 10915 9095 10918
rect 11646 10916 11652 10980
rect 11716 10978 11722 10980
rect 13670 10978 13676 10980
rect 11716 10918 13676 10978
rect 11716 10916 11722 10918
rect 13670 10916 13676 10918
rect 13740 10916 13746 10980
rect 14230 10978 14290 11054
rect 14365 11112 20227 11114
rect 14365 11056 14370 11112
rect 14426 11056 20166 11112
rect 20222 11056 20227 11112
rect 14365 11054 20227 11056
rect 14365 11051 14431 11054
rect 20161 11051 20227 11054
rect 15009 10978 15075 10981
rect 16757 10980 16823 10981
rect 16757 10978 16804 10980
rect 14230 10976 15075 10978
rect 14230 10920 15014 10976
rect 15070 10920 15075 10976
rect 14230 10918 15075 10920
rect 16712 10976 16804 10978
rect 16712 10920 16762 10976
rect 16712 10918 16804 10920
rect 15009 10915 15075 10918
rect 16757 10916 16804 10918
rect 16868 10916 16874 10980
rect 16757 10915 16823 10916
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 3693 10842 3759 10845
rect 0 10840 3759 10842
rect 0 10784 3698 10840
rect 3754 10784 3759 10840
rect 0 10782 3759 10784
rect 0 10752 480 10782
rect 3693 10779 3759 10782
rect 4889 10842 4955 10845
rect 8477 10842 8543 10845
rect 4889 10840 8543 10842
rect 4889 10784 4894 10840
rect 4950 10784 8482 10840
rect 8538 10784 8543 10840
rect 4889 10782 8543 10784
rect 4889 10779 4955 10782
rect 8477 10779 8543 10782
rect 12157 10842 12223 10845
rect 17677 10842 17743 10845
rect 22320 10842 22800 10872
rect 12157 10840 17743 10842
rect 12157 10784 12162 10840
rect 12218 10784 17682 10840
rect 17738 10784 17743 10840
rect 12157 10782 17743 10784
rect 12157 10779 12223 10782
rect 17677 10779 17743 10782
rect 19014 10782 22800 10842
rect 6821 10706 6887 10709
rect 7189 10706 7255 10709
rect 8334 10706 8340 10708
rect 6821 10704 8340 10706
rect 6821 10648 6826 10704
rect 6882 10648 7194 10704
rect 7250 10648 8340 10704
rect 6821 10646 8340 10648
rect 6821 10643 6887 10646
rect 7189 10643 7255 10646
rect 8334 10644 8340 10646
rect 8404 10644 8410 10708
rect 9305 10706 9371 10709
rect 13813 10706 13879 10709
rect 9305 10704 13879 10706
rect 9305 10648 9310 10704
rect 9366 10648 13818 10704
rect 13874 10648 13879 10704
rect 9305 10646 13879 10648
rect 9305 10643 9371 10646
rect 13813 10643 13879 10646
rect 16982 10644 16988 10708
rect 17052 10706 17058 10708
rect 18781 10706 18847 10709
rect 17052 10704 18847 10706
rect 17052 10648 18786 10704
rect 18842 10648 18847 10704
rect 17052 10646 18847 10648
rect 17052 10644 17058 10646
rect 18781 10643 18847 10646
rect 1853 10570 1919 10573
rect 5901 10570 5967 10573
rect 9949 10570 10015 10573
rect 11145 10570 11211 10573
rect 16297 10570 16363 10573
rect 1853 10568 5967 10570
rect 1853 10512 1858 10568
rect 1914 10512 5906 10568
rect 5962 10512 5967 10568
rect 1853 10510 5967 10512
rect 1853 10507 1919 10510
rect 5901 10507 5967 10510
rect 7652 10510 8264 10570
rect 0 10434 480 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 480 10374
rect 4061 10371 4127 10374
rect 6177 10298 6243 10301
rect 7652 10298 7712 10510
rect 8204 10434 8264 10510
rect 9949 10568 11211 10570
rect 9949 10512 9954 10568
rect 10010 10512 11150 10568
rect 11206 10512 11211 10568
rect 9949 10510 11211 10512
rect 9949 10507 10015 10510
rect 11145 10507 11211 10510
rect 11286 10568 16363 10570
rect 11286 10512 16302 10568
rect 16358 10512 16363 10568
rect 11286 10510 16363 10512
rect 11286 10434 11346 10510
rect 16297 10507 16363 10510
rect 17166 10508 17172 10572
rect 17236 10570 17242 10572
rect 19014 10570 19074 10782
rect 22320 10752 22800 10782
rect 17236 10510 19074 10570
rect 17236 10508 17242 10510
rect 8204 10374 11346 10434
rect 11513 10434 11579 10437
rect 14181 10434 14247 10437
rect 11513 10432 14247 10434
rect 11513 10376 11518 10432
rect 11574 10376 14186 10432
rect 14242 10376 14247 10432
rect 11513 10374 14247 10376
rect 11513 10371 11579 10374
rect 14181 10371 14247 10374
rect 16246 10372 16252 10436
rect 16316 10434 16322 10436
rect 18137 10434 18203 10437
rect 20110 10434 20116 10436
rect 16316 10432 18203 10434
rect 16316 10376 18142 10432
rect 18198 10376 18203 10432
rect 16316 10374 18203 10376
rect 16316 10372 16322 10374
rect 18137 10371 18203 10374
rect 18462 10374 20116 10434
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 12065 10298 12131 10301
rect 6177 10296 7712 10298
rect 6177 10240 6182 10296
rect 6238 10240 7712 10296
rect 6177 10238 7712 10240
rect 9078 10296 12131 10298
rect 9078 10240 12070 10296
rect 12126 10240 12131 10296
rect 9078 10238 12131 10240
rect 6177 10235 6243 10238
rect 6913 10162 6979 10165
rect 6870 10160 6979 10162
rect 6870 10104 6918 10160
rect 6974 10104 6979 10160
rect 6870 10099 6979 10104
rect 8109 10162 8175 10165
rect 9078 10162 9138 10238
rect 12065 10235 12131 10238
rect 12433 10298 12499 10301
rect 12617 10298 12683 10301
rect 13629 10298 13695 10301
rect 12433 10296 13695 10298
rect 12433 10240 12438 10296
rect 12494 10240 12622 10296
rect 12678 10240 13634 10296
rect 13690 10240 13695 10296
rect 12433 10238 13695 10240
rect 12433 10235 12499 10238
rect 12617 10235 12683 10238
rect 13629 10235 13695 10238
rect 15878 10236 15884 10300
rect 15948 10298 15954 10300
rect 18462 10298 18522 10374
rect 20110 10372 20116 10374
rect 20180 10434 20186 10436
rect 22320 10434 22800 10464
rect 20180 10374 22800 10434
rect 20180 10372 20186 10374
rect 22320 10344 22800 10374
rect 15948 10238 18522 10298
rect 15948 10236 15954 10238
rect 8109 10160 9138 10162
rect 8109 10104 8114 10160
rect 8170 10104 9138 10160
rect 8109 10102 9138 10104
rect 9213 10162 9279 10165
rect 12566 10162 12572 10164
rect 9213 10160 12572 10162
rect 9213 10104 9218 10160
rect 9274 10104 12572 10160
rect 9213 10102 12572 10104
rect 8109 10099 8175 10102
rect 9213 10099 9279 10102
rect 12566 10100 12572 10102
rect 12636 10100 12642 10164
rect 12750 10100 12756 10164
rect 12820 10162 12826 10164
rect 14365 10162 14431 10165
rect 12820 10160 14431 10162
rect 12820 10104 14370 10160
rect 14426 10104 14431 10160
rect 12820 10102 14431 10104
rect 12820 10100 12826 10102
rect 14365 10099 14431 10102
rect 14641 10162 14707 10165
rect 16941 10162 17007 10165
rect 14641 10160 17007 10162
rect 14641 10104 14646 10160
rect 14702 10104 16946 10160
rect 17002 10104 17007 10160
rect 14641 10102 17007 10104
rect 14641 10099 14707 10102
rect 16941 10099 17007 10102
rect 18137 10162 18203 10165
rect 19057 10162 19123 10165
rect 19926 10162 19932 10164
rect 18137 10160 19932 10162
rect 18137 10104 18142 10160
rect 18198 10104 19062 10160
rect 19118 10104 19932 10160
rect 18137 10102 19932 10104
rect 18137 10099 18203 10102
rect 19057 10099 19123 10102
rect 19926 10100 19932 10102
rect 19996 10100 20002 10164
rect 0 10026 480 10056
rect 5717 10026 5783 10029
rect 0 10024 5783 10026
rect 0 9968 5722 10024
rect 5778 9968 5783 10024
rect 0 9966 5783 9968
rect 0 9936 480 9966
rect 5717 9963 5783 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 0 9618 480 9648
rect 0 9558 3480 9618
rect 0 9528 480 9558
rect 3420 9482 3480 9558
rect 3550 9556 3556 9620
rect 3620 9618 3626 9620
rect 6361 9618 6427 9621
rect 3620 9616 6427 9618
rect 3620 9560 6366 9616
rect 6422 9560 6427 9616
rect 3620 9558 6427 9560
rect 3620 9556 3626 9558
rect 6361 9555 6427 9558
rect 6870 9485 6930 10099
rect 8702 9964 8708 10028
rect 8772 10026 8778 10028
rect 9029 10026 9095 10029
rect 10317 10028 10383 10029
rect 10317 10026 10364 10028
rect 8772 10024 9095 10026
rect 8772 9968 9034 10024
rect 9090 9968 9095 10024
rect 8772 9966 9095 9968
rect 10272 10024 10364 10026
rect 10428 10026 10434 10028
rect 12065 10026 12131 10029
rect 16941 10026 17007 10029
rect 10272 9968 10322 10024
rect 10272 9966 10364 9968
rect 8772 9964 8778 9966
rect 9029 9963 9095 9966
rect 10317 9964 10364 9966
rect 10428 9966 11944 10026
rect 10428 9964 10434 9966
rect 10317 9963 10383 9964
rect 8201 9890 8267 9893
rect 9857 9890 9923 9893
rect 11697 9892 11763 9893
rect 10726 9890 10732 9892
rect 8201 9888 10732 9890
rect 8201 9832 8206 9888
rect 8262 9832 9862 9888
rect 9918 9832 10732 9888
rect 8201 9830 10732 9832
rect 8201 9827 8267 9830
rect 9857 9827 9923 9830
rect 10726 9828 10732 9830
rect 10796 9828 10802 9892
rect 11646 9828 11652 9892
rect 11716 9890 11763 9892
rect 11884 9890 11944 9966
rect 12065 10024 17007 10026
rect 12065 9968 12070 10024
rect 12126 9968 16946 10024
rect 17002 9968 17007 10024
rect 12065 9966 17007 9968
rect 12065 9963 12131 9966
rect 16941 9963 17007 9966
rect 18045 10026 18111 10029
rect 20345 10026 20411 10029
rect 22320 10026 22800 10056
rect 18045 10024 22800 10026
rect 18045 9968 18050 10024
rect 18106 9968 20350 10024
rect 20406 9968 22800 10024
rect 18045 9966 22800 9968
rect 18045 9963 18111 9966
rect 20345 9963 20411 9966
rect 22320 9936 22800 9966
rect 15837 9890 15903 9893
rect 11716 9888 11808 9890
rect 11758 9832 11808 9888
rect 11716 9830 11808 9832
rect 11884 9888 15903 9890
rect 11884 9832 15842 9888
rect 15898 9832 15903 9888
rect 11884 9830 15903 9832
rect 11716 9828 11763 9830
rect 11697 9827 11763 9828
rect 15837 9827 15903 9830
rect 17585 9890 17651 9893
rect 17861 9890 17927 9893
rect 17585 9888 17927 9890
rect 17585 9832 17590 9888
rect 17646 9832 17866 9888
rect 17922 9832 17927 9888
rect 17585 9830 17927 9832
rect 17585 9827 17651 9830
rect 17861 9827 17927 9830
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 8661 9754 8727 9757
rect 10777 9754 10843 9757
rect 8661 9752 10843 9754
rect 8661 9696 8666 9752
rect 8722 9696 10782 9752
rect 10838 9696 10843 9752
rect 8661 9694 10843 9696
rect 8661 9691 8727 9694
rect 10777 9691 10843 9694
rect 11789 9754 11855 9757
rect 12750 9754 12756 9756
rect 11789 9752 12756 9754
rect 11789 9696 11794 9752
rect 11850 9696 12756 9752
rect 11789 9694 12756 9696
rect 11789 9691 11855 9694
rect 12750 9692 12756 9694
rect 12820 9692 12826 9756
rect 12893 9754 12959 9757
rect 13537 9754 13603 9757
rect 12893 9752 17970 9754
rect 12893 9696 12898 9752
rect 12954 9696 13542 9752
rect 13598 9696 17970 9752
rect 12893 9694 17970 9696
rect 12893 9691 12959 9694
rect 13537 9691 13603 9694
rect 9213 9618 9279 9621
rect 15929 9618 15995 9621
rect 9213 9616 15995 9618
rect 9213 9560 9218 9616
rect 9274 9560 15934 9616
rect 15990 9560 15995 9616
rect 9213 9558 15995 9560
rect 9213 9555 9279 9558
rect 15929 9555 15995 9558
rect 17125 9618 17191 9621
rect 17534 9618 17540 9620
rect 17125 9616 17540 9618
rect 17125 9560 17130 9616
rect 17186 9560 17540 9616
rect 17125 9558 17540 9560
rect 17125 9555 17191 9558
rect 17534 9556 17540 9558
rect 17604 9556 17610 9620
rect 17910 9618 17970 9694
rect 22320 9618 22800 9648
rect 17910 9558 22800 9618
rect 22320 9528 22800 9558
rect 4705 9482 4771 9485
rect 3420 9480 4771 9482
rect 3420 9424 4710 9480
rect 4766 9424 4771 9480
rect 3420 9422 4771 9424
rect 4705 9419 4771 9422
rect 5901 9482 5967 9485
rect 6361 9482 6427 9485
rect 5901 9480 6427 9482
rect 5901 9424 5906 9480
rect 5962 9424 6366 9480
rect 6422 9424 6427 9480
rect 5901 9422 6427 9424
rect 5901 9419 5967 9422
rect 6361 9419 6427 9422
rect 6821 9480 6930 9485
rect 9857 9482 9923 9485
rect 6821 9424 6826 9480
rect 6882 9424 6930 9480
rect 6821 9422 6930 9424
rect 7054 9480 9923 9482
rect 7054 9424 9862 9480
rect 9918 9424 9923 9480
rect 7054 9422 9923 9424
rect 6821 9419 6887 9422
rect 1853 9346 1919 9349
rect 5390 9346 5396 9348
rect 1853 9344 5396 9346
rect 1853 9288 1858 9344
rect 1914 9288 5396 9344
rect 1853 9286 5396 9288
rect 1853 9283 1919 9286
rect 5390 9284 5396 9286
rect 5460 9346 5466 9348
rect 6862 9346 6868 9348
rect 5460 9286 6868 9346
rect 5460 9284 5466 9286
rect 6862 9284 6868 9286
rect 6932 9346 6938 9348
rect 7054 9346 7114 9422
rect 9857 9419 9923 9422
rect 10041 9482 10107 9485
rect 11329 9482 11395 9485
rect 10041 9480 11395 9482
rect 10041 9424 10046 9480
rect 10102 9424 11334 9480
rect 11390 9424 11395 9480
rect 10041 9422 11395 9424
rect 10041 9419 10107 9422
rect 11329 9419 11395 9422
rect 11697 9482 11763 9485
rect 19374 9482 19380 9484
rect 11697 9480 19380 9482
rect 11697 9424 11702 9480
rect 11758 9424 19380 9480
rect 11697 9422 19380 9424
rect 11697 9419 11763 9422
rect 19374 9420 19380 9422
rect 19444 9420 19450 9484
rect 6932 9286 7114 9346
rect 8293 9346 8359 9349
rect 17585 9348 17651 9349
rect 14038 9346 14044 9348
rect 8293 9344 14044 9346
rect 8293 9288 8298 9344
rect 8354 9288 14044 9344
rect 8293 9286 14044 9288
rect 6932 9284 6938 9286
rect 8293 9283 8359 9286
rect 14038 9284 14044 9286
rect 14108 9284 14114 9348
rect 17534 9346 17540 9348
rect 17494 9286 17540 9346
rect 17604 9344 17651 9348
rect 17646 9288 17651 9344
rect 17534 9284 17540 9286
rect 17604 9284 17651 9288
rect 17718 9284 17724 9348
rect 17788 9346 17794 9348
rect 18597 9346 18663 9349
rect 17788 9344 18663 9346
rect 17788 9288 18602 9344
rect 18658 9288 18663 9344
rect 17788 9286 18663 9288
rect 17788 9284 17794 9286
rect 17585 9283 17651 9284
rect 18597 9283 18663 9286
rect 18822 9284 18828 9348
rect 18892 9346 18898 9348
rect 19701 9346 19767 9349
rect 18892 9344 19767 9346
rect 18892 9288 19706 9344
rect 19762 9288 19767 9344
rect 18892 9286 19767 9288
rect 18892 9284 18898 9286
rect 19701 9283 19767 9286
rect 7808 9280 8128 9281
rect 0 9210 480 9240
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 2037 9210 2103 9213
rect 0 9208 2103 9210
rect 0 9152 2042 9208
rect 2098 9152 2103 9208
rect 0 9150 2103 9152
rect 0 9120 480 9150
rect 2037 9147 2103 9150
rect 3049 9210 3115 9213
rect 3182 9210 3188 9212
rect 3049 9208 3188 9210
rect 3049 9152 3054 9208
rect 3110 9152 3188 9208
rect 3049 9150 3188 9152
rect 3049 9147 3115 9150
rect 3182 9148 3188 9150
rect 3252 9148 3258 9212
rect 8201 9210 8267 9213
rect 14406 9210 14412 9212
rect 8201 9208 14412 9210
rect 8201 9152 8206 9208
rect 8262 9152 14412 9208
rect 8201 9150 14412 9152
rect 8201 9147 8267 9150
rect 14406 9148 14412 9150
rect 14476 9148 14482 9212
rect 15510 9148 15516 9212
rect 15580 9210 15586 9212
rect 15929 9210 15995 9213
rect 22320 9210 22800 9240
rect 15580 9208 15995 9210
rect 15580 9152 15934 9208
rect 15990 9152 15995 9208
rect 15580 9150 15995 9152
rect 15580 9148 15586 9150
rect 15929 9147 15995 9150
rect 16070 9150 22800 9210
rect 5165 9074 5231 9077
rect 4110 9072 5231 9074
rect 4110 9016 5170 9072
rect 5226 9016 5231 9072
rect 4110 9014 5231 9016
rect 0 8802 480 8832
rect 4110 8802 4170 9014
rect 5165 9011 5231 9014
rect 6678 9012 6684 9076
rect 6748 9074 6754 9076
rect 6821 9074 6887 9077
rect 6748 9072 6887 9074
rect 6748 9016 6826 9072
rect 6882 9016 6887 9072
rect 6748 9014 6887 9016
rect 6748 9012 6754 9014
rect 6821 9011 6887 9014
rect 7189 9074 7255 9077
rect 7189 9072 9000 9074
rect 7189 9016 7194 9072
rect 7250 9016 9000 9072
rect 7189 9014 9000 9016
rect 7189 9011 7255 9014
rect 5073 8938 5139 8941
rect 8293 8938 8359 8941
rect 5073 8936 8359 8938
rect 5073 8880 5078 8936
rect 5134 8880 8298 8936
rect 8354 8880 8359 8936
rect 5073 8878 8359 8880
rect 8940 8938 9000 9014
rect 9070 9012 9076 9076
rect 9140 9074 9146 9076
rect 9489 9074 9555 9077
rect 9140 9072 9555 9074
rect 9140 9016 9494 9072
rect 9550 9016 9555 9072
rect 9140 9014 9555 9016
rect 9140 9012 9146 9014
rect 9489 9011 9555 9014
rect 9857 9074 9923 9077
rect 13629 9074 13695 9077
rect 16070 9074 16130 9150
rect 22320 9120 22800 9150
rect 9857 9072 13554 9074
rect 9857 9016 9862 9072
rect 9918 9016 13554 9072
rect 9857 9014 13554 9016
rect 9857 9011 9923 9014
rect 9213 8938 9279 8941
rect 10409 8938 10475 8941
rect 8940 8936 9279 8938
rect 8940 8880 9218 8936
rect 9274 8880 9279 8936
rect 8940 8878 9279 8880
rect 5073 8875 5139 8878
rect 8293 8875 8359 8878
rect 9213 8875 9279 8878
rect 10182 8936 10475 8938
rect 10182 8880 10414 8936
rect 10470 8880 10475 8936
rect 10182 8878 10475 8880
rect 0 8742 4170 8802
rect 5625 8802 5691 8805
rect 6637 8802 6703 8805
rect 6862 8802 6868 8804
rect 5625 8800 6868 8802
rect 5625 8744 5630 8800
rect 5686 8744 6642 8800
rect 6698 8744 6868 8800
rect 5625 8742 6868 8744
rect 0 8712 480 8742
rect 5625 8739 5691 8742
rect 6637 8739 6703 8742
rect 6862 8740 6868 8742
rect 6932 8740 6938 8804
rect 7230 8740 7236 8804
rect 7300 8802 7306 8804
rect 7373 8802 7439 8805
rect 7300 8800 7439 8802
rect 7300 8744 7378 8800
rect 7434 8744 7439 8800
rect 7300 8742 7439 8744
rect 7300 8740 7306 8742
rect 7373 8739 7439 8742
rect 8017 8802 8083 8805
rect 10041 8802 10107 8805
rect 8017 8800 10107 8802
rect 8017 8744 8022 8800
rect 8078 8744 10046 8800
rect 10102 8744 10107 8800
rect 8017 8742 10107 8744
rect 8017 8739 8083 8742
rect 10041 8739 10107 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 10182 8666 10242 8878
rect 10409 8875 10475 8878
rect 11329 8938 11395 8941
rect 13302 8938 13308 8940
rect 11329 8936 13308 8938
rect 11329 8880 11334 8936
rect 11390 8880 13308 8936
rect 11329 8878 13308 8880
rect 11329 8875 11395 8878
rect 13302 8876 13308 8878
rect 13372 8876 13378 8940
rect 13494 8938 13554 9014
rect 13629 9072 16130 9074
rect 13629 9016 13634 9072
rect 13690 9016 16130 9072
rect 13629 9014 16130 9016
rect 16389 9074 16455 9077
rect 16614 9074 16620 9076
rect 16389 9072 16620 9074
rect 16389 9016 16394 9072
rect 16450 9016 16620 9072
rect 16389 9014 16620 9016
rect 13629 9011 13695 9014
rect 16389 9011 16455 9014
rect 16614 9012 16620 9014
rect 16684 9012 16690 9076
rect 18597 9074 18663 9077
rect 19190 9074 19196 9076
rect 18597 9072 19196 9074
rect 18597 9016 18602 9072
rect 18658 9016 19196 9072
rect 18597 9014 19196 9016
rect 18597 9011 18663 9014
rect 19190 9012 19196 9014
rect 19260 9074 19266 9076
rect 19701 9074 19767 9077
rect 19260 9072 19767 9074
rect 19260 9016 19706 9072
rect 19762 9016 19767 9072
rect 19260 9014 19767 9016
rect 19260 9012 19266 9014
rect 19701 9011 19767 9014
rect 15510 8938 15516 8940
rect 13494 8878 15516 8938
rect 15510 8876 15516 8878
rect 15580 8876 15586 8940
rect 15929 8938 15995 8941
rect 21357 8938 21423 8941
rect 15929 8936 21423 8938
rect 15929 8880 15934 8936
rect 15990 8880 21362 8936
rect 21418 8880 21423 8936
rect 15929 8878 21423 8880
rect 15929 8875 15995 8878
rect 21357 8875 21423 8878
rect 12198 8740 12204 8804
rect 12268 8802 12274 8804
rect 12985 8802 13051 8805
rect 12268 8800 13051 8802
rect 12268 8744 12990 8800
rect 13046 8744 13051 8800
rect 12268 8742 13051 8744
rect 12268 8740 12274 8742
rect 12985 8739 13051 8742
rect 13353 8802 13419 8805
rect 17953 8802 18019 8805
rect 13353 8800 18019 8802
rect 13353 8744 13358 8800
rect 13414 8744 17958 8800
rect 18014 8744 18019 8800
rect 13353 8742 18019 8744
rect 13353 8739 13419 8742
rect 17953 8739 18019 8742
rect 18505 8802 18571 8805
rect 22320 8802 22800 8832
rect 18505 8800 22800 8802
rect 18505 8744 18510 8800
rect 18566 8744 22800 8800
rect 18505 8742 22800 8744
rect 18505 8739 18571 8742
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 22320 8712 22800 8742
rect 18104 8671 18424 8672
rect 5030 8606 10242 8666
rect 10317 8666 10383 8669
rect 10542 8666 10548 8668
rect 10317 8664 10548 8666
rect 10317 8608 10322 8664
rect 10378 8608 10548 8664
rect 10317 8606 10548 8608
rect 3141 8530 3207 8533
rect 5030 8530 5090 8606
rect 10317 8603 10383 8606
rect 10542 8604 10548 8606
rect 10612 8604 10618 8668
rect 10910 8604 10916 8668
rect 10980 8666 10986 8668
rect 11053 8666 11119 8669
rect 10980 8664 11119 8666
rect 10980 8608 11058 8664
rect 11114 8608 11119 8664
rect 10980 8606 11119 8608
rect 10980 8604 10986 8606
rect 11053 8603 11119 8606
rect 12525 8666 12591 8669
rect 13486 8666 13492 8668
rect 12525 8664 13492 8666
rect 12525 8608 12530 8664
rect 12586 8608 13492 8664
rect 12525 8606 13492 8608
rect 12525 8603 12591 8606
rect 13486 8604 13492 8606
rect 13556 8604 13562 8668
rect 14038 8604 14044 8668
rect 14108 8666 14114 8668
rect 14273 8666 14339 8669
rect 15009 8666 15075 8669
rect 14108 8664 15075 8666
rect 14108 8608 14278 8664
rect 14334 8608 15014 8664
rect 15070 8608 15075 8664
rect 14108 8606 15075 8608
rect 14108 8604 14114 8606
rect 14273 8603 14339 8606
rect 15009 8603 15075 8606
rect 15561 8666 15627 8669
rect 15561 8664 18016 8666
rect 15561 8608 15566 8664
rect 15622 8608 18016 8664
rect 15561 8606 18016 8608
rect 15561 8603 15627 8606
rect 3141 8528 5090 8530
rect 3141 8472 3146 8528
rect 3202 8472 5090 8528
rect 3141 8470 5090 8472
rect 5349 8530 5415 8533
rect 6177 8530 6243 8533
rect 5349 8528 6243 8530
rect 5349 8472 5354 8528
rect 5410 8472 6182 8528
rect 6238 8472 6243 8528
rect 5349 8470 6243 8472
rect 3141 8467 3207 8470
rect 5349 8467 5415 8470
rect 6177 8467 6243 8470
rect 6729 8530 6795 8533
rect 11830 8530 11836 8532
rect 6729 8528 11836 8530
rect 6729 8472 6734 8528
rect 6790 8472 11836 8528
rect 6729 8470 11836 8472
rect 6729 8467 6795 8470
rect 11830 8468 11836 8470
rect 11900 8468 11906 8532
rect 12433 8530 12499 8533
rect 15561 8530 15627 8533
rect 16941 8530 17007 8533
rect 12433 8528 17007 8530
rect 12433 8472 12438 8528
rect 12494 8472 15566 8528
rect 15622 8472 16946 8528
rect 17002 8472 17007 8528
rect 12433 8470 17007 8472
rect 17956 8530 18016 8606
rect 18822 8604 18828 8668
rect 18892 8666 18898 8668
rect 21081 8666 21147 8669
rect 18892 8664 21147 8666
rect 18892 8608 21086 8664
rect 21142 8608 21147 8664
rect 18892 8606 21147 8608
rect 18892 8604 18898 8606
rect 21081 8603 21147 8606
rect 19425 8530 19491 8533
rect 17956 8528 19491 8530
rect 17956 8472 19430 8528
rect 19486 8472 19491 8528
rect 17956 8470 19491 8472
rect 12433 8467 12499 8470
rect 15561 8467 15627 8470
rect 16941 8467 17007 8470
rect 19425 8467 19491 8470
rect 0 8394 480 8424
rect 4705 8394 4771 8397
rect 0 8392 4771 8394
rect 0 8336 4710 8392
rect 4766 8336 4771 8392
rect 0 8334 4771 8336
rect 0 8304 480 8334
rect 4705 8331 4771 8334
rect 5165 8392 5231 8397
rect 5165 8336 5170 8392
rect 5226 8336 5231 8392
rect 5165 8331 5231 8336
rect 6177 8394 6243 8397
rect 10409 8394 10475 8397
rect 11094 8394 11100 8396
rect 6177 8392 11100 8394
rect 6177 8336 6182 8392
rect 6238 8336 10414 8392
rect 10470 8336 11100 8392
rect 6177 8334 11100 8336
rect 6177 8331 6243 8334
rect 10409 8331 10475 8334
rect 11094 8332 11100 8334
rect 11164 8332 11170 8396
rect 11421 8394 11487 8397
rect 13118 8394 13124 8396
rect 11421 8392 13124 8394
rect 11421 8336 11426 8392
rect 11482 8336 13124 8392
rect 11421 8334 13124 8336
rect 11421 8331 11487 8334
rect 13118 8332 13124 8334
rect 13188 8332 13194 8396
rect 16021 8394 16087 8397
rect 16205 8394 16271 8397
rect 16021 8392 16271 8394
rect 16021 8336 16026 8392
rect 16082 8336 16210 8392
rect 16266 8336 16271 8392
rect 16021 8334 16271 8336
rect 16021 8331 16087 8334
rect 16205 8331 16271 8334
rect 16941 8394 17007 8397
rect 22320 8394 22800 8424
rect 16941 8392 22800 8394
rect 16941 8336 16946 8392
rect 17002 8336 22800 8392
rect 16941 8334 22800 8336
rect 16941 8331 17007 8334
rect 5168 8122 5228 8331
rect 22320 8304 22800 8334
rect 6361 8258 6427 8261
rect 6821 8258 6887 8261
rect 9029 8258 9095 8261
rect 13813 8258 13879 8261
rect 6361 8256 6887 8258
rect 6361 8200 6366 8256
rect 6422 8200 6826 8256
rect 6882 8200 6887 8256
rect 6361 8198 6887 8200
rect 6361 8195 6427 8198
rect 6821 8195 6887 8198
rect 8204 8256 13879 8258
rect 8204 8200 9034 8256
rect 9090 8200 13818 8256
rect 13874 8200 13879 8256
rect 8204 8198 13879 8200
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 7598 8122 7604 8124
rect 5168 8062 7604 8122
rect 7598 8060 7604 8062
rect 7668 8060 7674 8124
rect 0 7986 480 8016
rect 8204 7986 8264 8198
rect 9029 8195 9095 8198
rect 13813 8195 13879 8198
rect 15653 8258 15719 8261
rect 17033 8258 17099 8261
rect 18689 8258 18755 8261
rect 15653 8256 16084 8258
rect 15653 8200 15658 8256
rect 15714 8200 16084 8256
rect 15653 8198 16084 8200
rect 15653 8195 15719 8198
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 8661 8122 8727 8125
rect 9857 8122 9923 8125
rect 10501 8124 10567 8125
rect 9990 8122 9996 8124
rect 8661 8120 9690 8122
rect 8661 8064 8666 8120
rect 8722 8064 9690 8120
rect 8661 8062 9690 8064
rect 8661 8059 8727 8062
rect 0 7926 8264 7986
rect 8477 7986 8543 7989
rect 9070 7986 9076 7988
rect 8477 7984 9076 7986
rect 8477 7928 8482 7984
rect 8538 7928 9076 7984
rect 8477 7926 9076 7928
rect 0 7896 480 7926
rect 8477 7923 8543 7926
rect 9070 7924 9076 7926
rect 9140 7924 9146 7988
rect 9630 7986 9690 8062
rect 9857 8120 9996 8122
rect 9857 8064 9862 8120
rect 9918 8064 9996 8120
rect 9857 8062 9996 8064
rect 9857 8059 9923 8062
rect 9990 8060 9996 8062
rect 10060 8060 10066 8124
rect 10501 8122 10548 8124
rect 10456 8120 10548 8122
rect 10456 8064 10506 8120
rect 10456 8062 10548 8064
rect 10501 8060 10548 8062
rect 10612 8060 10618 8124
rect 11237 8122 11303 8125
rect 13077 8122 13143 8125
rect 11237 8120 13143 8122
rect 11237 8064 11242 8120
rect 11298 8064 13082 8120
rect 13138 8064 13143 8120
rect 11237 8062 13143 8064
rect 10501 8059 10567 8060
rect 11237 8059 11303 8062
rect 13077 8059 13143 8062
rect 15326 8060 15332 8124
rect 15396 8122 15402 8124
rect 15396 8062 15900 8122
rect 15396 8060 15402 8062
rect 15653 7986 15719 7989
rect 9630 7984 15719 7986
rect 9630 7928 15658 7984
rect 15714 7928 15719 7984
rect 9630 7926 15719 7928
rect 15653 7923 15719 7926
rect 3417 7850 3483 7853
rect 10317 7850 10383 7853
rect 10593 7850 10659 7853
rect 3417 7848 10383 7850
rect 3417 7792 3422 7848
rect 3478 7792 10322 7848
rect 10378 7792 10383 7848
rect 3417 7790 10383 7792
rect 3417 7787 3483 7790
rect 10317 7787 10383 7790
rect 10550 7848 10659 7850
rect 10550 7792 10598 7848
rect 10654 7792 10659 7848
rect 10550 7787 10659 7792
rect 10726 7788 10732 7852
rect 10796 7850 10802 7852
rect 11881 7850 11947 7853
rect 15469 7850 15535 7853
rect 10796 7790 11714 7850
rect 10796 7788 10802 7790
rect 0 7714 480 7744
rect 4061 7714 4127 7717
rect 0 7712 4127 7714
rect 0 7656 4066 7712
rect 4122 7656 4127 7712
rect 0 7654 4127 7656
rect 0 7624 480 7654
rect 4061 7651 4127 7654
rect 7649 7714 7715 7717
rect 10550 7714 10610 7787
rect 7649 7712 10610 7714
rect 7649 7656 7654 7712
rect 7710 7656 10610 7712
rect 7649 7654 10610 7656
rect 7649 7651 7715 7654
rect 10910 7652 10916 7716
rect 10980 7714 10986 7716
rect 11053 7714 11119 7717
rect 10980 7712 11119 7714
rect 10980 7656 11058 7712
rect 11114 7656 11119 7712
rect 10980 7654 11119 7656
rect 10980 7652 10986 7654
rect 11053 7651 11119 7654
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 6453 7578 6519 7581
rect 10685 7578 10751 7581
rect 6453 7576 10751 7578
rect 6453 7520 6458 7576
rect 6514 7520 10690 7576
rect 10746 7520 10751 7576
rect 6453 7518 10751 7520
rect 11654 7578 11714 7790
rect 11881 7848 15535 7850
rect 11881 7792 11886 7848
rect 11942 7792 15474 7848
rect 15530 7792 15535 7848
rect 11881 7790 15535 7792
rect 15840 7850 15900 8062
rect 16024 7986 16084 8198
rect 17033 8256 18755 8258
rect 17033 8200 17038 8256
rect 17094 8200 18694 8256
rect 18750 8200 18755 8256
rect 17033 8198 18755 8200
rect 17033 8195 17099 8198
rect 18689 8195 18755 8198
rect 18822 8196 18828 8260
rect 18892 8196 18898 8260
rect 19198 8198 20730 8258
rect 18229 8122 18295 8125
rect 18830 8122 18890 8196
rect 18229 8120 18890 8122
rect 18229 8064 18234 8120
rect 18290 8064 18890 8120
rect 18229 8062 18890 8064
rect 18229 8059 18295 8062
rect 19198 7986 19258 8198
rect 19333 8124 19399 8125
rect 19333 8120 19380 8124
rect 19444 8122 19450 8124
rect 19333 8064 19338 8120
rect 19333 8060 19380 8064
rect 19444 8062 19490 8122
rect 19444 8060 19450 8062
rect 19333 8059 19399 8060
rect 16024 7926 19258 7986
rect 19333 7986 19399 7989
rect 20110 7986 20116 7988
rect 19333 7984 20116 7986
rect 19333 7928 19338 7984
rect 19394 7928 20116 7984
rect 19333 7926 20116 7928
rect 19333 7923 19399 7926
rect 20110 7924 20116 7926
rect 20180 7924 20186 7988
rect 20670 7986 20730 8198
rect 22320 7986 22800 8016
rect 20670 7926 22800 7986
rect 22320 7896 22800 7926
rect 19977 7850 20043 7853
rect 15840 7848 20043 7850
rect 15840 7792 19982 7848
rect 20038 7792 20043 7848
rect 15840 7790 20043 7792
rect 11881 7787 11947 7790
rect 15469 7787 15535 7790
rect 19977 7787 20043 7790
rect 13813 7714 13879 7717
rect 15745 7714 15811 7717
rect 13813 7712 15811 7714
rect 13813 7656 13818 7712
rect 13874 7656 15750 7712
rect 15806 7656 15811 7712
rect 13813 7654 15811 7656
rect 13813 7651 13879 7654
rect 15745 7651 15811 7654
rect 17033 7714 17099 7717
rect 17166 7714 17172 7716
rect 17033 7712 17172 7714
rect 17033 7656 17038 7712
rect 17094 7656 17172 7712
rect 17033 7654 17172 7656
rect 17033 7651 17099 7654
rect 17166 7652 17172 7654
rect 17236 7652 17242 7716
rect 18689 7714 18755 7717
rect 19241 7714 19307 7717
rect 22320 7714 22800 7744
rect 18689 7712 19307 7714
rect 18689 7656 18694 7712
rect 18750 7656 19246 7712
rect 19302 7656 19307 7712
rect 18689 7654 19307 7656
rect 18689 7651 18755 7654
rect 19241 7651 19307 7654
rect 19382 7654 22800 7714
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 12893 7578 12959 7581
rect 11654 7576 12959 7578
rect 11654 7520 12898 7576
rect 12954 7520 12959 7576
rect 11654 7518 12959 7520
rect 6453 7515 6519 7518
rect 10685 7515 10751 7518
rect 12893 7515 12959 7518
rect 13353 7578 13419 7581
rect 13670 7578 13676 7580
rect 13353 7576 13676 7578
rect 13353 7520 13358 7576
rect 13414 7520 13676 7576
rect 13353 7518 13676 7520
rect 13353 7515 13419 7518
rect 13670 7516 13676 7518
rect 13740 7516 13746 7580
rect 14089 7578 14155 7581
rect 15326 7578 15332 7580
rect 14089 7576 15332 7578
rect 14089 7520 14094 7576
rect 14150 7520 15332 7576
rect 14089 7518 15332 7520
rect 14089 7515 14155 7518
rect 15326 7516 15332 7518
rect 15396 7516 15402 7580
rect 16021 7578 16087 7581
rect 17493 7578 17559 7581
rect 16021 7576 17559 7578
rect 16021 7520 16026 7576
rect 16082 7520 17498 7576
rect 17554 7520 17559 7576
rect 16021 7518 17559 7520
rect 16021 7515 16087 7518
rect 17493 7515 17559 7518
rect 18597 7578 18663 7581
rect 19006 7578 19012 7580
rect 18597 7576 19012 7578
rect 18597 7520 18602 7576
rect 18658 7520 19012 7576
rect 18597 7518 19012 7520
rect 18597 7515 18663 7518
rect 19006 7516 19012 7518
rect 19076 7516 19082 7580
rect 1669 7442 1735 7445
rect 4838 7442 4844 7444
rect 1669 7440 4844 7442
rect 1669 7384 1674 7440
rect 1730 7384 4844 7440
rect 1669 7382 4844 7384
rect 1669 7379 1735 7382
rect 4838 7380 4844 7382
rect 4908 7380 4914 7444
rect 7465 7442 7531 7445
rect 18689 7442 18755 7445
rect 7465 7440 18755 7442
rect 7465 7384 7470 7440
rect 7526 7384 18694 7440
rect 18750 7384 18755 7440
rect 7465 7382 18755 7384
rect 7465 7379 7531 7382
rect 18689 7379 18755 7382
rect 0 7306 480 7336
rect 5809 7306 5875 7309
rect 0 7304 5875 7306
rect 0 7248 5814 7304
rect 5870 7248 5875 7304
rect 0 7246 5875 7248
rect 0 7216 480 7246
rect 5809 7243 5875 7246
rect 6545 7306 6611 7309
rect 15142 7306 15148 7308
rect 6545 7304 15148 7306
rect 6545 7248 6550 7304
rect 6606 7248 15148 7304
rect 6545 7246 15148 7248
rect 6545 7243 6611 7246
rect 15142 7244 15148 7246
rect 15212 7244 15218 7308
rect 19382 7306 19442 7654
rect 22320 7624 22800 7654
rect 19701 7578 19767 7581
rect 19926 7578 19932 7580
rect 19701 7576 19932 7578
rect 19701 7520 19706 7576
rect 19762 7520 19932 7576
rect 19701 7518 19932 7520
rect 19701 7515 19767 7518
rect 19926 7516 19932 7518
rect 19996 7516 20002 7580
rect 19517 7442 19583 7445
rect 20805 7442 20871 7445
rect 19517 7440 20871 7442
rect 19517 7384 19522 7440
rect 19578 7384 20810 7440
rect 20866 7384 20871 7440
rect 19517 7382 20871 7384
rect 19517 7379 19583 7382
rect 20805 7379 20871 7382
rect 15288 7246 19442 7306
rect 19517 7304 19583 7309
rect 19517 7248 19522 7304
rect 19578 7248 19583 7304
rect 7649 7170 7715 7173
rect 2086 7168 7715 7170
rect 2086 7112 7654 7168
rect 7710 7112 7715 7168
rect 2086 7110 7715 7112
rect 0 6898 480 6928
rect 2086 6898 2146 7110
rect 7649 7107 7715 7110
rect 8334 7108 8340 7172
rect 8404 7170 8410 7172
rect 9305 7170 9371 7173
rect 8404 7168 9371 7170
rect 8404 7112 9310 7168
rect 9366 7112 9371 7168
rect 8404 7110 9371 7112
rect 8404 7108 8410 7110
rect 9305 7107 9371 7110
rect 11145 7170 11211 7173
rect 12382 7170 12388 7172
rect 11145 7168 12388 7170
rect 11145 7112 11150 7168
rect 11206 7112 12388 7168
rect 11145 7110 12388 7112
rect 11145 7107 11211 7110
rect 12382 7108 12388 7110
rect 12452 7108 12458 7172
rect 12525 7170 12591 7173
rect 12934 7170 12940 7172
rect 12525 7168 12940 7170
rect 12525 7112 12530 7168
rect 12586 7112 12940 7168
rect 12525 7110 12940 7112
rect 12525 7107 12591 7110
rect 12934 7108 12940 7110
rect 13004 7108 13010 7172
rect 13302 7108 13308 7172
rect 13372 7170 13378 7172
rect 13721 7170 13787 7173
rect 13372 7168 13787 7170
rect 13372 7112 13726 7168
rect 13782 7112 13787 7168
rect 13372 7110 13787 7112
rect 13372 7108 13378 7110
rect 13721 7107 13787 7110
rect 13854 7108 13860 7172
rect 13924 7170 13930 7172
rect 14457 7170 14523 7173
rect 13924 7168 14523 7170
rect 13924 7112 14462 7168
rect 14518 7112 14523 7168
rect 13924 7110 14523 7112
rect 13924 7108 13930 7110
rect 14457 7107 14523 7110
rect 15101 7170 15167 7173
rect 15288 7170 15348 7246
rect 19517 7243 19583 7248
rect 19977 7306 20043 7309
rect 22320 7306 22800 7336
rect 19977 7304 22800 7306
rect 19977 7248 19982 7304
rect 20038 7248 22800 7304
rect 19977 7246 22800 7248
rect 19977 7243 20043 7246
rect 15101 7168 15348 7170
rect 15101 7112 15106 7168
rect 15162 7112 15348 7168
rect 15101 7110 15348 7112
rect 15745 7170 15811 7173
rect 19149 7170 19215 7173
rect 19374 7170 19380 7172
rect 15745 7168 19074 7170
rect 15745 7112 15750 7168
rect 15806 7112 19074 7168
rect 15745 7110 19074 7112
rect 15101 7107 15167 7110
rect 15745 7107 15811 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 3734 6972 3740 7036
rect 3804 7034 3810 7036
rect 5533 7034 5599 7037
rect 3804 7032 5599 7034
rect 3804 6976 5538 7032
rect 5594 6976 5599 7032
rect 3804 6974 5599 6976
rect 3804 6972 3810 6974
rect 5533 6971 5599 6974
rect 6177 7034 6243 7037
rect 6310 7034 6316 7036
rect 6177 7032 6316 7034
rect 6177 6976 6182 7032
rect 6238 6976 6316 7032
rect 6177 6974 6316 6976
rect 6177 6971 6243 6974
rect 6310 6972 6316 6974
rect 6380 6972 6386 7036
rect 6729 7034 6795 7037
rect 7557 7034 7623 7037
rect 6729 7032 7623 7034
rect 6729 6976 6734 7032
rect 6790 6976 7562 7032
rect 7618 6976 7623 7032
rect 6729 6974 7623 6976
rect 6729 6971 6795 6974
rect 7557 6971 7623 6974
rect 8334 6972 8340 7036
rect 8404 7034 8410 7036
rect 9213 7034 9279 7037
rect 8404 7032 9279 7034
rect 8404 6976 9218 7032
rect 9274 6976 9279 7032
rect 8404 6974 9279 6976
rect 8404 6972 8410 6974
rect 9213 6971 9279 6974
rect 10685 7034 10751 7037
rect 11237 7034 11303 7037
rect 14089 7034 14155 7037
rect 10685 7032 14155 7034
rect 10685 6976 10690 7032
rect 10746 6976 11242 7032
rect 11298 6976 14094 7032
rect 14150 6976 14155 7032
rect 10685 6974 14155 6976
rect 10685 6971 10751 6974
rect 11237 6971 11303 6974
rect 14089 6971 14155 6974
rect 15929 7034 15995 7037
rect 19014 7036 19074 7110
rect 19149 7168 19380 7170
rect 19149 7112 19154 7168
rect 19210 7112 19380 7168
rect 19149 7110 19380 7112
rect 19149 7107 19215 7110
rect 19374 7108 19380 7110
rect 19444 7108 19450 7172
rect 19520 7170 19580 7243
rect 22320 7216 22800 7246
rect 19977 7170 20043 7173
rect 19520 7168 20043 7170
rect 19520 7112 19982 7168
rect 20038 7112 20043 7168
rect 19520 7110 20043 7112
rect 19977 7107 20043 7110
rect 15929 7032 18890 7034
rect 15929 6976 15934 7032
rect 15990 6976 18890 7032
rect 15929 6974 18890 6976
rect 15929 6971 15995 6974
rect 0 6838 2146 6898
rect 2221 6898 2287 6901
rect 8017 6898 8083 6901
rect 16849 6898 16915 6901
rect 2221 6896 7620 6898
rect 2221 6840 2226 6896
rect 2282 6840 7620 6896
rect 2221 6838 7620 6840
rect 0 6808 480 6838
rect 2221 6835 2287 6838
rect 3601 6762 3667 6765
rect 7560 6762 7620 6838
rect 8017 6896 16915 6898
rect 8017 6840 8022 6896
rect 8078 6840 16854 6896
rect 16910 6840 16915 6896
rect 8017 6838 16915 6840
rect 8017 6835 8083 6838
rect 16849 6835 16915 6838
rect 17217 6898 17283 6901
rect 17769 6898 17835 6901
rect 18597 6898 18663 6901
rect 18830 6900 18890 6974
rect 19006 6972 19012 7036
rect 19076 7034 19082 7036
rect 20989 7034 21055 7037
rect 19076 7032 21055 7034
rect 19076 6976 20994 7032
rect 21050 6976 21055 7032
rect 19076 6974 21055 6976
rect 19076 6972 19082 6974
rect 20989 6971 21055 6974
rect 17217 6896 17602 6898
rect 17217 6840 17222 6896
rect 17278 6840 17602 6896
rect 17217 6838 17602 6840
rect 17217 6835 17283 6838
rect 17401 6762 17467 6765
rect 3601 6760 7482 6762
rect 3601 6704 3606 6760
rect 3662 6704 7482 6760
rect 3601 6702 7482 6704
rect 7560 6760 17467 6762
rect 7560 6704 17406 6760
rect 17462 6704 17467 6760
rect 7560 6702 17467 6704
rect 17542 6762 17602 6838
rect 17769 6896 18663 6898
rect 17769 6840 17774 6896
rect 17830 6840 18602 6896
rect 18658 6840 18663 6896
rect 17769 6838 18663 6840
rect 17769 6835 17835 6838
rect 18597 6835 18663 6838
rect 18822 6836 18828 6900
rect 18892 6898 18898 6900
rect 19742 6898 19748 6900
rect 18892 6838 19748 6898
rect 18892 6836 18898 6838
rect 19742 6836 19748 6838
rect 19812 6836 19818 6900
rect 20069 6898 20135 6901
rect 22320 6898 22800 6928
rect 20069 6896 22800 6898
rect 20069 6840 20074 6896
rect 20130 6840 22800 6896
rect 20069 6838 22800 6840
rect 20069 6835 20135 6838
rect 22320 6808 22800 6838
rect 20161 6762 20227 6765
rect 17542 6760 20227 6762
rect 17542 6704 20166 6760
rect 20222 6704 20227 6760
rect 17542 6702 20227 6704
rect 3601 6699 3667 6702
rect 6453 6626 6519 6629
rect 7281 6626 7347 6629
rect 6453 6624 7347 6626
rect 6453 6568 6458 6624
rect 6514 6568 7286 6624
rect 7342 6568 7347 6624
rect 6453 6566 7347 6568
rect 7422 6626 7482 6702
rect 17401 6699 17467 6702
rect 20161 6699 20227 6702
rect 8017 6626 8083 6629
rect 7422 6624 8083 6626
rect 7422 6568 8022 6624
rect 8078 6568 8083 6624
rect 7422 6566 8083 6568
rect 6453 6563 6519 6566
rect 7281 6563 7347 6566
rect 8017 6563 8083 6566
rect 8661 6626 8727 6629
rect 10685 6626 10751 6629
rect 8661 6624 10751 6626
rect 8661 6568 8666 6624
rect 8722 6568 10690 6624
rect 10746 6568 10751 6624
rect 8661 6566 10751 6568
rect 8661 6563 8727 6566
rect 10685 6563 10751 6566
rect 11646 6564 11652 6628
rect 11716 6626 11722 6628
rect 11881 6626 11947 6629
rect 16941 6626 17007 6629
rect 11716 6624 17007 6626
rect 11716 6568 11886 6624
rect 11942 6568 16946 6624
rect 17002 6568 17007 6624
rect 11716 6566 17007 6568
rect 11716 6564 11722 6566
rect 11881 6563 11947 6566
rect 16941 6563 17007 6566
rect 18689 6626 18755 6629
rect 20713 6626 20779 6629
rect 18689 6624 20779 6626
rect 18689 6568 18694 6624
rect 18750 6568 20718 6624
rect 20774 6568 20779 6624
rect 18689 6566 20779 6568
rect 18689 6563 18755 6566
rect 20713 6563 20779 6566
rect 4376 6560 4696 6561
rect 0 6490 480 6520
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 2814 6490 2820 6492
rect 0 6430 2820 6490
rect 0 6400 480 6430
rect 2814 6428 2820 6430
rect 2884 6428 2890 6492
rect 6361 6490 6427 6493
rect 8334 6490 8340 6492
rect 6361 6488 8340 6490
rect 6361 6432 6366 6488
rect 6422 6432 8340 6488
rect 6361 6430 8340 6432
rect 6361 6427 6427 6430
rect 8334 6428 8340 6430
rect 8404 6428 8410 6492
rect 9121 6490 9187 6493
rect 9857 6492 9923 6493
rect 9438 6490 9444 6492
rect 9121 6488 9444 6490
rect 9121 6432 9126 6488
rect 9182 6432 9444 6488
rect 9121 6430 9444 6432
rect 9121 6427 9187 6430
rect 9438 6428 9444 6430
rect 9508 6428 9514 6492
rect 9806 6428 9812 6492
rect 9876 6490 9923 6492
rect 9876 6488 9968 6490
rect 9918 6432 9968 6488
rect 9876 6430 9968 6432
rect 9876 6428 9923 6430
rect 12382 6428 12388 6492
rect 12452 6490 12458 6492
rect 12525 6490 12591 6493
rect 12801 6492 12867 6493
rect 12750 6490 12756 6492
rect 12452 6488 12591 6490
rect 12452 6432 12530 6488
rect 12586 6432 12591 6488
rect 12452 6430 12591 6432
rect 12710 6430 12756 6490
rect 12820 6488 12867 6492
rect 12862 6432 12867 6488
rect 12452 6428 12458 6430
rect 9857 6427 9923 6428
rect 12525 6427 12591 6430
rect 12750 6428 12756 6430
rect 12820 6428 12867 6432
rect 13118 6428 13124 6492
rect 13188 6490 13194 6492
rect 13670 6490 13676 6492
rect 13188 6430 13676 6490
rect 13188 6428 13194 6430
rect 13670 6428 13676 6430
rect 13740 6428 13746 6492
rect 17166 6428 17172 6492
rect 17236 6490 17242 6492
rect 17677 6490 17743 6493
rect 17236 6488 17743 6490
rect 17236 6432 17682 6488
rect 17738 6432 17743 6488
rect 17236 6430 17743 6432
rect 17236 6428 17242 6430
rect 12801 6427 12867 6428
rect 17677 6427 17743 6430
rect 20529 6490 20595 6493
rect 22320 6490 22800 6520
rect 20529 6488 22800 6490
rect 20529 6432 20534 6488
rect 20590 6432 22800 6488
rect 20529 6430 22800 6432
rect 20529 6427 20595 6430
rect 22320 6400 22800 6430
rect 3366 6292 3372 6356
rect 3436 6354 3442 6356
rect 4613 6354 4679 6357
rect 3436 6352 4679 6354
rect 3436 6296 4618 6352
rect 4674 6296 4679 6352
rect 3436 6294 4679 6296
rect 3436 6292 3442 6294
rect 4613 6291 4679 6294
rect 4889 6354 4955 6357
rect 16430 6354 16436 6356
rect 4889 6352 16436 6354
rect 4889 6296 4894 6352
rect 4950 6296 16436 6352
rect 4889 6294 16436 6296
rect 4889 6291 4955 6294
rect 16430 6292 16436 6294
rect 16500 6292 16506 6356
rect 18413 6354 18479 6357
rect 19006 6354 19012 6356
rect 18413 6352 19012 6354
rect 18413 6296 18418 6352
rect 18474 6296 19012 6352
rect 18413 6294 19012 6296
rect 18413 6291 18479 6294
rect 19006 6292 19012 6294
rect 19076 6292 19082 6356
rect 3325 6218 3391 6221
rect 9765 6218 9831 6221
rect 18965 6220 19031 6221
rect 18965 6218 19012 6220
rect 3325 6216 9831 6218
rect 3325 6160 3330 6216
rect 3386 6160 9770 6216
rect 9826 6160 9831 6216
rect 3325 6158 9831 6160
rect 3325 6155 3391 6158
rect 9765 6155 9831 6158
rect 9998 6158 15762 6218
rect 18920 6216 19012 6218
rect 18920 6160 18970 6216
rect 18920 6158 19012 6160
rect 0 6082 480 6112
rect 5257 6082 5323 6085
rect 7097 6084 7163 6085
rect 7046 6082 7052 6084
rect 0 6080 5323 6082
rect 0 6024 5262 6080
rect 5318 6024 5323 6080
rect 0 6022 5323 6024
rect 7006 6022 7052 6082
rect 7116 6080 7163 6084
rect 7158 6024 7163 6080
rect 0 5992 480 6022
rect 5257 6019 5323 6022
rect 7046 6020 7052 6022
rect 7116 6020 7163 6024
rect 7097 6019 7163 6020
rect 8293 6082 8359 6085
rect 9998 6082 10058 6158
rect 8293 6080 10058 6082
rect 8293 6024 8298 6080
rect 8354 6024 10058 6080
rect 8293 6022 10058 6024
rect 10685 6082 10751 6085
rect 13169 6082 13235 6085
rect 10685 6080 13235 6082
rect 10685 6024 10690 6080
rect 10746 6024 13174 6080
rect 13230 6024 13235 6080
rect 10685 6022 13235 6024
rect 15702 6082 15762 6158
rect 18965 6156 19012 6158
rect 19076 6156 19082 6220
rect 18965 6155 19031 6156
rect 22320 6082 22800 6112
rect 15702 6022 22800 6082
rect 8293 6019 8359 6022
rect 10685 6019 10751 6022
rect 13169 6019 13235 6022
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 22320 5992 22800 6022
rect 14672 5951 14992 5952
rect 7046 5884 7052 5948
rect 7116 5946 7122 5948
rect 7281 5946 7347 5949
rect 7116 5944 7347 5946
rect 7116 5888 7286 5944
rect 7342 5888 7347 5944
rect 7116 5886 7347 5888
rect 7116 5884 7122 5886
rect 7281 5883 7347 5886
rect 8753 5946 8819 5949
rect 14365 5946 14431 5949
rect 8753 5944 14431 5946
rect 8753 5888 8758 5944
rect 8814 5888 14370 5944
rect 14426 5888 14431 5944
rect 8753 5886 14431 5888
rect 8753 5883 8819 5886
rect 14365 5883 14431 5886
rect 17718 5884 17724 5948
rect 17788 5946 17794 5948
rect 18965 5946 19031 5949
rect 17788 5944 19031 5946
rect 17788 5888 18970 5944
rect 19026 5888 19031 5944
rect 17788 5886 19031 5888
rect 17788 5884 17794 5886
rect 18965 5883 19031 5886
rect 6913 5810 6979 5813
rect 8937 5812 9003 5813
rect 8886 5810 8892 5812
rect 6913 5808 7850 5810
rect 6913 5752 6918 5808
rect 6974 5752 7850 5808
rect 6913 5750 7850 5752
rect 8846 5750 8892 5810
rect 8956 5808 9003 5812
rect 9397 5812 9463 5813
rect 9397 5810 9444 5812
rect 8998 5752 9003 5808
rect 6913 5747 6979 5750
rect 0 5674 480 5704
rect 4061 5674 4127 5677
rect 0 5672 4127 5674
rect 0 5616 4066 5672
rect 4122 5616 4127 5672
rect 0 5614 4127 5616
rect 0 5584 480 5614
rect 4061 5611 4127 5614
rect 5206 5612 5212 5676
rect 5276 5674 5282 5676
rect 7465 5674 7531 5677
rect 7598 5674 7604 5676
rect 5276 5614 7298 5674
rect 5276 5612 5282 5614
rect 7238 5538 7298 5614
rect 7465 5672 7604 5674
rect 7465 5616 7470 5672
rect 7526 5616 7604 5672
rect 7465 5614 7604 5616
rect 7465 5611 7531 5614
rect 7598 5612 7604 5614
rect 7668 5612 7674 5676
rect 7790 5674 7850 5750
rect 8886 5748 8892 5750
rect 8956 5748 9003 5752
rect 9352 5808 9444 5810
rect 9352 5752 9402 5808
rect 9352 5750 9444 5752
rect 8937 5747 9003 5748
rect 9397 5748 9444 5750
rect 9508 5748 9514 5812
rect 10542 5748 10548 5812
rect 10612 5810 10618 5812
rect 14457 5810 14523 5813
rect 18689 5810 18755 5813
rect 10612 5750 13922 5810
rect 10612 5748 10618 5750
rect 9397 5747 9463 5748
rect 13721 5674 13787 5677
rect 7790 5672 13787 5674
rect 7790 5616 13726 5672
rect 13782 5616 13787 5672
rect 7790 5614 13787 5616
rect 13862 5674 13922 5750
rect 14457 5808 18755 5810
rect 14457 5752 14462 5808
rect 14518 5752 18694 5808
rect 18750 5752 18755 5808
rect 14457 5750 18755 5752
rect 14457 5747 14523 5750
rect 18689 5747 18755 5750
rect 14641 5674 14707 5677
rect 13862 5672 14707 5674
rect 13862 5616 14646 5672
rect 14702 5616 14707 5672
rect 13862 5614 14707 5616
rect 13721 5611 13787 5614
rect 14641 5611 14707 5614
rect 17953 5674 18019 5677
rect 22320 5674 22800 5704
rect 17953 5672 22800 5674
rect 17953 5616 17958 5672
rect 18014 5616 22800 5672
rect 17953 5614 22800 5616
rect 17953 5611 18019 5614
rect 22320 5584 22800 5614
rect 10685 5538 10751 5541
rect 11697 5540 11763 5541
rect 7238 5536 10751 5538
rect 7238 5480 10690 5536
rect 10746 5480 10751 5536
rect 7238 5478 10751 5480
rect 10685 5475 10751 5478
rect 11646 5476 11652 5540
rect 11716 5538 11763 5540
rect 15837 5538 15903 5541
rect 11716 5536 15903 5538
rect 11758 5480 15842 5536
rect 15898 5480 15903 5536
rect 11716 5478 15903 5480
rect 11716 5476 11763 5478
rect 11697 5475 11763 5476
rect 15837 5475 15903 5478
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 6177 5402 6243 5405
rect 10869 5402 10935 5405
rect 6177 5400 10935 5402
rect 6177 5344 6182 5400
rect 6238 5344 10874 5400
rect 10930 5344 10935 5400
rect 6177 5342 10935 5344
rect 6177 5339 6243 5342
rect 10869 5339 10935 5342
rect 12433 5402 12499 5405
rect 17953 5402 18019 5405
rect 12433 5400 18019 5402
rect 12433 5344 12438 5400
rect 12494 5344 17958 5400
rect 18014 5344 18019 5400
rect 12433 5342 18019 5344
rect 12433 5339 12499 5342
rect 17953 5339 18019 5342
rect 19742 5340 19748 5404
rect 19812 5402 19818 5404
rect 19885 5402 19951 5405
rect 19812 5400 19951 5402
rect 19812 5344 19890 5400
rect 19946 5344 19951 5400
rect 19812 5342 19951 5344
rect 19812 5340 19818 5342
rect 19885 5339 19951 5342
rect 0 5266 480 5296
rect 6729 5266 6795 5269
rect 0 5264 6795 5266
rect 0 5208 6734 5264
rect 6790 5208 6795 5264
rect 0 5206 6795 5208
rect 0 5176 480 5206
rect 6729 5203 6795 5206
rect 7097 5266 7163 5269
rect 7097 5264 12450 5266
rect 7097 5208 7102 5264
rect 7158 5208 12450 5264
rect 7097 5206 12450 5208
rect 7097 5203 7163 5206
rect 4838 5068 4844 5132
rect 4908 5130 4914 5132
rect 10133 5130 10199 5133
rect 4908 5128 10199 5130
rect 4908 5072 10138 5128
rect 10194 5072 10199 5128
rect 4908 5070 10199 5072
rect 4908 5068 4914 5070
rect 10133 5067 10199 5070
rect 10317 5130 10383 5133
rect 12249 5130 12315 5133
rect 10317 5128 12315 5130
rect 10317 5072 10322 5128
rect 10378 5072 12254 5128
rect 12310 5072 12315 5128
rect 10317 5070 12315 5072
rect 12390 5130 12450 5206
rect 14222 5204 14228 5268
rect 14292 5266 14298 5268
rect 17493 5266 17559 5269
rect 14292 5264 17559 5266
rect 14292 5208 17498 5264
rect 17554 5208 17559 5264
rect 14292 5206 17559 5208
rect 14292 5204 14298 5206
rect 17493 5203 17559 5206
rect 17953 5266 18019 5269
rect 22320 5266 22800 5296
rect 17953 5264 22800 5266
rect 17953 5208 17958 5264
rect 18014 5208 22800 5264
rect 17953 5206 22800 5208
rect 17953 5203 18019 5206
rect 22320 5176 22800 5206
rect 14549 5130 14615 5133
rect 12390 5128 14615 5130
rect 12390 5072 14554 5128
rect 14610 5072 14615 5128
rect 12390 5070 14615 5072
rect 10317 5067 10383 5070
rect 12249 5067 12315 5070
rect 14549 5067 14615 5070
rect 3969 4994 4035 4997
rect 7557 4994 7623 4997
rect 12893 4994 12959 4997
rect 3969 4992 7623 4994
rect 3969 4936 3974 4992
rect 4030 4936 7562 4992
rect 7618 4936 7623 4992
rect 3969 4934 7623 4936
rect 3969 4931 4035 4934
rect 7557 4931 7623 4934
rect 8204 4992 12959 4994
rect 8204 4936 12898 4992
rect 12954 4936 12959 4992
rect 8204 4934 12959 4936
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 5533 4858 5599 4861
rect 0 4856 5599 4858
rect 0 4800 5538 4856
rect 5594 4800 5599 4856
rect 0 4798 5599 4800
rect 0 4768 480 4798
rect 5533 4795 5599 4798
rect 8204 4722 8264 4934
rect 12893 4931 12959 4934
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 8477 4858 8543 4861
rect 9213 4858 9279 4861
rect 9489 4860 9555 4861
rect 8477 4856 9279 4858
rect 8477 4800 8482 4856
rect 8538 4800 9218 4856
rect 9274 4800 9279 4856
rect 8477 4798 9279 4800
rect 8477 4795 8543 4798
rect 9213 4795 9279 4798
rect 9438 4796 9444 4860
rect 9508 4858 9555 4860
rect 11513 4858 11579 4861
rect 14365 4858 14431 4861
rect 9508 4856 9600 4858
rect 9550 4800 9600 4856
rect 9508 4798 9600 4800
rect 11513 4856 14431 4858
rect 11513 4800 11518 4856
rect 11574 4800 14370 4856
rect 14426 4800 14431 4856
rect 11513 4798 14431 4800
rect 9508 4796 9555 4798
rect 9489 4795 9555 4796
rect 11513 4795 11579 4798
rect 14365 4795 14431 4798
rect 15837 4858 15903 4861
rect 22320 4858 22800 4888
rect 15837 4856 22800 4858
rect 15837 4800 15842 4856
rect 15898 4800 22800 4856
rect 15837 4798 22800 4800
rect 15837 4795 15903 4798
rect 22320 4768 22800 4798
rect 13353 4722 13419 4725
rect 15009 4722 15075 4725
rect 4248 4662 8264 4722
rect 9446 4720 15075 4722
rect 9446 4664 13358 4720
rect 13414 4664 15014 4720
rect 15070 4664 15075 4720
rect 9446 4662 15075 4664
rect 0 4450 480 4480
rect 4248 4450 4308 4662
rect 7281 4586 7347 4589
rect 9254 4586 9260 4588
rect 7281 4584 9260 4586
rect 7281 4528 7286 4584
rect 7342 4528 9260 4584
rect 7281 4526 9260 4528
rect 7281 4523 7347 4526
rect 9254 4524 9260 4526
rect 9324 4524 9330 4588
rect 0 4390 4308 4450
rect 6269 4450 6335 4453
rect 9446 4450 9506 4662
rect 13353 4659 13419 4662
rect 15009 4659 15075 4662
rect 15377 4722 15443 4725
rect 16021 4722 16087 4725
rect 15377 4720 16087 4722
rect 15377 4664 15382 4720
rect 15438 4664 16026 4720
rect 16082 4664 16087 4720
rect 15377 4662 16087 4664
rect 15377 4659 15443 4662
rect 16021 4659 16087 4662
rect 10041 4586 10107 4589
rect 10317 4586 10383 4589
rect 17401 4586 17467 4589
rect 19198 4586 19396 4620
rect 10041 4584 17467 4586
rect 10041 4528 10046 4584
rect 10102 4528 10322 4584
rect 10378 4528 17406 4584
rect 17462 4528 17467 4584
rect 10041 4526 17467 4528
rect 10041 4523 10107 4526
rect 10317 4523 10383 4526
rect 17401 4523 17467 4526
rect 17542 4560 19994 4586
rect 17542 4526 19258 4560
rect 19336 4526 19994 4560
rect 6269 4448 9506 4450
rect 6269 4392 6274 4448
rect 6330 4392 9506 4448
rect 6269 4390 9506 4392
rect 0 4360 480 4390
rect 6269 4387 6335 4390
rect 12934 4388 12940 4452
rect 13004 4450 13010 4452
rect 17542 4450 17602 4526
rect 13004 4390 17602 4450
rect 19934 4450 19994 4526
rect 22320 4450 22800 4480
rect 19934 4390 22800 4450
rect 13004 4388 13010 4390
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 22320 4360 22800 4390
rect 18104 4319 18424 4320
rect 6862 4252 6868 4316
rect 6932 4314 6938 4316
rect 8017 4314 8083 4317
rect 8886 4314 8892 4316
rect 6932 4312 8892 4314
rect 6932 4256 8022 4312
rect 8078 4256 8892 4312
rect 6932 4254 8892 4256
rect 6932 4252 6938 4254
rect 8017 4251 8083 4254
rect 8886 4252 8892 4254
rect 8956 4252 8962 4316
rect 9121 4314 9187 4317
rect 10685 4314 10751 4317
rect 9121 4312 10751 4314
rect 9121 4256 9126 4312
rect 9182 4256 10690 4312
rect 10746 4256 10751 4312
rect 9121 4254 10751 4256
rect 9121 4251 9187 4254
rect 10685 4251 10751 4254
rect 12525 4314 12591 4317
rect 12750 4314 12756 4316
rect 12525 4312 12756 4314
rect 12525 4256 12530 4312
rect 12586 4256 12756 4312
rect 12525 4254 12756 4256
rect 12525 4251 12591 4254
rect 12750 4252 12756 4254
rect 12820 4252 12826 4316
rect 3141 4180 3207 4181
rect 3141 4176 3188 4180
rect 3252 4178 3258 4180
rect 5257 4178 5323 4181
rect 5390 4178 5396 4180
rect 3141 4120 3146 4176
rect 3141 4116 3188 4120
rect 3252 4118 3298 4178
rect 5257 4176 5396 4178
rect 5257 4120 5262 4176
rect 5318 4120 5396 4176
rect 5257 4118 5396 4120
rect 3252 4116 3258 4118
rect 3141 4115 3207 4116
rect 5257 4115 5323 4118
rect 5390 4116 5396 4118
rect 5460 4116 5466 4180
rect 5533 4178 5599 4181
rect 13629 4178 13695 4181
rect 19149 4178 19215 4181
rect 5533 4176 19215 4178
rect 5533 4120 5538 4176
rect 5594 4120 13634 4176
rect 13690 4120 19154 4176
rect 19210 4120 19215 4176
rect 5533 4118 19215 4120
rect 5533 4115 5599 4118
rect 0 4042 480 4072
rect 4061 4042 4127 4045
rect 0 4040 4127 4042
rect 0 3984 4066 4040
rect 4122 3984 4127 4040
rect 0 3982 4127 3984
rect 0 3952 480 3982
rect 4061 3979 4127 3982
rect 4429 4042 4495 4045
rect 5206 4042 5212 4044
rect 4429 4040 5212 4042
rect 4429 3984 4434 4040
rect 4490 3984 5212 4040
rect 4429 3982 5212 3984
rect 4429 3979 4495 3982
rect 5206 3980 5212 3982
rect 5276 3980 5282 4044
rect 6637 4042 6703 4045
rect 7414 4042 7420 4044
rect 6637 4040 7420 4042
rect 6637 3984 6642 4040
rect 6698 3984 7420 4040
rect 6637 3982 7420 3984
rect 6637 3979 6703 3982
rect 7414 3980 7420 3982
rect 7484 4042 7490 4044
rect 11973 4042 12039 4045
rect 12574 4044 12634 4118
rect 13629 4115 13695 4118
rect 19149 4115 19215 4118
rect 7484 4040 12039 4042
rect 7484 3984 11978 4040
rect 12034 3984 12039 4040
rect 7484 3982 12039 3984
rect 7484 3980 7490 3982
rect 11973 3979 12039 3982
rect 12566 3980 12572 4044
rect 12636 3980 12642 4044
rect 18638 3980 18644 4044
rect 18708 4042 18714 4044
rect 18873 4042 18939 4045
rect 22320 4042 22800 4072
rect 18708 4040 18939 4042
rect 18708 3984 18878 4040
rect 18934 3984 18939 4040
rect 19336 4008 22800 4042
rect 18708 3982 18939 3984
rect 18708 3980 18714 3982
rect 18873 3979 18939 3982
rect 19244 3982 22800 4008
rect 19244 3948 19396 3982
rect 22320 3952 22800 3982
rect 2405 3906 2471 3909
rect 7557 3906 7623 3909
rect 2405 3904 7623 3906
rect 2405 3848 2410 3904
rect 2466 3848 7562 3904
rect 7618 3848 7623 3904
rect 2405 3846 7623 3848
rect 2405 3843 2471 3846
rect 7557 3843 7623 3846
rect 8661 3906 8727 3909
rect 9070 3906 9076 3908
rect 8661 3904 9076 3906
rect 8661 3848 8666 3904
rect 8722 3848 9076 3904
rect 8661 3846 9076 3848
rect 8661 3843 8727 3846
rect 9070 3844 9076 3846
rect 9140 3844 9146 3908
rect 9305 3906 9371 3909
rect 12525 3906 12591 3909
rect 9305 3904 12591 3906
rect 9305 3848 9310 3904
rect 9366 3848 12530 3904
rect 12586 3848 12591 3904
rect 9305 3846 12591 3848
rect 9305 3843 9371 3846
rect 12525 3843 12591 3846
rect 13905 3906 13971 3909
rect 14038 3906 14044 3908
rect 13905 3904 14044 3906
rect 13905 3848 13910 3904
rect 13966 3848 14044 3904
rect 13905 3846 14044 3848
rect 13905 3843 13971 3846
rect 14038 3844 14044 3846
rect 14108 3844 14114 3908
rect 16614 3844 16620 3908
rect 16684 3906 16690 3908
rect 19244 3906 19304 3948
rect 16684 3846 19304 3906
rect 16684 3844 16690 3846
rect 7808 3840 8128 3841
rect 0 3770 480 3800
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 3182 3770 3188 3772
rect 0 3710 3188 3770
rect 0 3680 480 3710
rect 3182 3708 3188 3710
rect 3252 3708 3258 3772
rect 3918 3708 3924 3772
rect 3988 3770 3994 3772
rect 4245 3770 4311 3773
rect 14273 3770 14339 3773
rect 3988 3768 4311 3770
rect 3988 3712 4250 3768
rect 4306 3712 4311 3768
rect 3988 3710 4311 3712
rect 3988 3708 3994 3710
rect 4245 3707 4311 3710
rect 8204 3768 14339 3770
rect 8204 3712 14278 3768
rect 14334 3712 14339 3768
rect 8204 3710 14339 3712
rect 5533 3634 5599 3637
rect 8204 3634 8264 3710
rect 14273 3707 14339 3710
rect 20713 3770 20779 3773
rect 22320 3770 22800 3800
rect 20713 3768 22800 3770
rect 20713 3712 20718 3768
rect 20774 3712 22800 3768
rect 20713 3710 22800 3712
rect 20713 3707 20779 3710
rect 22320 3680 22800 3710
rect 5533 3632 8264 3634
rect 5533 3576 5538 3632
rect 5594 3576 8264 3632
rect 5533 3574 8264 3576
rect 8937 3634 9003 3637
rect 13997 3634 14063 3637
rect 8937 3632 14063 3634
rect 8937 3576 8942 3632
rect 8998 3576 14002 3632
rect 14058 3576 14063 3632
rect 8937 3574 14063 3576
rect 5533 3571 5599 3574
rect 8937 3571 9003 3574
rect 13997 3571 14063 3574
rect 2865 3498 2931 3501
rect 8109 3498 8175 3501
rect 8937 3498 9003 3501
rect 2865 3496 9003 3498
rect 2865 3440 2870 3496
rect 2926 3440 8114 3496
rect 8170 3440 8942 3496
rect 8998 3440 9003 3496
rect 2865 3438 9003 3440
rect 2865 3435 2931 3438
rect 8109 3435 8175 3438
rect 8937 3435 9003 3438
rect 9070 3436 9076 3500
rect 9140 3498 9146 3500
rect 10133 3498 10199 3501
rect 13537 3498 13603 3501
rect 9140 3496 13603 3498
rect 9140 3440 10138 3496
rect 10194 3440 13542 3496
rect 13598 3440 13603 3496
rect 9140 3438 13603 3440
rect 9140 3436 9146 3438
rect 10133 3435 10199 3438
rect 13537 3435 13603 3438
rect 13905 3498 13971 3501
rect 20713 3498 20779 3501
rect 13905 3496 20779 3498
rect 13905 3440 13910 3496
rect 13966 3440 20718 3496
rect 20774 3440 20779 3496
rect 13905 3438 20779 3440
rect 13905 3435 13971 3438
rect 20713 3435 20779 3438
rect 0 3362 480 3392
rect 2405 3362 2471 3365
rect 0 3360 2471 3362
rect 0 3304 2410 3360
rect 2466 3304 2471 3360
rect 0 3302 2471 3304
rect 0 3272 480 3302
rect 2405 3299 2471 3302
rect 6821 3362 6887 3365
rect 9622 3362 9628 3364
rect 6821 3360 9628 3362
rect 6821 3304 6826 3360
rect 6882 3304 9628 3360
rect 6821 3302 9628 3304
rect 6821 3299 6887 3302
rect 9622 3300 9628 3302
rect 9692 3362 9698 3364
rect 10501 3362 10567 3365
rect 9692 3360 10567 3362
rect 9692 3304 10506 3360
rect 10562 3304 10567 3360
rect 9692 3302 10567 3304
rect 9692 3300 9698 3302
rect 10501 3299 10567 3302
rect 14457 3362 14523 3365
rect 17166 3362 17172 3364
rect 14457 3360 17172 3362
rect 14457 3304 14462 3360
rect 14518 3304 17172 3360
rect 14457 3302 17172 3304
rect 14457 3299 14523 3302
rect 17166 3300 17172 3302
rect 17236 3300 17242 3364
rect 21909 3362 21975 3365
rect 22320 3362 22800 3392
rect 21909 3360 22800 3362
rect 21909 3304 21914 3360
rect 21970 3304 22800 3360
rect 21909 3302 22800 3304
rect 21909 3299 21975 3302
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 22320 3272 22800 3302
rect 18104 3231 18424 3232
rect 7598 3164 7604 3228
rect 7668 3226 7674 3228
rect 7741 3226 7807 3229
rect 7668 3224 7807 3226
rect 7668 3168 7746 3224
rect 7802 3168 7807 3224
rect 7668 3166 7807 3168
rect 7668 3164 7674 3166
rect 7741 3163 7807 3166
rect 8702 3164 8708 3228
rect 8772 3226 8778 3228
rect 15837 3226 15903 3229
rect 8772 3166 11162 3226
rect 8772 3164 8778 3166
rect 6821 3090 6887 3093
rect 8477 3090 8543 3093
rect 6821 3088 8543 3090
rect 6821 3032 6826 3088
rect 6882 3032 8482 3088
rect 8538 3032 8543 3088
rect 6821 3030 8543 3032
rect 6821 3027 6887 3030
rect 8477 3027 8543 3030
rect 9029 3090 9095 3093
rect 10133 3090 10199 3093
rect 10961 3090 11027 3093
rect 9029 3088 11027 3090
rect 9029 3032 9034 3088
rect 9090 3032 10138 3088
rect 10194 3032 10966 3088
rect 11022 3032 11027 3088
rect 9029 3030 11027 3032
rect 11102 3090 11162 3166
rect 11654 3224 15903 3226
rect 11654 3168 15842 3224
rect 15898 3168 15903 3224
rect 11654 3166 15903 3168
rect 11654 3090 11714 3166
rect 15837 3163 15903 3166
rect 17401 3226 17467 3229
rect 17534 3226 17540 3228
rect 17401 3224 17540 3226
rect 17401 3168 17406 3224
rect 17462 3168 17540 3224
rect 17401 3166 17540 3168
rect 17401 3163 17467 3166
rect 17534 3164 17540 3166
rect 17604 3164 17610 3228
rect 18689 3226 18755 3229
rect 19006 3226 19012 3228
rect 18689 3224 19012 3226
rect 18689 3168 18694 3224
rect 18750 3168 19012 3224
rect 18689 3166 19012 3168
rect 18689 3163 18755 3166
rect 19006 3164 19012 3166
rect 19076 3164 19082 3228
rect 19333 3226 19399 3229
rect 20805 3226 20871 3229
rect 19333 3224 20871 3226
rect 19333 3168 19338 3224
rect 19394 3168 20810 3224
rect 20866 3168 20871 3224
rect 19333 3166 20871 3168
rect 19333 3163 19399 3166
rect 20805 3163 20871 3166
rect 13077 3090 13143 3093
rect 11102 3030 11714 3090
rect 11792 3088 13143 3090
rect 11792 3032 13082 3088
rect 13138 3032 13143 3088
rect 11792 3030 13143 3032
rect 9029 3027 9095 3030
rect 10133 3027 10199 3030
rect 10961 3027 11027 3030
rect 0 2954 480 2984
rect 3233 2954 3299 2957
rect 0 2952 3299 2954
rect 0 2896 3238 2952
rect 3294 2896 3299 2952
rect 0 2894 3299 2896
rect 0 2864 480 2894
rect 3233 2891 3299 2894
rect 3877 2954 3943 2957
rect 7230 2954 7236 2956
rect 3877 2952 7236 2954
rect 3877 2896 3882 2952
rect 3938 2896 7236 2952
rect 3877 2894 7236 2896
rect 3877 2891 3943 2894
rect 7230 2892 7236 2894
rect 7300 2892 7306 2956
rect 8477 2954 8543 2957
rect 11646 2954 11652 2956
rect 7422 2894 8402 2954
rect 5717 2818 5783 2821
rect 6453 2818 6519 2821
rect 7422 2818 7482 2894
rect 5717 2816 7482 2818
rect 5717 2760 5722 2816
rect 5778 2760 6458 2816
rect 6514 2760 7482 2816
rect 5717 2758 7482 2760
rect 8342 2818 8402 2894
rect 8477 2952 11652 2954
rect 8477 2896 8482 2952
rect 8538 2896 11652 2952
rect 8477 2894 11652 2896
rect 8477 2891 8543 2894
rect 11646 2892 11652 2894
rect 11716 2892 11722 2956
rect 11792 2818 11852 3030
rect 13077 3027 13143 3030
rect 12341 2954 12407 2957
rect 20437 2954 20503 2957
rect 22320 2954 22800 2984
rect 12341 2952 20503 2954
rect 12341 2896 12346 2952
rect 12402 2896 20442 2952
rect 20498 2896 20503 2952
rect 12341 2894 20503 2896
rect 12341 2891 12407 2894
rect 20437 2891 20503 2894
rect 20670 2894 22800 2954
rect 8342 2758 11852 2818
rect 5717 2755 5783 2758
rect 6453 2755 6519 2758
rect 12382 2756 12388 2820
rect 12452 2818 12458 2820
rect 13997 2818 14063 2821
rect 12452 2816 14063 2818
rect 12452 2760 14002 2816
rect 14058 2760 14063 2816
rect 12452 2758 14063 2760
rect 12452 2756 12458 2758
rect 13997 2755 14063 2758
rect 17493 2818 17559 2821
rect 18965 2818 19031 2821
rect 17493 2816 19031 2818
rect 17493 2760 17498 2816
rect 17554 2760 18970 2816
rect 19026 2760 19031 2816
rect 17493 2758 19031 2760
rect 17493 2755 17559 2758
rect 18965 2755 19031 2758
rect 19149 2820 19215 2821
rect 19149 2816 19196 2820
rect 19260 2818 19266 2820
rect 20670 2818 20730 2894
rect 22320 2864 22800 2894
rect 19149 2760 19154 2816
rect 19149 2756 19196 2760
rect 19260 2758 20730 2818
rect 19260 2756 19266 2758
rect 19149 2755 19215 2756
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 2773 2682 2839 2685
rect 3601 2682 3667 2685
rect 2773 2680 3667 2682
rect 2773 2624 2778 2680
rect 2834 2624 3606 2680
rect 3662 2624 3667 2680
rect 2773 2622 3667 2624
rect 2773 2619 2839 2622
rect 3601 2619 3667 2622
rect 8334 2620 8340 2684
rect 8404 2682 8410 2684
rect 9121 2682 9187 2685
rect 8404 2680 9187 2682
rect 8404 2624 9126 2680
rect 9182 2624 9187 2680
rect 8404 2622 9187 2624
rect 8404 2620 8410 2622
rect 9121 2619 9187 2622
rect 16297 2682 16363 2685
rect 17902 2682 17908 2684
rect 16297 2680 17908 2682
rect 16297 2624 16302 2680
rect 16358 2624 17908 2680
rect 16297 2622 17908 2624
rect 16297 2619 16363 2622
rect 17902 2620 17908 2622
rect 17972 2620 17978 2684
rect 0 2546 480 2576
rect 2037 2546 2103 2549
rect 0 2544 2103 2546
rect 0 2488 2042 2544
rect 2098 2488 2103 2544
rect 0 2486 2103 2488
rect 0 2456 480 2486
rect 2037 2483 2103 2486
rect 8017 2546 8083 2549
rect 8702 2546 8708 2548
rect 8017 2544 8708 2546
rect 8017 2488 8022 2544
rect 8078 2488 8708 2544
rect 8017 2486 8708 2488
rect 8017 2483 8083 2486
rect 8702 2484 8708 2486
rect 8772 2484 8778 2548
rect 8937 2546 9003 2549
rect 11145 2546 11211 2549
rect 8937 2544 11211 2546
rect 8937 2488 8942 2544
rect 8998 2488 11150 2544
rect 11206 2488 11211 2544
rect 8937 2486 11211 2488
rect 8937 2483 9003 2486
rect 11145 2483 11211 2486
rect 11329 2546 11395 2549
rect 17585 2546 17651 2549
rect 11329 2544 17651 2546
rect 11329 2488 11334 2544
rect 11390 2488 17590 2544
rect 17646 2488 17651 2544
rect 11329 2486 17651 2488
rect 11329 2483 11395 2486
rect 17585 2483 17651 2486
rect 18781 2548 18847 2549
rect 18781 2544 18828 2548
rect 18892 2546 18898 2548
rect 20989 2546 21055 2549
rect 22320 2546 22800 2576
rect 18781 2488 18786 2544
rect 18781 2484 18828 2488
rect 18892 2486 18938 2546
rect 20989 2544 22800 2546
rect 20989 2488 20994 2544
rect 21050 2488 22800 2544
rect 20989 2486 22800 2488
rect 18892 2484 18898 2486
rect 18781 2483 18847 2484
rect 20989 2483 21055 2486
rect 22320 2456 22800 2486
rect 7189 2410 7255 2413
rect 9438 2410 9444 2412
rect 7189 2408 9444 2410
rect 7189 2352 7194 2408
rect 7250 2352 9444 2408
rect 7189 2350 9444 2352
rect 7189 2347 7255 2350
rect 9438 2348 9444 2350
rect 9508 2348 9514 2412
rect 17217 2410 17283 2413
rect 19558 2410 19564 2412
rect 17217 2408 19564 2410
rect 17217 2352 17222 2408
rect 17278 2352 19564 2408
rect 17217 2350 19564 2352
rect 17217 2347 17283 2350
rect 19558 2348 19564 2350
rect 19628 2348 19634 2412
rect 6678 2212 6684 2276
rect 6748 2274 6754 2276
rect 8753 2274 8819 2277
rect 6748 2272 8819 2274
rect 6748 2216 8758 2272
rect 8814 2216 8819 2272
rect 6748 2214 8819 2216
rect 6748 2212 6754 2214
rect 8753 2211 8819 2214
rect 18965 2274 19031 2277
rect 19742 2274 19748 2276
rect 18965 2272 19748 2274
rect 18965 2216 18970 2272
rect 19026 2216 19748 2272
rect 18965 2214 19748 2216
rect 18965 2211 19031 2214
rect 19742 2212 19748 2214
rect 19812 2212 19818 2276
rect 4376 2208 4696 2209
rect 0 2138 480 2168
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 3693 2138 3759 2141
rect 0 2136 3759 2138
rect 0 2080 3698 2136
rect 3754 2080 3759 2136
rect 0 2078 3759 2080
rect 0 2048 480 2078
rect 3693 2075 3759 2078
rect 7046 2076 7052 2140
rect 7116 2138 7122 2140
rect 8937 2138 9003 2141
rect 7116 2136 9003 2138
rect 7116 2080 8942 2136
rect 8998 2080 9003 2136
rect 7116 2078 9003 2080
rect 7116 2076 7122 2078
rect 8937 2075 9003 2078
rect 18597 2138 18663 2141
rect 22320 2138 22800 2168
rect 18597 2136 22800 2138
rect 18597 2080 18602 2136
rect 18658 2080 22800 2136
rect 18597 2078 22800 2080
rect 18597 2075 18663 2078
rect 22320 2048 22800 2078
rect 17033 2002 17099 2005
rect 19241 2002 19307 2005
rect 17033 2000 19307 2002
rect 17033 1944 17038 2000
rect 17094 1944 19246 2000
rect 19302 1944 19307 2000
rect 17033 1942 19307 1944
rect 17033 1939 17099 1942
rect 19241 1939 19307 1942
rect 0 1730 480 1760
rect 2773 1730 2839 1733
rect 0 1728 2839 1730
rect 0 1672 2778 1728
rect 2834 1672 2839 1728
rect 0 1670 2839 1672
rect 0 1640 480 1670
rect 2773 1667 2839 1670
rect 21173 1730 21239 1733
rect 22320 1730 22800 1760
rect 21173 1728 22800 1730
rect 21173 1672 21178 1728
rect 21234 1672 22800 1728
rect 21173 1670 22800 1672
rect 21173 1667 21239 1670
rect 22320 1640 22800 1670
rect 0 1322 480 1352
rect 3969 1322 4035 1325
rect 0 1320 4035 1322
rect 0 1264 3974 1320
rect 4030 1264 4035 1320
rect 0 1262 4035 1264
rect 0 1232 480 1262
rect 3969 1259 4035 1262
rect 18689 1322 18755 1325
rect 22320 1322 22800 1352
rect 18689 1320 22800 1322
rect 18689 1264 18694 1320
rect 18750 1264 22800 1320
rect 18689 1262 22800 1264
rect 18689 1259 18755 1262
rect 22320 1232 22800 1262
rect 0 914 480 944
rect 3325 914 3391 917
rect 0 912 3391 914
rect 0 856 3330 912
rect 3386 856 3391 912
rect 0 854 3391 856
rect 0 824 480 854
rect 3325 851 3391 854
rect 19374 852 19380 916
rect 19444 914 19450 916
rect 22320 914 22800 944
rect 19444 854 22800 914
rect 19444 852 19450 854
rect 22320 824 22800 854
rect 0 506 480 536
rect 3049 506 3115 509
rect 0 504 3115 506
rect 0 448 3054 504
rect 3110 448 3115 504
rect 0 446 3115 448
rect 0 416 480 446
rect 3049 443 3115 446
rect 17953 506 18019 509
rect 22320 506 22800 536
rect 17953 504 22800 506
rect 17953 448 17958 504
rect 18014 448 22800 504
rect 17953 446 22800 448
rect 17953 443 18019 446
rect 22320 416 22800 446
rect 0 234 480 264
rect 3417 234 3483 237
rect 0 232 3483 234
rect 0 176 3422 232
rect 3478 176 3483 232
rect 0 174 3483 176
rect 0 144 480 174
rect 3417 171 3483 174
rect 18781 234 18847 237
rect 22320 234 22800 264
rect 18781 232 22800 234
rect 18781 176 18786 232
rect 18842 176 22800 232
rect 18781 174 22800 176
rect 18781 171 18847 174
rect 22320 144 22800 174
<< via3 >>
rect 3556 22612 3620 22676
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 11836 19212 11900 19276
rect 12020 19212 12084 19276
rect 4844 19076 4908 19140
rect 9812 19076 9876 19140
rect 17724 19076 17788 19140
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 5396 18940 5460 19004
rect 14044 18940 14108 19004
rect 4844 18532 4908 18596
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 3924 18260 3988 18324
rect 10180 18396 10244 18460
rect 12756 18396 12820 18460
rect 9444 18260 9508 18324
rect 15148 18260 15212 18324
rect 11652 18124 11716 18188
rect 3740 17988 3804 18052
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 18644 17988 18708 18052
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 15332 17640 15396 17644
rect 15332 17584 15346 17640
rect 15346 17584 15396 17640
rect 15332 17580 15396 17584
rect 14412 17444 14476 17508
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 19012 17308 19076 17372
rect 7420 17172 7484 17236
rect 10548 17172 10612 17236
rect 12940 17036 13004 17100
rect 18828 17036 18892 17100
rect 4844 16900 4908 16964
rect 14228 16900 14292 16964
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 9996 16764 10060 16828
rect 17908 16764 17972 16828
rect 10180 16492 10244 16556
rect 17356 16492 17420 16556
rect 19564 16356 19628 16420
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 5212 16220 5276 16284
rect 11836 16220 11900 16284
rect 16436 16084 16500 16148
rect 19380 16008 19444 16012
rect 19380 15952 19394 16008
rect 19394 15952 19444 16008
rect 19380 15948 19444 15952
rect 16252 15872 16316 15876
rect 16252 15816 16266 15872
rect 16266 15816 16316 15872
rect 16252 15812 16316 15816
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 3372 15676 3436 15740
rect 10364 15736 10428 15740
rect 10364 15680 10414 15736
rect 10414 15680 10428 15736
rect 10364 15676 10428 15680
rect 8708 15540 8772 15604
rect 16252 15404 16316 15468
rect 8892 15268 8956 15332
rect 12572 15268 12636 15332
rect 19012 15268 19076 15332
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 10916 15132 10980 15196
rect 13492 15132 13556 15196
rect 19012 14860 19076 14924
rect 18828 14724 18892 14788
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 18828 14588 18892 14652
rect 14044 14452 14108 14516
rect 19932 14452 19996 14516
rect 13676 14316 13740 14380
rect 15884 14316 15948 14380
rect 16620 14316 16684 14380
rect 19380 14180 19444 14244
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 19748 14104 19812 14108
rect 19748 14048 19798 14104
rect 19798 14048 19812 14104
rect 19748 14044 19812 14048
rect 7420 13968 7484 13972
rect 7420 13912 7470 13968
rect 7470 13912 7484 13968
rect 7420 13908 7484 13912
rect 11100 13968 11164 13972
rect 11100 13912 11150 13968
rect 11150 13912 11164 13968
rect 11100 13908 11164 13912
rect 2820 13832 2884 13836
rect 2820 13776 2870 13832
rect 2870 13776 2884 13832
rect 2820 13772 2884 13776
rect 10916 13772 10980 13836
rect 16988 13772 17052 13836
rect 19564 13772 19628 13836
rect 13860 13636 13924 13700
rect 17540 13636 17604 13700
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 8340 13500 8404 13564
rect 15700 13560 15764 13564
rect 15700 13504 15714 13560
rect 15714 13504 15764 13560
rect 15700 13500 15764 13504
rect 16804 13500 16868 13564
rect 19012 13500 19076 13564
rect 6316 13228 6380 13292
rect 8524 13228 8588 13292
rect 8892 13228 8956 13292
rect 16068 13228 16132 13292
rect 10916 13092 10980 13156
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7236 12820 7300 12884
rect 9076 12956 9140 13020
rect 10180 13016 10244 13020
rect 10180 12960 10230 13016
rect 10230 12960 10244 13016
rect 10180 12956 10244 12960
rect 12940 13016 13004 13020
rect 12940 12960 12990 13016
rect 12990 12960 13004 13016
rect 12940 12956 13004 12960
rect 15332 13016 15396 13020
rect 15332 12960 15346 13016
rect 15346 12960 15396 13016
rect 15332 12956 15396 12960
rect 17172 13016 17236 13020
rect 17172 12960 17186 13016
rect 17186 12960 17236 13016
rect 17172 12956 17236 12960
rect 15332 12820 15396 12884
rect 19196 12684 19260 12748
rect 6684 12548 6748 12612
rect 9812 12548 9876 12612
rect 17724 12548 17788 12612
rect 19012 12608 19076 12612
rect 19012 12552 19062 12608
rect 19062 12552 19076 12608
rect 19012 12548 19076 12552
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 6868 12412 6932 12476
rect 6684 12276 6748 12340
rect 8708 12276 8772 12340
rect 7420 12200 7484 12204
rect 7420 12144 7470 12200
rect 7470 12144 7484 12200
rect 7420 12140 7484 12144
rect 8708 12140 8772 12204
rect 9812 12276 9876 12340
rect 10180 12412 10244 12476
rect 11836 12412 11900 12476
rect 16620 12412 16684 12476
rect 19932 12472 19996 12476
rect 19932 12416 19946 12472
rect 19946 12416 19996 12472
rect 19932 12412 19996 12416
rect 13676 12276 13740 12340
rect 16068 12276 16132 12340
rect 9260 12140 9324 12204
rect 18828 12140 18892 12204
rect 19196 12140 19260 12204
rect 3188 12064 3252 12068
rect 3188 12008 3238 12064
rect 3238 12008 3252 12064
rect 3188 12004 3252 12008
rect 7052 12004 7116 12068
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 17356 12004 17420 12068
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 12388 11732 12452 11796
rect 19380 11868 19444 11932
rect 7236 11596 7300 11660
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 9628 11324 9692 11388
rect 12020 11596 12084 11660
rect 13492 11460 13556 11524
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 9996 11384 10060 11388
rect 9996 11328 10010 11384
rect 10010 11328 10060 11384
rect 9996 11324 10060 11328
rect 15700 11324 15764 11388
rect 4844 11052 4908 11116
rect 9444 11052 9508 11116
rect 18828 11188 18892 11252
rect 19012 11188 19076 11252
rect 4844 10916 4908 10980
rect 5396 10916 5460 10980
rect 12756 11052 12820 11116
rect 11652 10916 11716 10980
rect 13676 10916 13740 10980
rect 16804 10976 16868 10980
rect 16804 10920 16818 10976
rect 16818 10920 16868 10976
rect 16804 10916 16868 10920
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 8340 10644 8404 10708
rect 16988 10644 17052 10708
rect 17172 10508 17236 10572
rect 16252 10372 16316 10436
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 15884 10236 15948 10300
rect 20116 10372 20180 10436
rect 12572 10100 12636 10164
rect 12756 10100 12820 10164
rect 19932 10100 19996 10164
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 3556 9556 3620 9620
rect 8708 9964 8772 10028
rect 10364 10024 10428 10028
rect 10364 9968 10378 10024
rect 10378 9968 10428 10024
rect 10364 9964 10428 9968
rect 10732 9828 10796 9892
rect 11652 9888 11716 9892
rect 11652 9832 11702 9888
rect 11702 9832 11716 9888
rect 11652 9828 11716 9832
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 12756 9692 12820 9756
rect 17540 9556 17604 9620
rect 5396 9284 5460 9348
rect 6868 9284 6932 9348
rect 19380 9420 19444 9484
rect 14044 9284 14108 9348
rect 17540 9344 17604 9348
rect 17540 9288 17590 9344
rect 17590 9288 17604 9344
rect 17540 9284 17604 9288
rect 17724 9284 17788 9348
rect 18828 9284 18892 9348
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 3188 9148 3252 9212
rect 14412 9148 14476 9212
rect 15516 9148 15580 9212
rect 6684 9012 6748 9076
rect 9076 9012 9140 9076
rect 6868 8740 6932 8804
rect 7236 8740 7300 8804
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 13308 8876 13372 8940
rect 16620 9012 16684 9076
rect 19196 9012 19260 9076
rect 15516 8876 15580 8940
rect 12204 8740 12268 8804
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 10548 8604 10612 8668
rect 10916 8604 10980 8668
rect 13492 8604 13556 8668
rect 14044 8604 14108 8668
rect 11836 8468 11900 8532
rect 18828 8604 18892 8668
rect 11100 8332 11164 8396
rect 13124 8332 13188 8396
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 7604 8060 7668 8124
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 9076 7924 9140 7988
rect 9996 8060 10060 8124
rect 10548 8120 10612 8124
rect 10548 8064 10562 8120
rect 10562 8064 10612 8120
rect 10548 8060 10612 8064
rect 15332 8060 15396 8124
rect 10732 7788 10796 7852
rect 10916 7652 10980 7716
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18828 8196 18892 8260
rect 19380 8120 19444 8124
rect 19380 8064 19394 8120
rect 19394 8064 19444 8120
rect 19380 8060 19444 8064
rect 20116 7924 20180 7988
rect 17172 7652 17236 7716
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 13676 7516 13740 7580
rect 15332 7516 15396 7580
rect 19012 7516 19076 7580
rect 4844 7380 4908 7444
rect 15148 7244 15212 7308
rect 19932 7516 19996 7580
rect 8340 7108 8404 7172
rect 12388 7108 12452 7172
rect 12940 7108 13004 7172
rect 13308 7108 13372 7172
rect 13860 7108 13924 7172
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 3740 6972 3804 7036
rect 6316 6972 6380 7036
rect 8340 6972 8404 7036
rect 19380 7108 19444 7172
rect 19012 6972 19076 7036
rect 18828 6836 18892 6900
rect 19748 6836 19812 6900
rect 11652 6564 11716 6628
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 2820 6428 2884 6492
rect 8340 6428 8404 6492
rect 9444 6428 9508 6492
rect 9812 6488 9876 6492
rect 9812 6432 9862 6488
rect 9862 6432 9876 6488
rect 9812 6428 9876 6432
rect 12388 6428 12452 6492
rect 12756 6488 12820 6492
rect 12756 6432 12806 6488
rect 12806 6432 12820 6488
rect 12756 6428 12820 6432
rect 13124 6428 13188 6492
rect 13676 6428 13740 6492
rect 17172 6428 17236 6492
rect 3372 6292 3436 6356
rect 16436 6292 16500 6356
rect 19012 6292 19076 6356
rect 19012 6216 19076 6220
rect 19012 6160 19026 6216
rect 19026 6160 19076 6216
rect 7052 6080 7116 6084
rect 7052 6024 7102 6080
rect 7102 6024 7116 6080
rect 7052 6020 7116 6024
rect 19012 6156 19076 6160
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 7052 5884 7116 5948
rect 17724 5884 17788 5948
rect 8892 5808 8956 5812
rect 8892 5752 8942 5808
rect 8942 5752 8956 5808
rect 5212 5612 5276 5676
rect 7604 5612 7668 5676
rect 8892 5748 8956 5752
rect 9444 5808 9508 5812
rect 9444 5752 9458 5808
rect 9458 5752 9508 5808
rect 9444 5748 9508 5752
rect 10548 5748 10612 5812
rect 11652 5536 11716 5540
rect 11652 5480 11702 5536
rect 11702 5480 11716 5536
rect 11652 5476 11716 5480
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 19748 5340 19812 5404
rect 4844 5068 4908 5132
rect 14228 5204 14292 5268
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 9444 4856 9508 4860
rect 9444 4800 9494 4856
rect 9494 4800 9508 4856
rect 9444 4796 9508 4800
rect 9260 4524 9324 4588
rect 12940 4388 13004 4452
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 6868 4252 6932 4316
rect 8892 4252 8956 4316
rect 12756 4252 12820 4316
rect 3188 4176 3252 4180
rect 3188 4120 3202 4176
rect 3202 4120 3252 4176
rect 3188 4116 3252 4120
rect 5396 4116 5460 4180
rect 5212 3980 5276 4044
rect 7420 3980 7484 4044
rect 12572 3980 12636 4044
rect 18644 3980 18708 4044
rect 9076 3844 9140 3908
rect 14044 3844 14108 3908
rect 16620 3844 16684 3908
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 3188 3708 3252 3772
rect 3924 3708 3988 3772
rect 9076 3436 9140 3500
rect 9628 3300 9692 3364
rect 17172 3300 17236 3364
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7604 3164 7668 3228
rect 8708 3164 8772 3228
rect 17540 3164 17604 3228
rect 19012 3164 19076 3228
rect 7236 2892 7300 2956
rect 11652 2892 11716 2956
rect 12388 2756 12452 2820
rect 19196 2816 19260 2820
rect 19196 2760 19210 2816
rect 19210 2760 19260 2816
rect 19196 2756 19260 2760
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 8340 2620 8404 2684
rect 17908 2620 17972 2684
rect 8708 2484 8772 2548
rect 18828 2544 18892 2548
rect 18828 2488 18842 2544
rect 18842 2488 18892 2544
rect 18828 2484 18892 2488
rect 9444 2348 9508 2412
rect 19564 2348 19628 2412
rect 6684 2212 6748 2276
rect 19748 2212 19812 2276
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
rect 7052 2076 7116 2140
rect 19380 852 19444 916
<< metal4 >>
rect 3555 22676 3621 22677
rect 3555 22612 3556 22676
rect 3620 22612 3621 22676
rect 3555 22611 3621 22612
rect 3371 15740 3437 15741
rect 3371 15676 3372 15740
rect 3436 15676 3437 15740
rect 3371 15675 3437 15676
rect 2819 13836 2885 13837
rect 2819 13772 2820 13836
rect 2884 13772 2885 13836
rect 2819 13771 2885 13772
rect 2822 6493 2882 13771
rect 3187 12068 3253 12069
rect 3187 12004 3188 12068
rect 3252 12004 3253 12068
rect 3187 12003 3253 12004
rect 3190 9213 3250 12003
rect 3187 9212 3253 9213
rect 3187 9148 3188 9212
rect 3252 9148 3253 9212
rect 3187 9147 3253 9148
rect 2819 6492 2885 6493
rect 2819 6428 2820 6492
rect 2884 6428 2885 6492
rect 2819 6427 2885 6428
rect 3374 6357 3434 15675
rect 3558 9621 3618 22611
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 4843 19140 4909 19141
rect 4843 19076 4844 19140
rect 4908 19076 4909 19140
rect 4843 19075 4909 19076
rect 4846 18597 4906 19075
rect 7808 19072 8128 20096
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 9811 19140 9877 19141
rect 9811 19076 9812 19140
rect 9876 19076 9877 19140
rect 9811 19075 9877 19076
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 5395 19004 5461 19005
rect 5395 18940 5396 19004
rect 5460 18940 5461 19004
rect 5395 18939 5461 18940
rect 4843 18596 4909 18597
rect 4843 18532 4844 18596
rect 4908 18532 4909 18596
rect 4843 18531 4909 18532
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 3923 18324 3989 18325
rect 3923 18260 3924 18324
rect 3988 18260 3989 18324
rect 3923 18259 3989 18260
rect 3739 18052 3805 18053
rect 3739 17988 3740 18052
rect 3804 17988 3805 18052
rect 3739 17987 3805 17988
rect 3555 9620 3621 9621
rect 3555 9556 3556 9620
rect 3620 9556 3621 9620
rect 3555 9555 3621 9556
rect 3742 7037 3802 17987
rect 3739 7036 3805 7037
rect 3739 6972 3740 7036
rect 3804 6972 3805 7036
rect 3739 6971 3805 6972
rect 3371 6356 3437 6357
rect 3371 6292 3372 6356
rect 3436 6292 3437 6356
rect 3371 6291 3437 6292
rect 3187 4180 3253 4181
rect 3187 4116 3188 4180
rect 3252 4116 3253 4180
rect 3187 4115 3253 4116
rect 3190 3773 3250 4115
rect 3926 3773 3986 18259
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4843 16964 4909 16965
rect 4843 16900 4844 16964
rect 4908 16900 4909 16964
rect 4843 16899 4909 16900
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4846 11117 4906 16899
rect 5211 16284 5277 16285
rect 5211 16220 5212 16284
rect 5276 16220 5277 16284
rect 5211 16219 5277 16220
rect 4843 11116 4909 11117
rect 4843 11052 4844 11116
rect 4908 11052 4909 11116
rect 4843 11051 4909 11052
rect 4843 10980 4909 10981
rect 4843 10916 4844 10980
rect 4908 10916 4909 10980
rect 4843 10915 4909 10916
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4846 7445 4906 10915
rect 4843 7444 4909 7445
rect 4843 7380 4844 7444
rect 4908 7380 4909 7444
rect 4843 7379 4909 7380
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4846 5133 4906 7379
rect 5214 5677 5274 16219
rect 5398 10981 5458 18939
rect 7808 17984 8128 19008
rect 9443 18324 9509 18325
rect 9443 18260 9444 18324
rect 9508 18260 9509 18324
rect 9443 18259 9509 18260
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7419 17236 7485 17237
rect 7419 17172 7420 17236
rect 7484 17172 7485 17236
rect 7419 17171 7485 17172
rect 7422 13973 7482 17171
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 8707 15604 8773 15605
rect 8707 15540 8708 15604
rect 8772 15540 8773 15604
rect 8707 15539 8773 15540
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7419 13972 7485 13973
rect 7419 13908 7420 13972
rect 7484 13908 7485 13972
rect 7419 13907 7485 13908
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 6315 13292 6381 13293
rect 6315 13228 6316 13292
rect 6380 13228 6381 13292
rect 6315 13227 6381 13228
rect 5395 10980 5461 10981
rect 5395 10916 5396 10980
rect 5460 10916 5461 10980
rect 5395 10915 5461 10916
rect 5395 9348 5461 9349
rect 5395 9284 5396 9348
rect 5460 9284 5461 9348
rect 5395 9283 5461 9284
rect 5211 5676 5277 5677
rect 5211 5612 5212 5676
rect 5276 5612 5277 5676
rect 5211 5611 5277 5612
rect 4843 5132 4909 5133
rect 4843 5068 4844 5132
rect 4908 5068 4909 5132
rect 4843 5067 4909 5068
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 3187 3772 3253 3773
rect 3187 3708 3188 3772
rect 3252 3708 3253 3772
rect 3187 3707 3253 3708
rect 3923 3772 3989 3773
rect 3923 3708 3924 3772
rect 3988 3708 3989 3772
rect 3923 3707 3989 3708
rect 4376 3296 4696 4320
rect 5214 4045 5274 5611
rect 5398 4181 5458 9283
rect 6318 7037 6378 13227
rect 7235 12884 7301 12885
rect 7235 12820 7236 12884
rect 7300 12820 7301 12884
rect 7235 12819 7301 12820
rect 6683 12612 6749 12613
rect 6683 12548 6684 12612
rect 6748 12548 6749 12612
rect 6683 12547 6749 12548
rect 6686 12341 6746 12547
rect 6867 12476 6933 12477
rect 6867 12412 6868 12476
rect 6932 12412 6933 12476
rect 6867 12411 6933 12412
rect 6683 12340 6749 12341
rect 6683 12276 6684 12340
rect 6748 12276 6749 12340
rect 6683 12275 6749 12276
rect 6870 9349 6930 12411
rect 7051 12068 7117 12069
rect 7051 12004 7052 12068
rect 7116 12004 7117 12068
rect 7051 12003 7117 12004
rect 6867 9348 6933 9349
rect 6867 9284 6868 9348
rect 6932 9284 6933 9348
rect 6867 9283 6933 9284
rect 6683 9076 6749 9077
rect 6683 9012 6684 9076
rect 6748 9012 6749 9076
rect 6683 9011 6749 9012
rect 6315 7036 6381 7037
rect 6315 6972 6316 7036
rect 6380 6972 6381 7036
rect 6315 6971 6381 6972
rect 5395 4180 5461 4181
rect 5395 4116 5396 4180
rect 5460 4116 5461 4180
rect 5395 4115 5461 4116
rect 5211 4044 5277 4045
rect 5211 3980 5212 4044
rect 5276 3980 5277 4044
rect 5211 3979 5277 3980
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 6686 2277 6746 9011
rect 6867 8804 6933 8805
rect 6867 8740 6868 8804
rect 6932 8740 6933 8804
rect 6867 8739 6933 8740
rect 6870 4317 6930 8739
rect 7054 6085 7114 12003
rect 7238 11661 7298 12819
rect 7808 12544 8128 13568
rect 8339 13564 8405 13565
rect 8339 13500 8340 13564
rect 8404 13500 8405 13564
rect 8339 13499 8405 13500
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7419 12204 7485 12205
rect 7419 12140 7420 12204
rect 7484 12140 7485 12204
rect 7419 12139 7485 12140
rect 7235 11660 7301 11661
rect 7235 11596 7236 11660
rect 7300 11596 7301 11660
rect 7235 11595 7301 11596
rect 7235 8804 7301 8805
rect 7235 8740 7236 8804
rect 7300 8740 7301 8804
rect 7235 8739 7301 8740
rect 7051 6084 7117 6085
rect 7051 6020 7052 6084
rect 7116 6020 7117 6084
rect 7051 6019 7117 6020
rect 7051 5948 7117 5949
rect 7051 5884 7052 5948
rect 7116 5884 7117 5948
rect 7051 5883 7117 5884
rect 6867 4316 6933 4317
rect 6867 4252 6868 4316
rect 6932 4252 6933 4316
rect 6867 4251 6933 4252
rect 6683 2276 6749 2277
rect 6683 2212 6684 2276
rect 6748 2212 6749 2276
rect 6683 2211 6749 2212
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7054 2141 7114 5883
rect 7238 2957 7298 8739
rect 7422 4045 7482 12139
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 8342 10709 8402 13499
rect 8523 13292 8589 13293
rect 8523 13228 8524 13292
rect 8588 13228 8589 13292
rect 8523 13227 8589 13228
rect 8339 10708 8405 10709
rect 8339 10644 8340 10708
rect 8404 10644 8405 10708
rect 8339 10643 8405 10644
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 8526 9890 8586 13227
rect 8710 12341 8770 15539
rect 8891 15332 8957 15333
rect 8891 15268 8892 15332
rect 8956 15268 8957 15332
rect 8891 15267 8957 15268
rect 8894 13293 8954 15267
rect 8891 13292 8957 13293
rect 8891 13228 8892 13292
rect 8956 13228 8957 13292
rect 8891 13227 8957 13228
rect 8707 12340 8773 12341
rect 8707 12276 8708 12340
rect 8772 12276 8773 12340
rect 8707 12275 8773 12276
rect 8707 12204 8773 12205
rect 8707 12140 8708 12204
rect 8772 12140 8773 12204
rect 8707 12139 8773 12140
rect 8710 10029 8770 12139
rect 8707 10028 8773 10029
rect 8707 9964 8708 10028
rect 8772 9964 8773 10028
rect 8707 9963 8773 9964
rect 8526 9830 8770 9890
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7603 8124 7669 8125
rect 7603 8060 7604 8124
rect 7668 8060 7669 8124
rect 7603 8059 7669 8060
rect 7606 5677 7666 8059
rect 7808 7104 8128 8128
rect 8339 7172 8405 7173
rect 8339 7170 8340 7172
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 8204 7110 8340 7170
rect 8204 6218 8264 7110
rect 8339 7108 8340 7110
rect 8404 7108 8405 7172
rect 8339 7107 8405 7108
rect 8339 7036 8405 7037
rect 8339 6972 8340 7036
rect 8404 6972 8405 7036
rect 8339 6971 8405 6972
rect 8342 6493 8402 6971
rect 8339 6492 8405 6493
rect 8339 6428 8340 6492
rect 8404 6428 8405 6492
rect 8339 6427 8405 6428
rect 8204 6158 8402 6218
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7603 5676 7669 5677
rect 7603 5612 7604 5676
rect 7668 5612 7669 5676
rect 7603 5611 7669 5612
rect 7419 4044 7485 4045
rect 7419 3980 7420 4044
rect 7484 3980 7485 4044
rect 7419 3979 7485 3980
rect 7606 3229 7666 5611
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7603 3228 7669 3229
rect 7603 3164 7604 3228
rect 7668 3164 7669 3228
rect 7603 3163 7669 3164
rect 7235 2956 7301 2957
rect 7235 2892 7236 2956
rect 7300 2892 7301 2956
rect 7235 2891 7301 2892
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7051 2140 7117 2141
rect 7051 2076 7052 2140
rect 7116 2076 7117 2140
rect 7808 2128 8128 2688
rect 8342 2685 8402 6158
rect 8710 3229 8770 9830
rect 8894 5813 8954 13227
rect 9075 13020 9141 13021
rect 9075 12956 9076 13020
rect 9140 12956 9141 13020
rect 9075 12955 9141 12956
rect 9078 9077 9138 12955
rect 9259 12204 9325 12205
rect 9259 12140 9260 12204
rect 9324 12140 9325 12204
rect 9259 12139 9325 12140
rect 9075 9076 9141 9077
rect 9075 9012 9076 9076
rect 9140 9012 9141 9076
rect 9075 9011 9141 9012
rect 9075 7988 9141 7989
rect 9075 7924 9076 7988
rect 9140 7924 9141 7988
rect 9075 7923 9141 7924
rect 8891 5812 8957 5813
rect 8891 5748 8892 5812
rect 8956 5748 8957 5812
rect 8891 5747 8957 5748
rect 8891 4316 8957 4317
rect 8891 4252 8892 4316
rect 8956 4252 8957 4316
rect 8891 4251 8957 4252
rect 8894 3498 8954 4251
rect 9078 3909 9138 7923
rect 9262 4589 9322 12139
rect 9446 11117 9506 18259
rect 9814 12613 9874 19075
rect 11240 18528 11560 19552
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 11835 19276 11901 19277
rect 11835 19212 11836 19276
rect 11900 19212 11901 19276
rect 11835 19211 11901 19212
rect 12019 19276 12085 19277
rect 12019 19212 12020 19276
rect 12084 19212 12085 19276
rect 12019 19211 12085 19212
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 10179 18460 10245 18461
rect 10179 18396 10180 18460
rect 10244 18396 10245 18460
rect 10179 18395 10245 18396
rect 9995 16828 10061 16829
rect 9995 16764 9996 16828
rect 10060 16764 10061 16828
rect 9995 16763 10061 16764
rect 9811 12612 9877 12613
rect 9811 12548 9812 12612
rect 9876 12548 9877 12612
rect 9811 12547 9877 12548
rect 9811 12340 9877 12341
rect 9811 12276 9812 12340
rect 9876 12276 9877 12340
rect 9811 12275 9877 12276
rect 9627 11388 9693 11389
rect 9627 11324 9628 11388
rect 9692 11324 9693 11388
rect 9627 11323 9693 11324
rect 9443 11116 9509 11117
rect 9443 11052 9444 11116
rect 9508 11052 9509 11116
rect 9443 11051 9509 11052
rect 9443 6492 9509 6493
rect 9443 6428 9444 6492
rect 9508 6428 9509 6492
rect 9443 6427 9509 6428
rect 9446 5813 9506 6427
rect 9443 5812 9509 5813
rect 9443 5748 9444 5812
rect 9508 5748 9509 5812
rect 9443 5747 9509 5748
rect 9443 4860 9509 4861
rect 9443 4796 9444 4860
rect 9508 4796 9509 4860
rect 9443 4795 9509 4796
rect 9259 4588 9325 4589
rect 9259 4524 9260 4588
rect 9324 4524 9325 4588
rect 9259 4523 9325 4524
rect 9075 3908 9141 3909
rect 9075 3844 9076 3908
rect 9140 3844 9141 3908
rect 9075 3843 9141 3844
rect 9075 3500 9141 3501
rect 9075 3498 9076 3500
rect 8894 3438 9076 3498
rect 9075 3436 9076 3438
rect 9140 3436 9141 3500
rect 9075 3435 9141 3436
rect 8707 3228 8773 3229
rect 8707 3164 8708 3228
rect 8772 3164 8773 3228
rect 8707 3163 8773 3164
rect 8339 2684 8405 2685
rect 8339 2620 8340 2684
rect 8404 2620 8405 2684
rect 8339 2619 8405 2620
rect 8710 2549 8770 3163
rect 8707 2548 8773 2549
rect 8707 2484 8708 2548
rect 8772 2484 8773 2548
rect 8707 2483 8773 2484
rect 9446 2413 9506 4795
rect 9630 3365 9690 11323
rect 9814 6493 9874 12275
rect 9998 11389 10058 16763
rect 10182 16557 10242 18395
rect 11240 17440 11560 18464
rect 11651 18188 11717 18189
rect 11651 18124 11652 18188
rect 11716 18124 11717 18188
rect 11651 18123 11717 18124
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 10547 17236 10613 17237
rect 10547 17172 10548 17236
rect 10612 17172 10613 17236
rect 10547 17171 10613 17172
rect 10179 16556 10245 16557
rect 10179 16492 10180 16556
rect 10244 16492 10245 16556
rect 10179 16491 10245 16492
rect 10182 13021 10242 16491
rect 10363 15740 10429 15741
rect 10363 15676 10364 15740
rect 10428 15676 10429 15740
rect 10363 15675 10429 15676
rect 10179 13020 10245 13021
rect 10179 12956 10180 13020
rect 10244 12956 10245 13020
rect 10179 12955 10245 12956
rect 10179 12476 10245 12477
rect 10179 12412 10180 12476
rect 10244 12412 10245 12476
rect 10179 12411 10245 12412
rect 9995 11388 10061 11389
rect 9995 11324 9996 11388
rect 10060 11324 10061 11388
rect 9995 11323 10061 11324
rect 10182 8530 10242 12411
rect 10366 10029 10426 15675
rect 10363 10028 10429 10029
rect 10363 9964 10364 10028
rect 10428 9964 10429 10028
rect 10363 9963 10429 9964
rect 10550 8669 10610 17171
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 10915 15196 10981 15197
rect 10915 15132 10916 15196
rect 10980 15132 10981 15196
rect 10915 15131 10981 15132
rect 10918 13837 10978 15131
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11099 13972 11165 13973
rect 11099 13908 11100 13972
rect 11164 13908 11165 13972
rect 11099 13907 11165 13908
rect 10915 13836 10981 13837
rect 10915 13772 10916 13836
rect 10980 13772 10981 13836
rect 10915 13771 10981 13772
rect 10918 13157 10978 13771
rect 10915 13156 10981 13157
rect 10915 13092 10916 13156
rect 10980 13092 10981 13156
rect 10915 13091 10981 13092
rect 10731 9892 10797 9893
rect 10731 9828 10732 9892
rect 10796 9828 10797 9892
rect 10731 9827 10797 9828
rect 10547 8668 10613 8669
rect 10547 8604 10548 8668
rect 10612 8604 10613 8668
rect 10547 8603 10613 8604
rect 9998 8470 10242 8530
rect 9998 8125 10058 8470
rect 9995 8124 10061 8125
rect 9995 8060 9996 8124
rect 10060 8060 10061 8124
rect 9995 8059 10061 8060
rect 10547 8124 10613 8125
rect 10547 8060 10548 8124
rect 10612 8060 10613 8124
rect 10547 8059 10613 8060
rect 9811 6492 9877 6493
rect 9811 6428 9812 6492
rect 9876 6428 9877 6492
rect 9811 6427 9877 6428
rect 10550 5813 10610 8059
rect 10734 7853 10794 9827
rect 10915 8668 10981 8669
rect 10915 8604 10916 8668
rect 10980 8604 10981 8668
rect 10915 8603 10981 8604
rect 10731 7852 10797 7853
rect 10731 7788 10732 7852
rect 10796 7788 10797 7852
rect 10731 7787 10797 7788
rect 10918 7717 10978 8603
rect 11102 8397 11162 13907
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11654 10981 11714 18123
rect 11838 16285 11898 19211
rect 11835 16284 11901 16285
rect 11835 16220 11836 16284
rect 11900 16220 11901 16284
rect 11835 16219 11901 16220
rect 11838 12477 11898 16219
rect 11835 12476 11901 12477
rect 11835 12412 11836 12476
rect 11900 12412 11901 12476
rect 11835 12411 11901 12412
rect 12022 11661 12082 19211
rect 14672 19072 14992 20096
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 17723 19140 17789 19141
rect 17723 19076 17724 19140
rect 17788 19076 17789 19140
rect 17723 19075 17789 19076
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14043 19004 14109 19005
rect 14043 18940 14044 19004
rect 14108 18940 14109 19004
rect 14043 18939 14109 18940
rect 12755 18460 12821 18461
rect 12755 18396 12756 18460
rect 12820 18396 12821 18460
rect 12755 18395 12821 18396
rect 12571 15332 12637 15333
rect 12571 15268 12572 15332
rect 12636 15268 12637 15332
rect 12571 15267 12637 15268
rect 12387 11796 12453 11797
rect 12387 11732 12388 11796
rect 12452 11732 12453 11796
rect 12387 11731 12453 11732
rect 12019 11660 12085 11661
rect 12019 11596 12020 11660
rect 12084 11596 12085 11660
rect 12019 11595 12085 11596
rect 11651 10980 11717 10981
rect 11651 10916 11652 10980
rect 11716 10916 11717 10980
rect 11651 10915 11717 10916
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11651 9892 11717 9893
rect 11651 9828 11652 9892
rect 11716 9828 11717 9892
rect 11651 9827 11717 9828
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11099 8396 11165 8397
rect 11099 8332 11100 8396
rect 11164 8332 11165 8396
rect 11099 8331 11165 8332
rect 10915 7716 10981 7717
rect 10915 7652 10916 7716
rect 10980 7652 10981 7716
rect 10915 7651 10981 7652
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11654 6629 11714 9827
rect 12203 8804 12269 8805
rect 12203 8740 12204 8804
rect 12268 8740 12269 8804
rect 12203 8739 12269 8740
rect 11835 8532 11901 8533
rect 11835 8468 11836 8532
rect 11900 8530 11901 8532
rect 12206 8530 12266 8739
rect 11900 8470 12266 8530
rect 11900 8468 11901 8470
rect 11835 8467 11901 8468
rect 12390 7173 12450 11731
rect 12574 10165 12634 15267
rect 12758 11117 12818 18395
rect 12939 17100 13005 17101
rect 12939 17036 12940 17100
rect 13004 17036 13005 17100
rect 12939 17035 13005 17036
rect 12942 16282 13002 17035
rect 12942 16222 13186 16282
rect 12939 13020 13005 13021
rect 12939 12956 12940 13020
rect 13004 12956 13005 13020
rect 12939 12955 13005 12956
rect 12755 11116 12821 11117
rect 12755 11052 12756 11116
rect 12820 11052 12821 11116
rect 12755 11051 12821 11052
rect 12571 10164 12637 10165
rect 12571 10100 12572 10164
rect 12636 10100 12637 10164
rect 12571 10099 12637 10100
rect 12755 10164 12821 10165
rect 12755 10100 12756 10164
rect 12820 10100 12821 10164
rect 12755 10099 12821 10100
rect 12758 9757 12818 10099
rect 12755 9756 12821 9757
rect 12755 9692 12756 9756
rect 12820 9692 12821 9756
rect 12755 9691 12821 9692
rect 12942 9618 13002 12955
rect 12574 9558 13002 9618
rect 12387 7172 12453 7173
rect 12387 7108 12388 7172
rect 12452 7108 12453 7172
rect 12387 7107 12453 7108
rect 11651 6628 11717 6629
rect 11651 6564 11652 6628
rect 11716 6564 11717 6628
rect 11651 6563 11717 6564
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 10547 5812 10613 5813
rect 10547 5748 10548 5812
rect 10612 5748 10613 5812
rect 10547 5747 10613 5748
rect 11240 5472 11560 6496
rect 12387 6492 12453 6493
rect 12387 6428 12388 6492
rect 12452 6428 12453 6492
rect 12387 6427 12453 6428
rect 11651 5540 11717 5541
rect 11651 5476 11652 5540
rect 11716 5476 11717 5540
rect 11651 5475 11717 5476
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 9627 3364 9693 3365
rect 9627 3300 9628 3364
rect 9692 3300 9693 3364
rect 9627 3299 9693 3300
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 9443 2412 9509 2413
rect 9443 2348 9444 2412
rect 9508 2348 9509 2412
rect 9443 2347 9509 2348
rect 11240 2208 11560 3232
rect 11654 2957 11714 5475
rect 11651 2956 11717 2957
rect 11651 2892 11652 2956
rect 11716 2892 11717 2956
rect 11651 2891 11717 2892
rect 12390 2821 12450 6427
rect 12574 4045 12634 9558
rect 13126 8397 13186 16222
rect 13491 15196 13557 15197
rect 13491 15132 13492 15196
rect 13556 15132 13557 15196
rect 13491 15131 13557 15132
rect 13494 11525 13554 15131
rect 14046 14517 14106 18939
rect 14672 17984 14992 19008
rect 15147 18324 15213 18325
rect 15147 18260 15148 18324
rect 15212 18260 15213 18324
rect 15147 18259 15213 18260
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14411 17508 14477 17509
rect 14411 17444 14412 17508
rect 14476 17444 14477 17508
rect 14411 17443 14477 17444
rect 14227 16964 14293 16965
rect 14227 16900 14228 16964
rect 14292 16900 14293 16964
rect 14227 16899 14293 16900
rect 14043 14516 14109 14517
rect 14043 14452 14044 14516
rect 14108 14452 14109 14516
rect 14043 14451 14109 14452
rect 13675 14380 13741 14381
rect 13675 14316 13676 14380
rect 13740 14316 13741 14380
rect 13675 14315 13741 14316
rect 13678 12341 13738 14315
rect 13859 13700 13925 13701
rect 13859 13636 13860 13700
rect 13924 13636 13925 13700
rect 13859 13635 13925 13636
rect 13675 12340 13741 12341
rect 13675 12276 13676 12340
rect 13740 12276 13741 12340
rect 13675 12275 13741 12276
rect 13491 11524 13557 11525
rect 13491 11460 13492 11524
rect 13556 11460 13557 11524
rect 13491 11459 13557 11460
rect 13307 8940 13373 8941
rect 13307 8876 13308 8940
rect 13372 8876 13373 8940
rect 13307 8875 13373 8876
rect 13123 8396 13189 8397
rect 13123 8332 13124 8396
rect 13188 8332 13189 8396
rect 13123 8331 13189 8332
rect 12939 7172 13005 7173
rect 12939 7108 12940 7172
rect 13004 7108 13005 7172
rect 12939 7107 13005 7108
rect 12755 6492 12821 6493
rect 12755 6428 12756 6492
rect 12820 6428 12821 6492
rect 12755 6427 12821 6428
rect 12758 4317 12818 6427
rect 12942 4453 13002 7107
rect 13126 6493 13186 8331
rect 13310 7173 13370 8875
rect 13494 8669 13554 11459
rect 13675 10980 13741 10981
rect 13675 10916 13676 10980
rect 13740 10916 13741 10980
rect 13675 10915 13741 10916
rect 13491 8668 13557 8669
rect 13491 8604 13492 8668
rect 13556 8604 13557 8668
rect 13491 8603 13557 8604
rect 13678 7581 13738 10915
rect 13675 7580 13741 7581
rect 13675 7516 13676 7580
rect 13740 7516 13741 7580
rect 13675 7515 13741 7516
rect 13862 7173 13922 13635
rect 14043 9348 14109 9349
rect 14043 9284 14044 9348
rect 14108 9284 14109 9348
rect 14043 9283 14109 9284
rect 14046 8669 14106 9283
rect 14043 8668 14109 8669
rect 14043 8604 14044 8668
rect 14108 8604 14109 8668
rect 14043 8603 14109 8604
rect 13307 7172 13373 7173
rect 13307 7108 13308 7172
rect 13372 7108 13373 7172
rect 13307 7107 13373 7108
rect 13859 7172 13925 7173
rect 13859 7108 13860 7172
rect 13924 7108 13925 7172
rect 13859 7107 13925 7108
rect 13123 6492 13189 6493
rect 13123 6428 13124 6492
rect 13188 6428 13189 6492
rect 13123 6427 13189 6428
rect 13675 6492 13741 6493
rect 13675 6428 13676 6492
rect 13740 6428 13741 6492
rect 13675 6427 13741 6428
rect 13678 5538 13738 6427
rect 13678 5478 14106 5538
rect 12939 4452 13005 4453
rect 12939 4388 12940 4452
rect 13004 4388 13005 4452
rect 12939 4387 13005 4388
rect 12755 4316 12821 4317
rect 12755 4252 12756 4316
rect 12820 4252 12821 4316
rect 12755 4251 12821 4252
rect 12571 4044 12637 4045
rect 12571 3980 12572 4044
rect 12636 3980 12637 4044
rect 12571 3979 12637 3980
rect 14046 3909 14106 5478
rect 14230 5269 14290 16899
rect 14414 9213 14474 17443
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14411 9212 14477 9213
rect 14411 9148 14412 9212
rect 14476 9148 14477 9212
rect 14411 9147 14477 9148
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 15150 7309 15210 18259
rect 15331 17644 15397 17645
rect 15331 17580 15332 17644
rect 15396 17580 15397 17644
rect 15331 17579 15397 17580
rect 15334 13021 15394 17579
rect 17355 16556 17421 16557
rect 17355 16492 17356 16556
rect 17420 16492 17421 16556
rect 17355 16491 17421 16492
rect 16435 16148 16501 16149
rect 16435 16084 16436 16148
rect 16500 16084 16501 16148
rect 16435 16083 16501 16084
rect 16251 15876 16317 15877
rect 16251 15812 16252 15876
rect 16316 15812 16317 15876
rect 16251 15811 16317 15812
rect 16254 15469 16314 15811
rect 16251 15468 16317 15469
rect 16251 15404 16252 15468
rect 16316 15404 16317 15468
rect 16251 15403 16317 15404
rect 15883 14380 15949 14381
rect 15883 14316 15884 14380
rect 15948 14316 15949 14380
rect 15883 14315 15949 14316
rect 15699 13564 15765 13565
rect 15699 13500 15700 13564
rect 15764 13500 15765 13564
rect 15699 13499 15765 13500
rect 15331 13020 15397 13021
rect 15331 12956 15332 13020
rect 15396 12956 15397 13020
rect 15331 12955 15397 12956
rect 15331 12884 15397 12885
rect 15331 12820 15332 12884
rect 15396 12820 15397 12884
rect 15331 12819 15397 12820
rect 15334 8125 15394 12819
rect 15702 11389 15762 13499
rect 15699 11388 15765 11389
rect 15699 11324 15700 11388
rect 15764 11324 15765 11388
rect 15699 11323 15765 11324
rect 15886 10301 15946 14315
rect 16067 13292 16133 13293
rect 16067 13228 16068 13292
rect 16132 13228 16133 13292
rect 16067 13227 16133 13228
rect 16070 12341 16130 13227
rect 16067 12340 16133 12341
rect 16067 12276 16068 12340
rect 16132 12276 16133 12340
rect 16067 12275 16133 12276
rect 16254 10437 16314 15403
rect 16251 10436 16317 10437
rect 16251 10372 16252 10436
rect 16316 10372 16317 10436
rect 16251 10371 16317 10372
rect 15883 10300 15949 10301
rect 15883 10236 15884 10300
rect 15948 10236 15949 10300
rect 15883 10235 15949 10236
rect 15515 9212 15581 9213
rect 15515 9148 15516 9212
rect 15580 9148 15581 9212
rect 15515 9147 15581 9148
rect 15518 8941 15578 9147
rect 15515 8940 15581 8941
rect 15515 8876 15516 8940
rect 15580 8876 15581 8940
rect 15515 8875 15581 8876
rect 15331 8124 15397 8125
rect 15331 8060 15332 8124
rect 15396 8060 15397 8124
rect 15331 8059 15397 8060
rect 15334 7581 15394 8059
rect 15331 7580 15397 7581
rect 15331 7516 15332 7580
rect 15396 7516 15397 7580
rect 15331 7515 15397 7516
rect 15147 7308 15213 7309
rect 15147 7244 15148 7308
rect 15212 7244 15213 7308
rect 15147 7243 15213 7244
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 16438 6357 16498 16083
rect 16619 14380 16685 14381
rect 16619 14316 16620 14380
rect 16684 14316 16685 14380
rect 16619 14315 16685 14316
rect 16622 12477 16682 14315
rect 16987 13836 17053 13837
rect 16987 13772 16988 13836
rect 17052 13772 17053 13836
rect 16987 13771 17053 13772
rect 16803 13564 16869 13565
rect 16803 13500 16804 13564
rect 16868 13500 16869 13564
rect 16803 13499 16869 13500
rect 16619 12476 16685 12477
rect 16619 12412 16620 12476
rect 16684 12412 16685 12476
rect 16619 12411 16685 12412
rect 16806 10981 16866 13499
rect 16803 10980 16869 10981
rect 16803 10916 16804 10980
rect 16868 10916 16869 10980
rect 16803 10915 16869 10916
rect 16990 10709 17050 13771
rect 17171 13020 17237 13021
rect 17171 12956 17172 13020
rect 17236 12956 17237 13020
rect 17171 12955 17237 12956
rect 16987 10708 17053 10709
rect 16987 10644 16988 10708
rect 17052 10644 17053 10708
rect 16987 10643 17053 10644
rect 17174 10573 17234 12955
rect 17358 12069 17418 16491
rect 17539 13700 17605 13701
rect 17539 13636 17540 13700
rect 17604 13636 17605 13700
rect 17539 13635 17605 13636
rect 17355 12068 17421 12069
rect 17355 12004 17356 12068
rect 17420 12004 17421 12068
rect 17355 12003 17421 12004
rect 17171 10572 17237 10573
rect 17171 10508 17172 10572
rect 17236 10508 17237 10572
rect 17171 10507 17237 10508
rect 16619 9076 16685 9077
rect 16619 9012 16620 9076
rect 16684 9012 16685 9076
rect 16619 9011 16685 9012
rect 16435 6356 16501 6357
rect 16435 6292 16436 6356
rect 16500 6292 16501 6356
rect 16435 6291 16501 6292
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14227 5268 14293 5269
rect 14227 5204 14228 5268
rect 14292 5204 14293 5268
rect 14227 5203 14293 5204
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14043 3908 14109 3909
rect 14043 3844 14044 3908
rect 14108 3844 14109 3908
rect 14043 3843 14109 3844
rect 14672 3840 14992 4864
rect 16622 3909 16682 9011
rect 17174 7717 17234 10507
rect 17542 9621 17602 13635
rect 17726 12613 17786 19075
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18643 18052 18709 18053
rect 18643 17988 18644 18052
rect 18708 17988 18709 18052
rect 18643 17987 18709 17988
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 17907 16828 17973 16829
rect 17907 16764 17908 16828
rect 17972 16764 17973 16828
rect 17907 16763 17973 16764
rect 17723 12612 17789 12613
rect 17723 12548 17724 12612
rect 17788 12548 17789 12612
rect 17723 12547 17789 12548
rect 17539 9620 17605 9621
rect 17539 9556 17540 9620
rect 17604 9556 17605 9620
rect 17539 9555 17605 9556
rect 17539 9348 17605 9349
rect 17539 9284 17540 9348
rect 17604 9284 17605 9348
rect 17539 9283 17605 9284
rect 17723 9348 17789 9349
rect 17723 9284 17724 9348
rect 17788 9284 17789 9348
rect 17723 9283 17789 9284
rect 17171 7716 17237 7717
rect 17171 7652 17172 7716
rect 17236 7652 17237 7716
rect 17171 7651 17237 7652
rect 17171 6492 17237 6493
rect 17171 6428 17172 6492
rect 17236 6428 17237 6492
rect 17171 6427 17237 6428
rect 16619 3908 16685 3909
rect 16619 3844 16620 3908
rect 16684 3844 16685 3908
rect 16619 3843 16685 3844
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 12387 2820 12453 2821
rect 12387 2756 12388 2820
rect 12452 2756 12453 2820
rect 12387 2755 12453 2756
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 2752 14992 3776
rect 17174 3365 17234 6427
rect 17171 3364 17237 3365
rect 17171 3300 17172 3364
rect 17236 3300 17237 3364
rect 17171 3299 17237 3300
rect 17542 3229 17602 9283
rect 17726 5949 17786 9283
rect 17723 5948 17789 5949
rect 17723 5884 17724 5948
rect 17788 5884 17789 5948
rect 17723 5883 17789 5884
rect 17539 3228 17605 3229
rect 17539 3164 17540 3228
rect 17604 3164 17605 3228
rect 17539 3163 17605 3164
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 17910 2685 17970 16763
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18646 8122 18706 17987
rect 19011 17372 19077 17373
rect 19011 17308 19012 17372
rect 19076 17308 19077 17372
rect 19011 17307 19077 17308
rect 18827 17100 18893 17101
rect 18827 17036 18828 17100
rect 18892 17036 18893 17100
rect 18827 17035 18893 17036
rect 18830 14789 18890 17035
rect 19014 15333 19074 17307
rect 19563 16420 19629 16421
rect 19563 16356 19564 16420
rect 19628 16356 19629 16420
rect 19563 16355 19629 16356
rect 19379 16012 19445 16013
rect 19379 15948 19380 16012
rect 19444 15948 19445 16012
rect 19379 15947 19445 15948
rect 19011 15332 19077 15333
rect 19011 15268 19012 15332
rect 19076 15268 19077 15332
rect 19011 15267 19077 15268
rect 19011 14924 19077 14925
rect 19011 14860 19012 14924
rect 19076 14860 19077 14924
rect 19011 14859 19077 14860
rect 18827 14788 18893 14789
rect 18827 14724 18828 14788
rect 18892 14724 18893 14788
rect 18827 14723 18893 14724
rect 18827 14652 18893 14653
rect 18827 14588 18828 14652
rect 18892 14588 18893 14652
rect 18827 14587 18893 14588
rect 18830 12205 18890 14587
rect 19014 13565 19074 14859
rect 19382 14245 19442 15947
rect 19379 14244 19445 14245
rect 19379 14180 19380 14244
rect 19444 14180 19445 14244
rect 19379 14179 19445 14180
rect 19566 13970 19626 16355
rect 19931 14516 19997 14517
rect 19931 14452 19932 14516
rect 19996 14452 19997 14516
rect 19931 14451 19997 14452
rect 19747 14108 19813 14109
rect 19747 14044 19748 14108
rect 19812 14044 19813 14108
rect 19747 14043 19813 14044
rect 19382 13910 19626 13970
rect 19011 13564 19077 13565
rect 19011 13500 19012 13564
rect 19076 13500 19077 13564
rect 19011 13499 19077 13500
rect 19195 12748 19261 12749
rect 19195 12684 19196 12748
rect 19260 12684 19261 12748
rect 19195 12683 19261 12684
rect 19011 12612 19077 12613
rect 19011 12548 19012 12612
rect 19076 12548 19077 12612
rect 19011 12547 19077 12548
rect 18827 12204 18893 12205
rect 18827 12140 18828 12204
rect 18892 12140 18893 12204
rect 18827 12139 18893 12140
rect 19014 11253 19074 12547
rect 19198 12205 19258 12683
rect 19195 12204 19261 12205
rect 19195 12140 19196 12204
rect 19260 12140 19261 12204
rect 19195 12139 19261 12140
rect 19382 12066 19442 13910
rect 19563 13836 19629 13837
rect 19563 13772 19564 13836
rect 19628 13772 19629 13836
rect 19563 13771 19629 13772
rect 19198 12006 19442 12066
rect 18827 11252 18893 11253
rect 18827 11188 18828 11252
rect 18892 11188 18893 11252
rect 18827 11187 18893 11188
rect 19011 11252 19077 11253
rect 19011 11188 19012 11252
rect 19076 11188 19077 11252
rect 19011 11187 19077 11188
rect 18830 9349 18890 11187
rect 18827 9348 18893 9349
rect 18827 9284 18828 9348
rect 18892 9284 18893 9348
rect 18827 9283 18893 9284
rect 19198 9077 19258 12006
rect 19379 11932 19445 11933
rect 19379 11868 19380 11932
rect 19444 11868 19445 11932
rect 19379 11867 19445 11868
rect 19382 9485 19442 11867
rect 19379 9484 19445 9485
rect 19379 9420 19380 9484
rect 19444 9420 19445 9484
rect 19379 9419 19445 9420
rect 19195 9076 19261 9077
rect 19195 9074 19196 9076
rect 19014 9014 19196 9074
rect 18827 8668 18893 8669
rect 18827 8604 18828 8668
rect 18892 8604 18893 8668
rect 18827 8603 18893 8604
rect 18830 8261 18890 8603
rect 18827 8260 18893 8261
rect 18827 8196 18828 8260
rect 18892 8196 18893 8260
rect 18827 8195 18893 8196
rect 18646 8062 18890 8122
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18830 7034 18890 8062
rect 19014 7581 19074 9014
rect 19195 9012 19196 9014
rect 19260 9012 19261 9076
rect 19195 9011 19261 9012
rect 19379 8124 19445 8125
rect 19379 8122 19380 8124
rect 19198 8062 19380 8122
rect 19011 7580 19077 7581
rect 19011 7516 19012 7580
rect 19076 7516 19077 7580
rect 19011 7515 19077 7516
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18646 6974 18890 7034
rect 19011 7036 19077 7037
rect 18646 4045 18706 6974
rect 19011 6972 19012 7036
rect 19076 6972 19077 7036
rect 19011 6971 19077 6972
rect 18827 6900 18893 6901
rect 18827 6836 18828 6900
rect 18892 6836 18893 6900
rect 18827 6835 18893 6836
rect 18643 4044 18709 4045
rect 18643 3980 18644 4044
rect 18708 3980 18709 4044
rect 18643 3979 18709 3980
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 17907 2684 17973 2685
rect 17907 2620 17908 2684
rect 17972 2620 17973 2684
rect 17907 2619 17973 2620
rect 18104 2208 18424 3232
rect 18830 2549 18890 6835
rect 19014 6357 19074 6971
rect 19011 6356 19077 6357
rect 19011 6292 19012 6356
rect 19076 6292 19077 6356
rect 19011 6291 19077 6292
rect 19011 6220 19077 6221
rect 19011 6156 19012 6220
rect 19076 6156 19077 6220
rect 19011 6155 19077 6156
rect 19014 3229 19074 6155
rect 19011 3228 19077 3229
rect 19011 3164 19012 3228
rect 19076 3164 19077 3228
rect 19011 3163 19077 3164
rect 19198 2821 19258 8062
rect 19379 8060 19380 8062
rect 19444 8060 19445 8124
rect 19379 8059 19445 8060
rect 19379 7172 19445 7173
rect 19379 7108 19380 7172
rect 19444 7108 19445 7172
rect 19379 7107 19445 7108
rect 19195 2820 19261 2821
rect 19195 2756 19196 2820
rect 19260 2756 19261 2820
rect 19195 2755 19261 2756
rect 18827 2548 18893 2549
rect 18827 2484 18828 2548
rect 18892 2484 18893 2548
rect 18827 2483 18893 2484
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
rect 7051 2075 7117 2076
rect 19382 917 19442 7107
rect 19566 2413 19626 13771
rect 19750 6901 19810 14043
rect 19934 12477 19994 14451
rect 19931 12476 19997 12477
rect 19931 12412 19932 12476
rect 19996 12412 19997 12476
rect 19931 12411 19997 12412
rect 20115 10436 20181 10437
rect 20115 10372 20116 10436
rect 20180 10372 20181 10436
rect 20115 10371 20181 10372
rect 19931 10164 19997 10165
rect 19931 10100 19932 10164
rect 19996 10100 19997 10164
rect 19931 10099 19997 10100
rect 19934 7581 19994 10099
rect 20118 7989 20178 10371
rect 20115 7988 20181 7989
rect 20115 7924 20116 7988
rect 20180 7924 20181 7988
rect 20115 7923 20181 7924
rect 19931 7580 19997 7581
rect 19931 7516 19932 7580
rect 19996 7516 19997 7580
rect 19931 7515 19997 7516
rect 19747 6900 19813 6901
rect 19747 6836 19748 6900
rect 19812 6836 19813 6900
rect 19747 6835 19813 6836
rect 19747 5404 19813 5405
rect 19747 5340 19748 5404
rect 19812 5340 19813 5404
rect 19747 5339 19813 5340
rect 19563 2412 19629 2413
rect 19563 2348 19564 2412
rect 19628 2348 19629 2412
rect 19563 2347 19629 2348
rect 19750 2277 19810 5339
rect 19747 2276 19813 2277
rect 19747 2212 19748 2276
rect 19812 2212 19813 2276
rect 19747 2211 19813 2212
rect 19379 916 19445 917
rect 19379 852 19380 916
rect 19444 852 19445 916
rect 19379 851 19445 852
use sky130_fd_sc_hd__decap_3  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1932 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1606821651
transform 1 0 1656 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18
timestamp 1606821651
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1606821651
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3864 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1606821651
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1606821651
transform 1 0 5796 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1606821651
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48
timestamp 1606821651
transform 1 0 5520 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1606821651
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1606821651
transform 1 0 5336 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1606821651
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8464 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1606821651
transform 1 0 7912 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1606821651
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1606821651
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_78
timestamp 1606821651
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 9108 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _145_
timestamp 1606821651
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 10672 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1606821651
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1606821651
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_96
timestamp 1606821651
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1606821651
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1606821651
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10764 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_123
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1606821651
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1606821651
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 11776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1606821651
transform 1 0 12604 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13800 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1606821651
transform 1 0 13340 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1606821651
transform 1 0 14352 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1606821651
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_142
timestamp 1606821651
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_134
timestamp 1606821651
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1606821651
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1606821651
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 14812 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_164
timestamp 1606821651
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_162
timestamp 1606821651
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1606821651
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1606821651
transform 1 0 16192 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606821651
transform 1 0 15824 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1606821651
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1606821651
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1606821651
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1606821651
transform 1 0 17204 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1606821651
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606821651
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1606821651
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1606821651
transform 1 0 18216 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606821651
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1606821651
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1606821651
transform 1 0 19412 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 19320 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1606821651
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_207
timestamp 1606821651
transform 1 0 20148 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1606821651
transform 1 0 19044 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_208
timestamp 1606821651
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1606821651
transform 1 0 20424 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_S_FTB01
timestamp 1606821651
transform 1 0 20332 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1606821651
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606821651
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_216
timestamp 1606821651
transform 1 0 20976 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _051_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1472 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1932 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1606821651
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4416 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1606821651
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_25
timestamp 1606821651
transform 1 0 3404 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1606821651
transform 1 0 6624 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5428 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1606821651
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_56
timestamp 1606821651
transform 1 0 6256 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1606821651
transform 1 0 7636 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_69
timestamp 1606821651
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1606821651
transform 1 0 8464 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 8832 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1606821651
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_102
timestamp 1606821651
transform 1 0 10488 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10764 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1606821651
transform 1 0 12420 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_121
timestamp 1606821651
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14444 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1606821651
transform 1 0 13432 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_132
timestamp 1606821651
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_143
timestamp 1606821651
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15824 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1606821651
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_158
timestamp 1606821651
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606821651
transform 1 0 17480 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 18032 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_176
timestamp 1606821651
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1606821651
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606821651
transform 1 0 20148 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1606821651
transform 1 0 19136 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp 1606821651
transform 1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_205
timestamp 1606821651
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606821651
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_211
timestamp 1606821651
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_218
timestamp 1606821651
transform 1 0 21160 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2852 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1840 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_6
timestamp 1606821651
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1606821651
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4876 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1606821651
transform 1 0 3864 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_28
timestamp 1606821651
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_39
timestamp 1606821651
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1606821651
transform 1 0 6164 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_50
timestamp 1606821651
transform 1 0 5704 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_54
timestamp 1606821651
transform 1 0 6072 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606821651
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1606821651
transform 1 0 8004 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8556 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1606821651
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_79
timestamp 1606821651
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 10212 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_97
timestamp 1606821651
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606821651
transform 1 0 12512 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_105
timestamp 1606821651
transform 1 0 10764 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1606821651
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13064 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_128
timestamp 1606821651
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 14720 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1606821651
transform 1 0 15732 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_146
timestamp 1606821651
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1606821651
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 18032 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16744 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_168
timestamp 1606821651
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1606821651
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1606821651
transform 1 0 19688 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1606821651
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _138_
timestamp 1606821651
transform 1 0 20700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1606821651
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 1606821651
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1472 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_20
timestamp 1606821651
transform 1 0 2944 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1606821651
transform 1 0 3404 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_24
timestamp 1606821651
transform 1 0 3312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1606821651
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 1606821651
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1606821651
transform 1 0 5060 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 5612 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_47
timestamp 1606821651
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8280 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 7268 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_65
timestamp 1606821651
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_76
timestamp 1606821651
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606821651
transform 1 0 9844 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1606821651
transform 1 0 10396 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1606821651
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1606821651
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_99
timestamp 1606821651
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12420 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11408 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_110
timestamp 1606821651
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_121
timestamp 1606821651
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13432 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_132
timestamp 1606821651
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_143
timestamp 1606821651
transform 1 0 14260 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606821651
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 16284 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1606821651
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1606821651
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 17112 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_4_171
timestamp 1606821651
transform 1 0 16836 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  clk_2_S_FTB01
timestamp 1606821651
transform 1 0 20056 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1606821651
transform 1 0 19044 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_190
timestamp 1606821651
transform 1 0 18584 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_194
timestamp 1606821651
transform 1 0 18952 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_204
timestamp 1606821651
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1606821651
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1606821651
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_218
timestamp 1606821651
transform 1 0 21160 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1606821651
transform 1 0 2116 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_9
timestamp 1606821651
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_20
timestamp 1606821651
transform 1 0 2944 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1606821651
transform 1 0 4324 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1606821651
transform 1 0 3312 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_33
timestamp 1606821651
transform 1 0 4140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1606821651
transform 1 0 5704 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_44
timestamp 1606821651
transform 1 0 5152 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606821651
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8740 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1606821651
transform 1 0 8280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_82
timestamp 1606821651
transform 1 0 8648 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606821651
transform 1 0 10396 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_99
timestamp 1606821651
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10948 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_105
timestamp 1606821651
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_116
timestamp 1606821651
transform 1 0 11776 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13616 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606821651
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1606821651
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_145
timestamp 1606821651
transform 1 0 14444 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15732 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1606821651
transform 1 0 14720 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_157
timestamp 1606821651
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606821651
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_3_S_FTB01
timestamp 1606821651
transform 1 0 18032 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1606821651
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1606821651
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 18768 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_190
timestamp 1606821651
transform 1 0 18584 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_208
timestamp 1606821651
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 20424 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_216
timestamp 1606821651
transform 1 0 20976 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606821651
transform 1 0 1748 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 1932 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2208 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_10
timestamp 1606821651
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1606821651
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1606821651
transform 1 0 4692 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1606821651
transform 1 0 3588 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_28
timestamp 1606821651
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_25
timestamp 1606821651
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_36
timestamp 1606821651
transform 1 0 4416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 1606821651
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1606821651
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5244 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606821651
transform 1 0 5704 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606821651
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1606821651
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_53
timestamp 1606821651
transform 1 0 5980 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1606821651
transform 1 0 6164 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606821651
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_68
timestamp 1606821651
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_64
timestamp 1606821651
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1606821651
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1606821651
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7728 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1606821651
transform 1 0 6992 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_81
timestamp 1606821651
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_75
timestamp 1606821651
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1606821651
transform 1 0 8188 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1606821651
transform 1 0 8740 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9752 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_86
timestamp 1606821651
transform 1 0 9016 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1606821651
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_110
timestamp 1606821651
transform 1 0 11224 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1606821651
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1606821651
transform 1 0 11316 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1606821651
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_120
timestamp 1606821651
transform 1 0 12144 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1606821651
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1606821651
transform 1 0 12512 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 12604 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _148_
timestamp 1606821651
transform 1 0 14444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13064 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1606821651
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_141
timestamp 1606821651
transform 1 0 14076 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606821651
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 14996 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 15456 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1606821651
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1606821651
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_165
timestamp 1606821651
transform 1 0 16284 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_149
timestamp 1606821651
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 16652 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 18124 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_167
timestamp 1606821651
transform 1 0 16468 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_171
timestamp 1606821651
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606821651
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19320 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1606821651
transform 1 0 19320 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1606821651
transform 1 0 19136 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1606821651
transform 1 0 18952 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_207
timestamp 1606821651
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1606821651
transform 1 0 18860 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_197
timestamp 1606821651
transform 1 0 19228 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1606821651
transform 1 0 20332 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1606821651
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606821651
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606821651
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_214
timestamp 1606821651
transform 1 0 20792 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1606821651
transform 1 0 1564 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1606821651
transform 1 0 2116 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_9
timestamp 1606821651
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_20
timestamp 1606821651
transform 1 0 2944 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1606821651
transform 1 0 3404 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_24
timestamp 1606821651
transform 1 0 3312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1606821651
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1606821651
transform 1 0 4876 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1606821651
transform 1 0 5244 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1606821651
transform 1 0 6072 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1606821651
transform 1 0 8556 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1606821651
transform 1 0 7268 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8280 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1606821651
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_63
timestamp 1606821651
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_76
timestamp 1606821651
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1606821651
transform 1 0 9844 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1606821651
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_104
timestamp 1606821651
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10856 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11868 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_115
timestamp 1606821651
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1606821651
transform 1 0 13892 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_126
timestamp 1606821651
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_137
timestamp 1606821651
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _141_
timestamp 1606821651
transform 1 0 16284 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1606821651
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1606821651
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1606821651
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 17848 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 16836 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_169
timestamp 1606821651
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_180
timestamp 1606821651
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 19136 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_191
timestamp 1606821651
transform 1 0 18676 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1606821651
transform 1 0 19044 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606821651
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1606821651
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_218
timestamp 1606821651
transform 1 0 21160 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1748 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 3772 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_9_23
timestamp 1606821651
transform 1 0 3220 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5428 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_45
timestamp 1606821651
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_56
timestamp 1606821651
transform 1 0 6256 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1606821651
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_62
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7084 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp 1606821651
transform 1 0 8556 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9844 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8832 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1606821651
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_104
timestamp 1606821651
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1606821651
transform 1 0 11868 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10856 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_115
timestamp 1606821651
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1606821651
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1606821651
transform 1 0 14076 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_139
timestamp 1606821651
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1606821651
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15364 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_150
timestamp 1606821651
transform 1 0 14904 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_154
timestamp 1606821651
transform 1 0 15272 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_164
timestamp 1606821651
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606821651
transform 1 0 17388 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1606821651
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1606821651
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1606821651
transform 1 0 19044 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1606821651
transform 1 0 20056 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1606821651
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_204
timestamp 1606821651
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1606821651
transform 1 0 20884 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1606821651
transform 1 0 21252 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2300 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1606821651
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1606821651
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1606821651
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1606821651
transform 1 0 6348 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 5060 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 6072 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1606821651
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_61
timestamp 1606821651
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7912 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6900 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_72
timestamp 1606821651
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1606821651
transform 1 0 9936 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10580 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606821651
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_93
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_100
timestamp 1606821651
transform 1 0 10304 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1606821651
transform 1 0 12236 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_119
timestamp 1606821651
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13524 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 13248 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_130
timestamp 1606821651
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 16284 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606821651
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_163
timestamp 1606821651
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606821651
transform 1 0 16560 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 17112 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_172
timestamp 1606821651
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1606821651
transform 1 0 19780 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1606821651
transform 1 0 18584 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1606821651
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_199
timestamp 1606821651
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1606821651
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606821651
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606821651
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1606821651
transform 1 0 2392 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_12
timestamp 1606821651
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606821651
transform 1 0 3404 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3956 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_23
timestamp 1606821651
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_29
timestamp 1606821651
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_47
timestamp 1606821651
transform 1 0 5428 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606821651
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1606821651
transform 1 0 8464 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1606821651
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10488 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1606821651
transform 1 0 9476 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_89
timestamp 1606821651
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_100
timestamp 1606821651
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1606821651
transform 1 0 11776 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_111
timestamp 1606821651
transform 1 0 11316 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_115
timestamp 1606821651
transform 1 0 11684 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606821651
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14444 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1606821651
transform 1 0 13432 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1606821651
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_143
timestamp 1606821651
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _147_
timestamp 1606821651
transform 1 0 15548 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16100 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_154
timestamp 1606821651
transform 1 0 15272 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_161
timestamp 1606821651
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1606821651
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1606821651
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1606821651
transform 1 0 20056 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1606821651
transform 1 0 19044 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1606821651
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_204
timestamp 1606821651
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1606821651
transform 1 0 20884 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_219
timestamp 1606821651
transform 1 0 21252 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1606821651
transform 1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1606821651
transform 1 0 1932 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1606821651
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_18
timestamp 1606821651
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1606821651
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1606821651
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1606821651
transform 1 0 6808 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5060 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_12_59
timestamp 1606821651
transform 1 0 6532 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7360 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_66
timestamp 1606821651
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1606821651
transform 1 0 10580 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1606821651
transform 1 0 9016 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1606821651
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1606821651
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_102
timestamp 1606821651
transform 1 0 10488 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 10948 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1606821651
transform 1 0 12604 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_123
timestamp 1606821651
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1606821651
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_134
timestamp 1606821651
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_145
timestamp 1606821651
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1606821651
transform 1 0 14628 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16284 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1606821651
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1606821651
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 18308 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1606821651
transform 1 0 17296 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_174
timestamp 1606821651
transform 1 0 17112 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_185
timestamp 1606821651
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19964 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_203
timestamp 1606821651
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606821651
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1606821651
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_218
timestamp 1606821651
transform 1 0 21160 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_8
timestamp 1606821651
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1606821651
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606821651
transform 1 0 1564 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606821651
transform 1 0 1472 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_19
timestamp 1606821651
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1606821651
transform 1 0 2024 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1606821651
transform 1 0 2116 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_20
timestamp 1606821651
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606821651
transform 1 0 3036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1606821651
transform 1 0 3128 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1606821651
transform 1 0 4140 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_31
timestamp 1606821651
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_25
timestamp 1606821651
transform 1 0 3404 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_48
timestamp 1606821651
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_42
timestamp 1606821651
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1606821651
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1606821651
transform 1 0 5704 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606821651
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1606821651
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6532 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _149_
timestamp 1606821651
transform 1 0 6164 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 7820 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1606821651
transform 1 0 7728 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 8740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1606821651
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1606821651
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_68
timestamp 1606821651
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_81
timestamp 1606821651
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1606821651
transform 1 0 9016 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10488 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1606821651
transform 1 0 9476 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_89
timestamp 1606821651
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_100
timestamp 1606821651
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606821651
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1606821651
transform 1 0 11408 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12420 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1606821651
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_109
timestamp 1606821651
transform 1 0 11132 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_121
timestamp 1606821651
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1606821651
transform 1 0 13432 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 14352 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_139
timestamp 1606821651
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_132
timestamp 1606821651
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_143
timestamp 1606821651
transform 1 0 14260 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606821651
transform 1 0 14628 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15732 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_153
timestamp 1606821651
transform 1 0 15180 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1606821651
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_170
timestamp 1606821651
transform 1 0 16744 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1606821651
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1606821651
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1606821651
transform 1 0 17296 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_185
timestamp 1606821651
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1606821651
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1606821651
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606821651
transform 1 0 17388 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18308 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606821651
transform 1 0 19044 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1606821651
transform 1 0 20056 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1606821651
transform 1 0 19044 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1606821651
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1606821651
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_193
timestamp 1606821651
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1606821651
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1606821651
transform 1 0 20884 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1606821651
transform 1 0 21252 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1606821651
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_218
timestamp 1606821651
transform 1 0 21160 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1840 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_6
timestamp 1606821651
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1606821651
transform 1 0 3496 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4416 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1606821651
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_30
timestamp 1606821651
transform 1 0 3864 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5428 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_45
timestamp 1606821651
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_56
timestamp 1606821651
transform 1 0 6256 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1606821651
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 7820 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1606821651
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_82
timestamp 1606821651
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1606821651
transform 1 0 9108 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 8832 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_91
timestamp 1606821651
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606821651
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1606821651
transform 1 0 13432 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1606821651
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_143
timestamp 1606821651
transform 1 0 14260 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1606821651
transform 1 0 14720 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15916 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_147
timestamp 1606821651
transform 1 0 14628 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_157
timestamp 1606821651
transform 1 0 15548 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18124 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1606821651
transform 1 0 16928 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_170
timestamp 1606821651
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1606821651
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_184
timestamp 1606821651
transform 1 0 18032 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1606821651
transform 1 0 19780 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_201
timestamp 1606821651
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606821651
transform 1 0 20792 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1606821651
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1606821651
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606821651
transform 1 0 1840 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_6
timestamp 1606821651
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1606821651
transform 1 0 3496 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_24
timestamp 1606821651
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1606821651
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1606821651
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606821651
transform 1 0 5060 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 5796 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_47
timestamp 1606821651
transform 1 0 5428 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7452 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_67
timestamp 1606821651
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606821651
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1606821651
transform 1 0 9936 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10488 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1606821651
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606821651
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_100
timestamp 1606821651
transform 1 0 10304 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12420 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_122
timestamp 1606821651
transform 1 0 12328 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1606821651
transform 1 0 14076 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_139
timestamp 1606821651
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1606821651
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1606821651
transform 1 0 16100 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16560 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1606821651
transform 1 0 17572 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_167
timestamp 1606821651
transform 1 0 16468 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_177
timestamp 1606821651
transform 1 0 17388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1606821651
transform 1 0 18584 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19136 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_188
timestamp 1606821651
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1606821651
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1606821651
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1606821651
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_218
timestamp 1606821651
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1606821651
transform 1 0 2208 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1472 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_10
timestamp 1606821651
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606821651
transform 1 0 4784 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3312 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_21
timestamp 1606821651
transform 1 0 3036 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1606821651
transform 1 0 5520 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1606821651
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_44
timestamp 1606821651
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1606821651
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1606821651
transform 1 0 7820 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1606821651
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_82
timestamp 1606821651
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 10580 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1606821651
transform 1 0 9660 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1606821651
transform 1 0 8832 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_102
timestamp 1606821651
transform 1 0 10488 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_119
timestamp 1606821651
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 14352 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 14076 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1606821651
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16284 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_160
timestamp 1606821651
transform 1 0 15824 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_164
timestamp 1606821651
transform 1 0 16192 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606821651
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606821651
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1606821651
transform 1 0 19780 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1606821651
transform 1 0 18768 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_190
timestamp 1606821651
transform 1 0 18584 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_201
timestamp 1606821651
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606821651
transform 1 0 20792 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1606821651
transform 1 0 20608 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1606821651
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1606821651
transform 1 0 1932 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1606821651
transform 1 0 2944 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_7
timestamp 1606821651
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_18
timestamp 1606821651
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4692 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1606821651
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_36
timestamp 1606821651
transform 1 0 4416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6348 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_55
timestamp 1606821651
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1606821651
transform 1 0 8372 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1606821651
transform 1 0 7360 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_66
timestamp 1606821651
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 1606821651
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 9844 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1606821651
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11500 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_111
timestamp 1606821651
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_122
timestamp 1606821651
transform 1 0 12328 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1606821651
transform 1 0 12696 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1606821651
transform 1 0 13708 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_135
timestamp 1606821651
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606821651
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15456 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_146
timestamp 1606821651
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1606821651
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_165
timestamp 1606821651
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 16468 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 18124 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_183
timestamp 1606821651
transform 1 0 17940 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1606821651
transform 1 0 19780 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_201
timestamp 1606821651
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606821651
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606821651
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1606821651
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_218
timestamp 1606821651
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1564 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1606821651
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_14
timestamp 1606821651
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2300 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2576 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1606821651
transform 1 0 4232 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4140 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_32
timestamp 1606821651
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1606821651
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_32
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_42
timestamp 1606821651
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_43
timestamp 1606821651
transform 1 0 5060 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5152 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5428 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_58
timestamp 1606821651
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_53
timestamp 1606821651
transform 1 0 5980 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_56
timestamp 1606821651
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1606821651
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1606821651
transform 1 0 6072 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 6808 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7268 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7820 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1606821651
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_83
timestamp 1606821651
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_71
timestamp 1606821651
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1606821651
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _146_
timestamp 1606821651
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1606821651
transform 1 0 9936 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8924 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10672 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_94
timestamp 1606821651
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1606821651
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1606821651
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1606821651
transform 1 0 10948 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1606821651
transform 1 0 11684 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_105
timestamp 1606821651
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_116
timestamp 1606821651
transform 1 0 11776 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_123
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_113
timestamp 1606821651
transform 1 0 11500 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_124
timestamp 1606821651
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606821651
transform 1 0 12972 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13524 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12696 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14352 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 12696 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_142
timestamp 1606821651
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 1606821651
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1606821651
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_153
timestamp 1606821651
transform 1 0 15180 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 15364 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_163
timestamp 1606821651
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1606821651
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1606821651
transform 1 0 16192 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606821651
transform 1 0 15640 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1606821651
transform 1 0 16376 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1606821651
transform 1 0 17388 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1606821651
transform 1 0 18308 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1606821651
transform 1 0 18216 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 17204 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606821651
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp 1606821651
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1606821651
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_184
timestamp 1606821651
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_175
timestamp 1606821651
transform 1 0 17204 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1606821651
transform 1 0 19412 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1606821651
transform 1 0 19320 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1606821651
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_196
timestamp 1606821651
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1606821651
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_195
timestamp 1606821651
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_208
timestamp 1606821651
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1606821651
transform 1 0 20332 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606821651
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_218
timestamp 1606821651
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606821651
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606821651
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1606821651
transform 1 0 1932 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2944 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1606821651
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_18
timestamp 1606821651
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3956 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1606821651
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5612 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_47
timestamp 1606821651
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_58
timestamp 1606821651
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7820 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1606821651
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _144_
timestamp 1606821651
transform 1 0 9568 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10120 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_89
timestamp 1606821651
transform 1 0 9292 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_96
timestamp 1606821651
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11132 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_107
timestamp 1606821651
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1606821651
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_123
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 12696 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_142
timestamp 1606821651
transform 1 0 14168 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606821651
transform 1 0 14536 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15088 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_150
timestamp 1606821651
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18032 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16744 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606821651
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_168
timestamp 1606821651
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1606821651
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 19688 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1606821651
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606821651
transform 1 0 20700 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1606821651
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_217
timestamp 1606821651
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1606821651
transform 1 0 1840 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2852 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_6
timestamp 1606821651
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_17
timestamp 1606821651
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_28
timestamp 1606821651
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1606821651
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5888 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 5060 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_49
timestamp 1606821651
transform 1 0 5612 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1606821651
transform 1 0 7544 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 8556 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_68
timestamp 1606821651
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_79
timestamp 1606821651
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9936 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606821651
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1606821651
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1606821651
transform 1 0 10948 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1606821651
transform 1 0 11960 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_105
timestamp 1606821651
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1606821651
transform 1 0 11776 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13984 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12972 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_127
timestamp 1606821651
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1606821651
transform 1 0 13800 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1606821651
transform 1 0 16008 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15272 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606821651
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1606821651
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_160
timestamp 1606821651
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 17020 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_171
timestamp 1606821651
transform 1 0 16836 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1606821651
transform 1 0 18676 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1606821651
transform 1 0 19688 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_189
timestamp 1606821651
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_200
timestamp 1606821651
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1606821651
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606821651
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1606821651
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1606821651
transform 1 0 21160 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1748 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1606821651
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 3404 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1606821651
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_41
timestamp 1606821651
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5060 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606821651
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606821651
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1606821651
transform 1 0 7820 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8740 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1606821651
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_77
timestamp 1606821651
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_82
timestamp 1606821651
transform 1 0 8648 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 10396 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_99
timestamp 1606821651
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606821651
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_117
timestamp 1606821651
transform 1 0 11868 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606821651
transform 1 0 13616 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 14168 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_132
timestamp 1606821651
transform 1 0 13248 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_140
timestamp 1606821651
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 16192 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_23_158
timestamp 1606821651
transform 1 0 15640 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606821651
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1606821651
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1606821651
transform 1 0 19044 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1606821651
transform 1 0 20056 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_193
timestamp 1606821651
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_204
timestamp 1606821651
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1606821651
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1606821651
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1606821651
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2944 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1606821651
transform 1 0 1932 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1606821651
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_18
timestamp 1606821651
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4232 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606821651
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1606821651
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1606821651
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5336 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 6532 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_43
timestamp 1606821651
transform 1 0 5060 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_55
timestamp 1606821651
transform 1 0 6164 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7544 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 8556 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_68
timestamp 1606821651
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_79
timestamp 1606821651
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 10028 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606821651
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1606821651
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1606821651
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11224 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_106
timestamp 1606821651
transform 1 0 10856 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12880 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_126
timestamp 1606821651
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_144
timestamp 1606821651
transform 1 0 14352 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606821651
transform 1 0 14628 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1606821651
transform 1 0 16284 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1606821651
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606821651
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606821651
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1606821651
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1606821651
transform 1 0 17296 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18308 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_174
timestamp 1606821651
transform 1 0 17112 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_185
timestamp 1606821651
transform 1 0 18124 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1606821651
transform 1 0 19320 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_196
timestamp 1606821651
transform 1 0 19136 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_207
timestamp 1606821651
transform 1 0 20148 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606821651
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1606821651
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606821651
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606821651
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1606821651
transform 1 0 1472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2024 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1606821651
transform 1 0 2760 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1606821651
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_8
timestamp 1606821651
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_16
timestamp 1606821651
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1606821651
transform 1 0 4784 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1606821651
transform 1 0 3772 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_27
timestamp 1606821651
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1606821651
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1606821651
transform 1 0 5796 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606821651
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 6348 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_49
timestamp 1606821651
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_55
timestamp 1606821651
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1606821651
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1606821651
transform 1 0 8464 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1606821651
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10488 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1606821651
transform 1 0 9476 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_89
timestamp 1606821651
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1606821651
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606821651
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1606821651
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13432 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1606821651
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_143
timestamp 1606821651
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15548 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1606821651
transform 1 0 14536 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1606821651
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1606821651
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1606821651
transform 1 0 16560 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606821651
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_177
timestamp 1606821651
transform 1 0 17388 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 19044 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1606821651
transform 1 0 20056 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1606821651
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_204
timestamp 1606821651
transform 1 0 19872 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1606821651
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1606821651
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2116 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1380 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1606821651
transform 1 0 2576 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1606821651
transform 1 0 1564 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1606821651
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_14
timestamp 1606821651
transform 1 0 2392 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1606821651
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606821651
transform 1 0 3772 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1606821651
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1606821651
transform 1 0 4232 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606821651
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_25
timestamp 1606821651
transform 1 0 3404 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 1606821651
transform 1 0 4876 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_27
timestamp 1606821651
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_32
timestamp 1606821651
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606821651
transform 1 0 5244 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5244 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606821651
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_61
timestamp 1606821651
transform 1 0 6716 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_43
timestamp 1606821651
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_48
timestamp 1606821651
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1606821651
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_62
timestamp 1606821651
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 6900 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7912 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 6900 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_72
timestamp 1606821651
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_79
timestamp 1606821651
transform 1 0 8372 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_83
timestamp 1606821651
transform 1 0 8740 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_88
timestamp 1606821651
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1606821651
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1606821651
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606821651
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1606821651
transform 1 0 9384 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _135_
timestamp 1606821651
transform 1 0 8832 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1606821651
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_100
timestamp 1606821651
transform 1 0 10304 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10396 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1606821651
transform 1 0 9936 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10488 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _131_
timestamp 1606821651
transform 1 0 11408 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _132_
timestamp 1606821651
transform 1 0 12144 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606821651
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_118
timestamp 1606821651
transform 1 0 11960 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_124
timestamp 1606821651
transform 1 0 12512 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1606821651
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_116
timestamp 1606821651
transform 1 0 11776 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13800 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12972 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_26_128
timestamp 1606821651
transform 1 0 12880 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1606821651
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_132
timestamp 1606821651
transform 1 0 13248 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _143_
timestamp 1606821651
transform 1 0 14628 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15456 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1606821651
transform 1 0 16284 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606821651
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1606821651
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1606821651
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_154
timestamp 1606821651
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_176
timestamp 1606821651
transform 1 0 17296 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_172
timestamp 1606821651
transform 1 0 16928 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_174
timestamp 1606821651
transform 1 0 17112 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1606821651
transform 1 0 17296 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1606821651
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_185
timestamp 1606821651
transform 1 0 18124 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606821651
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606821651
transform 1 0 17388 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1606821651
transform 1 0 18308 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1606821651
transform 1 0 20240 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1606821651
transform 1 0 19044 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 19412 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_26_196
timestamp 1606821651
transform 1 0 19136 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_208
timestamp 1606821651
transform 1 0 20240 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1606821651
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_204
timestamp 1606821651
transform 1 0 19872 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606821651
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606821651
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606821651
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_217
timestamp 1606821651
transform 1 0 21068 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 1380 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1606821651
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606821651
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_12
timestamp 1606821651
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1606821651
transform 1 0 3404 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606821651
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1606821651
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1606821651
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1606821651
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6440 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1606821651
transform 1 0 5060 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_28_52
timestamp 1606821651
transform 1 0 5888 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 7452 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1606821651
transform 1 0 8556 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_67
timestamp 1606821651
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_78
timestamp 1606821651
transform 1 0 8280 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10672 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606821651
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1606821651
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1606821651
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1606821651
transform 1 0 11776 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_28_113
timestamp 1606821651
transform 1 0 11500 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_125
timestamp 1606821651
transform 1 0 12604 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _129_
timestamp 1606821651
transform 1 0 12880 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _142_
timestamp 1606821651
transform 1 0 14444 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13432 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_132
timestamp 1606821651
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_143
timestamp 1606821651
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1606821651
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 15732 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606821651
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1606821651
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_157
timestamp 1606821651
transform 1 0 15548 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1606821651
transform 1 0 17388 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_175
timestamp 1606821651
transform 1 0 17204 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_186
timestamp 1606821651
transform 1 0 18216 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1606821651
transform 1 0 19780 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1606821651
transform 1 0 18768 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_201
timestamp 1606821651
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606821651
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606821651
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1606821651
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606821651
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606821651
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1606821651
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2392 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606821651
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1606821651
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_11
timestamp 1606821651
transform 1 0 2116 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4048 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_30
timestamp 1606821651
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_41
timestamp 1606821651
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _139_
timestamp 1606821651
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5060 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606821651
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606821651
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8464 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1606821651
transform 1 0 7452 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_66
timestamp 1606821651
transform 1 0 7176 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1606821651
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10672 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1606821651
transform 1 0 9476 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_89
timestamp 1606821651
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_100
timestamp 1606821651
transform 1 0 10304 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606821651
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1606821651
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13432 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1606821651
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_143
timestamp 1606821651
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _136_
timestamp 1606821651
transform 1 0 14536 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1606821651
transform 1 0 16100 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1606821651
transform 1 0 15088 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_150
timestamp 1606821651
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_161
timestamp 1606821651
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606821651
transform 1 0 17388 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606821651
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606821651
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_172
timestamp 1606821651
transform 1 0 16928 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_176
timestamp 1606821651
transform 1 0 17296 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1606821651
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_184
timestamp 1606821651
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01
timestamp 1606821651
transform 1 0 18492 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19320 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 20056 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_195
timestamp 1606821651
transform 1 0 19044 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_204
timestamp 1606821651
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606821651
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1606821651
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1606821651
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1606821651
transform 1 0 2392 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_2_W_FTB01
timestamp 1606821651
transform 1 0 1656 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606821651
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1606821651
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1606821651
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1606821651
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606821651
transform 1 0 4048 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606821651
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1606821651
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 6716 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5704 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_48
timestamp 1606821651
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1606821651
transform 1 0 6532 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7452 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_67
timestamp 1606821651
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606821651
transform 1 0 9108 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 10672 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606821651
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1606821651
transform 1 0 8924 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1606821651
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1606821651
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 11408 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_110
timestamp 1606821651
transform 1 0 11224 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13064 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_128
timestamp 1606821651
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606821651
transform 1 0 14720 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16284 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606821651
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1606821651
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_146
timestamp 1606821651
transform 1 0 14536 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1606821651
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_154 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 15272 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_162
timestamp 1606821651
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606821651
transform 1 0 17296 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_W_FTB01
timestamp 1606821651
transform 1 0 17848 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_174
timestamp 1606821651
transform 1 0 17112 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_180
timestamp 1606821651
transform 1 0 17664 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  clk_1_W_FTB01
timestamp 1606821651
transform 1 0 18584 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01
timestamp 1606821651
transform 1 0 20056 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1606821651
transform 1 0 19320 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_188
timestamp 1606821651
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_196
timestamp 1606821651
transform 1 0 19136 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_204
timestamp 1606821651
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606821651
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606821651
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1606821651
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606821651
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606821651
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2484 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1606821651
transform 1 0 1656 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606821651
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1606821651
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_12
timestamp 1606821651
transform 1 0 2208 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4784 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 3772 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_24
timestamp 1606821651
transform 1 0 3312 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_28
timestamp 1606821651
transform 1 0 3680 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_38
timestamp 1606821651
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606821651
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_56
timestamp 1606821651
transform 1 0 6256 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1606821651
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1606821651
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 6992 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_80
timestamp 1606821651
transform 1 0 8464 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8832 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 10488 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_100
timestamp 1606821651
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1606821651
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606821651
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_108
timestamp 1606821651
transform 1 0 11040 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1606821651
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13616 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_132
timestamp 1606821651
transform 1 0 13248 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1606821651
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1606821651
transform 1 0 14628 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1606821651
transform 1 0 15456 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_165
timestamp 1606821651
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606821651
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_2_E_FTB01
timestamp 1606821651
transform 1 0 17204 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_E_FTB01
timestamp 1606821651
transform 1 0 16468 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606821651
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_173
timestamp 1606821651
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1606821651
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606821651
transform 1 0 19872 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 18584 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_188
timestamp 1606821651
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_202
timestamp 1606821651
transform 1 0 19688 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_208
timestamp 1606821651
transform 1 0 20240 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_E_FTB01
timestamp 1606821651
transform 1 0 20424 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606821651
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_216
timestamp 1606821651
transform 1 0 20976 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_3_W_FTB01
timestamp 1606821651
transform 1 0 2392 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_W_FTB01
timestamp 1606821651
transform 1 0 1656 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606821651
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1606821651
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_12
timestamp 1606821651
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_20
timestamp 1606821651
transform 1 0 2944 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _133_
timestamp 1606821651
transform 1 0 3404 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606821651
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_24
timestamp 1606821651
transform 1 0 3312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1606821651
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_41
timestamp 1606821651
transform 1 0 4876 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5060 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 6072 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606821651
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_52
timestamp 1606821651
transform 1 0 5888 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_60
timestamp 1606821651
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6900 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_79
timestamp 1606821651
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9752 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606821651
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_90
timestamp 1606821651
transform 1 0 9384 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_103
timestamp 1606821651
transform 1 0 10580 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _130_
timestamp 1606821651
transform 1 0 10948 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1606821651
transform 1 0 11500 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12604 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606821651
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_111
timestamp 1606821651
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1606821651
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _127_
timestamp 1606821651
transform 1 0 13340 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _128_
timestamp 1606821651
transform 1 0 13892 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14444 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_131
timestamp 1606821651
transform 1 0 13156 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_137
timestamp 1606821651
transform 1 0 13708 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_143
timestamp 1606821651
transform 1 0 14260 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _137_
timestamp 1606821651
transform 1 0 16192 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _140_
timestamp 1606821651
transform 1 0 14996 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15640 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606821651
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_156
timestamp 1606821651
transform 1 0 15456 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606821651
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_2_N_FTB01
timestamp 1606821651
transform 1 0 17480 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1606821651
transform 1 0 16744 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606821651
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_168
timestamp 1606821651
transform 1 0 16560 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_176
timestamp 1606821651
transform 1 0 17296 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1606821651
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  clk_1_E_FTB01
timestamp 1606821651
transform 1 0 18860 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1606821651
transform 1 0 19596 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp 1606821651
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_199
timestamp 1606821651
transform 1 0 19412 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_207
timestamp 1606821651
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_E_FTB01
timestamp 1606821651
transform 1 0 20332 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606821651
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606821651
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1606821651
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606821651
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 18418 22320 18474 22800 6 Test_en_N_out
port 0 nsew default tristate
rlabel metal2 s 18878 0 18934 480 6 Test_en_S_in
port 1 nsew default input
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 2 nsew default input
rlabel metal2 s 570 0 626 480 6 bottom_left_grid_pin_43_
port 3 nsew default input
rlabel metal2 s 938 0 994 480 6 bottom_left_grid_pin_44_
port 4 nsew default input
rlabel metal2 s 1306 0 1362 480 6 bottom_left_grid_pin_45_
port 5 nsew default input
rlabel metal2 s 1674 0 1730 480 6 bottom_left_grid_pin_46_
port 6 nsew default input
rlabel metal2 s 2042 0 2098 480 6 bottom_left_grid_pin_47_
port 7 nsew default input
rlabel metal2 s 2410 0 2466 480 6 bottom_left_grid_pin_48_
port 8 nsew default input
rlabel metal2 s 2778 0 2834 480 6 bottom_left_grid_pin_49_
port 9 nsew default input
rlabel metal2 s 3146 0 3202 480 6 ccff_head
port 10 nsew default input
rlabel metal2 s 3514 0 3570 480 6 ccff_tail
port 11 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_in[0]
port 12 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[10]
port 13 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[11]
port 14 nsew default input
rlabel metal3 s 0 7896 480 8016 6 chanx_left_in[12]
port 15 nsew default input
rlabel metal3 s 0 8304 480 8424 6 chanx_left_in[13]
port 16 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[14]
port 17 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[15]
port 18 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[16]
port 19 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[17]
port 20 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[18]
port 21 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[19]
port 22 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[1]
port 23 nsew default input
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[2]
port 24 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[3]
port 25 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[4]
port 26 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[5]
port 27 nsew default input
rlabel metal3 s 0 5584 480 5704 6 chanx_left_in[6]
port 28 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[7]
port 29 nsew default input
rlabel metal3 s 0 6400 480 6520 6 chanx_left_in[8]
port 30 nsew default input
rlabel metal3 s 0 6808 480 6928 6 chanx_left_in[9]
port 31 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_out[0]
port 32 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 chanx_left_out[10]
port 33 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[11]
port 34 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 chanx_left_out[12]
port 35 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 chanx_left_out[13]
port 36 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[14]
port 37 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chanx_left_out[15]
port 38 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[16]
port 39 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[17]
port 40 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[18]
port 41 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chanx_left_out[19]
port 42 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[1]
port 43 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 chanx_left_out[2]
port 44 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 12656 480 12776 6 chanx_left_out[4]
port 46 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 chanx_left_out[5]
port 47 nsew default tristate
rlabel metal3 s 0 13472 480 13592 6 chanx_left_out[6]
port 48 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[7]
port 49 nsew default tristate
rlabel metal3 s 0 14288 480 14408 6 chanx_left_out[8]
port 50 nsew default tristate
rlabel metal3 s 0 14696 480 14816 6 chanx_left_out[9]
port 51 nsew default tristate
rlabel metal3 s 22320 3272 22800 3392 6 chanx_right_in[0]
port 52 nsew default input
rlabel metal3 s 22320 7216 22800 7336 6 chanx_right_in[10]
port 53 nsew default input
rlabel metal3 s 22320 7624 22800 7744 6 chanx_right_in[11]
port 54 nsew default input
rlabel metal3 s 22320 7896 22800 8016 6 chanx_right_in[12]
port 55 nsew default input
rlabel metal3 s 22320 8304 22800 8424 6 chanx_right_in[13]
port 56 nsew default input
rlabel metal3 s 22320 8712 22800 8832 6 chanx_right_in[14]
port 57 nsew default input
rlabel metal3 s 22320 9120 22800 9240 6 chanx_right_in[15]
port 58 nsew default input
rlabel metal3 s 22320 9528 22800 9648 6 chanx_right_in[16]
port 59 nsew default input
rlabel metal3 s 22320 9936 22800 10056 6 chanx_right_in[17]
port 60 nsew default input
rlabel metal3 s 22320 10344 22800 10464 6 chanx_right_in[18]
port 61 nsew default input
rlabel metal3 s 22320 10752 22800 10872 6 chanx_right_in[19]
port 62 nsew default input
rlabel metal3 s 22320 3680 22800 3800 6 chanx_right_in[1]
port 63 nsew default input
rlabel metal3 s 22320 3952 22800 4072 6 chanx_right_in[2]
port 64 nsew default input
rlabel metal3 s 22320 4360 22800 4480 6 chanx_right_in[3]
port 65 nsew default input
rlabel metal3 s 22320 4768 22800 4888 6 chanx_right_in[4]
port 66 nsew default input
rlabel metal3 s 22320 5176 22800 5296 6 chanx_right_in[5]
port 67 nsew default input
rlabel metal3 s 22320 5584 22800 5704 6 chanx_right_in[6]
port 68 nsew default input
rlabel metal3 s 22320 5992 22800 6112 6 chanx_right_in[7]
port 69 nsew default input
rlabel metal3 s 22320 6400 22800 6520 6 chanx_right_in[8]
port 70 nsew default input
rlabel metal3 s 22320 6808 22800 6928 6 chanx_right_in[9]
port 71 nsew default input
rlabel metal3 s 22320 11160 22800 11280 6 chanx_right_out[0]
port 72 nsew default tristate
rlabel metal3 s 22320 15104 22800 15224 6 chanx_right_out[10]
port 73 nsew default tristate
rlabel metal3 s 22320 15376 22800 15496 6 chanx_right_out[11]
port 74 nsew default tristate
rlabel metal3 s 22320 15784 22800 15904 6 chanx_right_out[12]
port 75 nsew default tristate
rlabel metal3 s 22320 16192 22800 16312 6 chanx_right_out[13]
port 76 nsew default tristate
rlabel metal3 s 22320 16600 22800 16720 6 chanx_right_out[14]
port 77 nsew default tristate
rlabel metal3 s 22320 17008 22800 17128 6 chanx_right_out[15]
port 78 nsew default tristate
rlabel metal3 s 22320 17416 22800 17536 6 chanx_right_out[16]
port 79 nsew default tristate
rlabel metal3 s 22320 17824 22800 17944 6 chanx_right_out[17]
port 80 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[18]
port 81 nsew default tristate
rlabel metal3 s 22320 18640 22800 18760 6 chanx_right_out[19]
port 82 nsew default tristate
rlabel metal3 s 22320 11568 22800 11688 6 chanx_right_out[1]
port 83 nsew default tristate
rlabel metal3 s 22320 11840 22800 11960 6 chanx_right_out[2]
port 84 nsew default tristate
rlabel metal3 s 22320 12248 22800 12368 6 chanx_right_out[3]
port 85 nsew default tristate
rlabel metal3 s 22320 12656 22800 12776 6 chanx_right_out[4]
port 86 nsew default tristate
rlabel metal3 s 22320 13064 22800 13184 6 chanx_right_out[5]
port 87 nsew default tristate
rlabel metal3 s 22320 13472 22800 13592 6 chanx_right_out[6]
port 88 nsew default tristate
rlabel metal3 s 22320 13880 22800 14000 6 chanx_right_out[7]
port 89 nsew default tristate
rlabel metal3 s 22320 14288 22800 14408 6 chanx_right_out[8]
port 90 nsew default tristate
rlabel metal3 s 22320 14696 22800 14816 6 chanx_right_out[9]
port 91 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 chany_bottom_in[0]
port 92 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[10]
port 93 nsew default input
rlabel metal2 s 8022 0 8078 480 6 chany_bottom_in[11]
port 94 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[12]
port 95 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chany_bottom_in[13]
port 96 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[14]
port 97 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[15]
port 98 nsew default input
rlabel metal2 s 9862 0 9918 480 6 chany_bottom_in[16]
port 99 nsew default input
rlabel metal2 s 10230 0 10286 480 6 chany_bottom_in[17]
port 100 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[18]
port 101 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[19]
port 102 nsew default input
rlabel metal2 s 4250 0 4306 480 6 chany_bottom_in[1]
port 103 nsew default input
rlabel metal2 s 4618 0 4674 480 6 chany_bottom_in[2]
port 104 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[3]
port 105 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_in[4]
port 106 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[5]
port 107 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[6]
port 108 nsew default input
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[7]
port 109 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[8]
port 110 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[9]
port 111 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_out[0]
port 112 nsew default tristate
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_out[10]
port 113 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[11]
port 114 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[12]
port 115 nsew default tristate
rlabel metal2 s 16210 0 16266 480 6 chany_bottom_out[13]
port 116 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[14]
port 117 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chany_bottom_out[15]
port 118 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[16]
port 119 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_out[17]
port 120 nsew default tristate
rlabel metal2 s 18142 0 18198 480 6 chany_bottom_out[18]
port 121 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 chany_bottom_out[19]
port 122 nsew default tristate
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_out[1]
port 123 nsew default tristate
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_out[2]
port 124 nsew default tristate
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_out[3]
port 125 nsew default tristate
rlabel metal2 s 12898 0 12954 480 6 chany_bottom_out[4]
port 126 nsew default tristate
rlabel metal2 s 13266 0 13322 480 6 chany_bottom_out[5]
port 127 nsew default tristate
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_out[6]
port 128 nsew default tristate
rlabel metal2 s 14002 0 14058 480 6 chany_bottom_out[7]
port 129 nsew default tristate
rlabel metal2 s 14370 0 14426 480 6 chany_bottom_out[8]
port 130 nsew default tristate
rlabel metal2 s 14738 0 14794 480 6 chany_bottom_out[9]
port 131 nsew default tristate
rlabel metal2 s 3238 22320 3294 22800 6 chany_top_in[0]
port 132 nsew default input
rlabel metal2 s 7010 22320 7066 22800 6 chany_top_in[10]
port 133 nsew default input
rlabel metal2 s 7378 22320 7434 22800 6 chany_top_in[11]
port 134 nsew default input
rlabel metal2 s 7746 22320 7802 22800 6 chany_top_in[12]
port 135 nsew default input
rlabel metal2 s 8114 22320 8170 22800 6 chany_top_in[13]
port 136 nsew default input
rlabel metal2 s 8482 22320 8538 22800 6 chany_top_in[14]
port 137 nsew default input
rlabel metal2 s 8942 22320 8998 22800 6 chany_top_in[15]
port 138 nsew default input
rlabel metal2 s 9310 22320 9366 22800 6 chany_top_in[16]
port 139 nsew default input
rlabel metal2 s 9678 22320 9734 22800 6 chany_top_in[17]
port 140 nsew default input
rlabel metal2 s 10046 22320 10102 22800 6 chany_top_in[18]
port 141 nsew default input
rlabel metal2 s 10414 22320 10470 22800 6 chany_top_in[19]
port 142 nsew default input
rlabel metal2 s 3606 22320 3662 22800 6 chany_top_in[1]
port 143 nsew default input
rlabel metal2 s 3974 22320 4030 22800 6 chany_top_in[2]
port 144 nsew default input
rlabel metal2 s 4342 22320 4398 22800 6 chany_top_in[3]
port 145 nsew default input
rlabel metal2 s 4710 22320 4766 22800 6 chany_top_in[4]
port 146 nsew default input
rlabel metal2 s 5078 22320 5134 22800 6 chany_top_in[5]
port 147 nsew default input
rlabel metal2 s 5446 22320 5502 22800 6 chany_top_in[6]
port 148 nsew default input
rlabel metal2 s 5906 22320 5962 22800 6 chany_top_in[7]
port 149 nsew default input
rlabel metal2 s 6274 22320 6330 22800 6 chany_top_in[8]
port 150 nsew default input
rlabel metal2 s 6642 22320 6698 22800 6 chany_top_in[9]
port 151 nsew default input
rlabel metal2 s 10782 22320 10838 22800 6 chany_top_out[0]
port 152 nsew default tristate
rlabel metal2 s 14646 22320 14702 22800 6 chany_top_out[10]
port 153 nsew default tristate
rlabel metal2 s 15014 22320 15070 22800 6 chany_top_out[11]
port 154 nsew default tristate
rlabel metal2 s 15382 22320 15438 22800 6 chany_top_out[12]
port 155 nsew default tristate
rlabel metal2 s 15750 22320 15806 22800 6 chany_top_out[13]
port 156 nsew default tristate
rlabel metal2 s 16118 22320 16174 22800 6 chany_top_out[14]
port 157 nsew default tristate
rlabel metal2 s 16486 22320 16542 22800 6 chany_top_out[15]
port 158 nsew default tristate
rlabel metal2 s 16854 22320 16910 22800 6 chany_top_out[16]
port 159 nsew default tristate
rlabel metal2 s 17314 22320 17370 22800 6 chany_top_out[17]
port 160 nsew default tristate
rlabel metal2 s 17682 22320 17738 22800 6 chany_top_out[18]
port 161 nsew default tristate
rlabel metal2 s 18050 22320 18106 22800 6 chany_top_out[19]
port 162 nsew default tristate
rlabel metal2 s 11150 22320 11206 22800 6 chany_top_out[1]
port 163 nsew default tristate
rlabel metal2 s 11610 22320 11666 22800 6 chany_top_out[2]
port 164 nsew default tristate
rlabel metal2 s 11978 22320 12034 22800 6 chany_top_out[3]
port 165 nsew default tristate
rlabel metal2 s 12346 22320 12402 22800 6 chany_top_out[4]
port 166 nsew default tristate
rlabel metal2 s 12714 22320 12770 22800 6 chany_top_out[5]
port 167 nsew default tristate
rlabel metal2 s 13082 22320 13138 22800 6 chany_top_out[6]
port 168 nsew default tristate
rlabel metal2 s 13450 22320 13506 22800 6 chany_top_out[7]
port 169 nsew default tristate
rlabel metal2 s 13818 22320 13874 22800 6 chany_top_out[8]
port 170 nsew default tristate
rlabel metal2 s 14186 22320 14242 22800 6 chany_top_out[9]
port 171 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 clk_1_E_out
port 172 nsew default tristate
rlabel metal2 s 18786 22320 18842 22800 6 clk_1_N_in
port 173 nsew default input
rlabel metal2 s 19246 0 19302 480 6 clk_1_S_in
port 174 nsew default input
rlabel metal3 s 0 19048 480 19168 6 clk_1_W_out
port 175 nsew default tristate
rlabel metal3 s 22320 19048 22800 19168 6 clk_2_E_in
port 176 nsew default input
rlabel metal3 s 22320 20952 22800 21072 6 clk_2_E_out
port 177 nsew default tristate
rlabel metal2 s 19154 22320 19210 22800 6 clk_2_N_in
port 178 nsew default input
rlabel metal2 s 21454 22320 21510 22800 6 clk_2_N_out
port 179 nsew default tristate
rlabel metal2 s 19614 0 19670 480 6 clk_2_S_in
port 180 nsew default input
rlabel metal2 s 20350 0 20406 480 6 clk_2_S_out
port 181 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 clk_2_W_in
port 182 nsew default input
rlabel metal3 s 0 19320 480 19440 6 clk_2_W_out
port 183 nsew default tristate
rlabel metal3 s 22320 19320 22800 19440 6 clk_3_E_in
port 184 nsew default input
rlabel metal3 s 22320 21360 22800 21480 6 clk_3_E_out
port 185 nsew default tristate
rlabel metal2 s 19522 22320 19578 22800 6 clk_3_N_in
port 186 nsew default input
rlabel metal2 s 21822 22320 21878 22800 6 clk_3_N_out
port 187 nsew default tristate
rlabel metal2 s 19982 0 20038 480 6 clk_3_S_in
port 188 nsew default input
rlabel metal2 s 20718 0 20774 480 6 clk_3_S_out
port 189 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 clk_3_W_in
port 190 nsew default input
rlabel metal3 s 0 19728 480 19848 6 clk_3_W_out
port 191 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 192 nsew default input
rlabel metal3 s 0 416 480 536 6 left_bottom_grid_pin_35_
port 193 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_36_
port 194 nsew default input
rlabel metal3 s 0 1232 480 1352 6 left_bottom_grid_pin_37_
port 195 nsew default input
rlabel metal3 s 0 1640 480 1760 6 left_bottom_grid_pin_38_
port 196 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_39_
port 197 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_40_
port 198 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_41_
port 199 nsew default input
rlabel metal2 s 19890 22320 19946 22800 6 prog_clk_0_N_in
port 200 nsew default input
rlabel metal3 s 22320 21768 22800 21888 6 prog_clk_1_E_out
port 201 nsew default tristate
rlabel metal2 s 20350 22320 20406 22800 6 prog_clk_1_N_in
port 202 nsew default input
rlabel metal2 s 21086 0 21142 480 6 prog_clk_1_S_in
port 203 nsew default input
rlabel metal3 s 0 20136 480 20256 6 prog_clk_1_W_out
port 204 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 prog_clk_2_E_in
port 205 nsew default input
rlabel metal3 s 22320 22176 22800 22296 6 prog_clk_2_E_out
port 206 nsew default tristate
rlabel metal2 s 20718 22320 20774 22800 6 prog_clk_2_N_in
port 207 nsew default input
rlabel metal2 s 22190 22320 22246 22800 6 prog_clk_2_N_out
port 208 nsew default tristate
rlabel metal2 s 21454 0 21510 480 6 prog_clk_2_S_in
port 209 nsew default input
rlabel metal2 s 22190 0 22246 480 6 prog_clk_2_S_out
port 210 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 prog_clk_2_W_in
port 211 nsew default input
rlabel metal3 s 0 20544 480 20664 6 prog_clk_2_W_out
port 212 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 prog_clk_3_E_in
port 213 nsew default input
rlabel metal3 s 22320 22584 22800 22704 6 prog_clk_3_E_out
port 214 nsew default tristate
rlabel metal2 s 21086 22320 21142 22800 6 prog_clk_3_N_in
port 215 nsew default input
rlabel metal2 s 22558 22320 22614 22800 6 prog_clk_3_N_out
port 216 nsew default tristate
rlabel metal2 s 21822 0 21878 480 6 prog_clk_3_S_in
port 217 nsew default input
rlabel metal2 s 22558 0 22614 480 6 prog_clk_3_S_out
port 218 nsew default tristate
rlabel metal3 s 0 22584 480 22704 6 prog_clk_3_W_in
port 219 nsew default input
rlabel metal3 s 0 20952 480 21072 6 prog_clk_3_W_out
port 220 nsew default tristate
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_34_
port 221 nsew default input
rlabel metal3 s 22320 416 22800 536 6 right_bottom_grid_pin_35_
port 222 nsew default input
rlabel metal3 s 22320 824 22800 944 6 right_bottom_grid_pin_36_
port 223 nsew default input
rlabel metal3 s 22320 1232 22800 1352 6 right_bottom_grid_pin_37_
port 224 nsew default input
rlabel metal3 s 22320 1640 22800 1760 6 right_bottom_grid_pin_38_
port 225 nsew default input
rlabel metal3 s 22320 2048 22800 2168 6 right_bottom_grid_pin_39_
port 226 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_40_
port 227 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_41_
port 228 nsew default input
rlabel metal2 s 202 22320 258 22800 6 top_left_grid_pin_42_
port 229 nsew default input
rlabel metal2 s 570 22320 626 22800 6 top_left_grid_pin_43_
port 230 nsew default input
rlabel metal2 s 938 22320 994 22800 6 top_left_grid_pin_44_
port 231 nsew default input
rlabel metal2 s 1306 22320 1362 22800 6 top_left_grid_pin_45_
port 232 nsew default input
rlabel metal2 s 1674 22320 1730 22800 6 top_left_grid_pin_46_
port 233 nsew default input
rlabel metal2 s 2042 22320 2098 22800 6 top_left_grid_pin_47_
port 234 nsew default input
rlabel metal2 s 2410 22320 2466 22800 6 top_left_grid_pin_48_
port 235 nsew default input
rlabel metal2 s 2778 22320 2834 22800 6 top_left_grid_pin_49_
port 236 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 237 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 238 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
