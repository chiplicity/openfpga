magic
tech sky130A
magscale 1 2
timestamp 1606224842
<< locali >>
rect 3433 14467 3467 14569
rect 9505 11067 9539 11169
rect 9781 3995 9815 4165
rect 12265 2975 12299 3077
rect 6101 1479 6135 1853
<< viali >>
rect 1593 15657 1627 15691
rect 5733 15657 5767 15691
rect 9965 15657 9999 15691
rect 10977 15657 11011 15691
rect 13737 15657 13771 15691
rect 14473 15657 14507 15691
rect 4813 15589 4847 15623
rect 7297 15589 7331 15623
rect 8493 15589 8527 15623
rect 12909 15589 12943 15623
rect 1409 15521 1443 15555
rect 2412 15521 2446 15555
rect 4721 15521 4755 15555
rect 5549 15521 5583 15555
rect 7389 15521 7423 15555
rect 8585 15521 8619 15555
rect 9781 15521 9815 15555
rect 11345 15521 11379 15555
rect 12633 15521 12667 15555
rect 13553 15521 13587 15555
rect 14289 15521 14323 15555
rect 2145 15453 2179 15487
rect 4997 15453 5031 15487
rect 7481 15453 7515 15487
rect 8677 15453 8711 15487
rect 11437 15453 11471 15487
rect 11621 15453 11655 15487
rect 4353 15385 4387 15419
rect 3525 15317 3559 15351
rect 6929 15317 6963 15351
rect 8125 15317 8159 15351
rect 1685 15113 1719 15147
rect 4813 15113 4847 15147
rect 6193 15113 6227 15147
rect 8033 15113 8067 15147
rect 8585 15113 8619 15147
rect 9965 15113 9999 15147
rect 2973 15045 3007 15079
rect 13829 15045 13863 15079
rect 4077 14977 4111 15011
rect 4261 14977 4295 15011
rect 5457 14977 5491 15011
rect 9229 14977 9263 15011
rect 11713 14977 11747 15011
rect 13093 14977 13127 15011
rect 1501 14909 1535 14943
rect 2789 14909 2823 14943
rect 6009 14909 6043 14943
rect 6837 14909 6871 14943
rect 7849 14909 7883 14943
rect 9781 14909 9815 14943
rect 11437 14909 11471 14943
rect 13645 14909 13679 14943
rect 14381 14909 14415 14943
rect 5273 14841 5307 14875
rect 9045 14841 9079 14875
rect 3617 14773 3651 14807
rect 3985 14773 4019 14807
rect 5181 14773 5215 14807
rect 7021 14773 7055 14807
rect 8953 14773 8987 14807
rect 11069 14773 11103 14807
rect 11529 14773 11563 14807
rect 12449 14773 12483 14807
rect 12817 14773 12851 14807
rect 12909 14773 12943 14807
rect 14565 14773 14599 14807
rect 1961 14569 1995 14603
rect 3433 14569 3467 14603
rect 3525 14569 3559 14603
rect 6561 14569 6595 14603
rect 7757 14569 7791 14603
rect 12449 14569 12483 14603
rect 12541 14569 12575 14603
rect 2789 14501 2823 14535
rect 8861 14501 8895 14535
rect 13553 14501 13587 14535
rect 1777 14433 1811 14467
rect 2513 14433 2547 14467
rect 3433 14433 3467 14467
rect 3709 14433 3743 14467
rect 4609 14433 4643 14467
rect 7849 14433 7883 14467
rect 8585 14433 8619 14467
rect 9956 14433 9990 14467
rect 13277 14433 13311 14467
rect 14197 14433 14231 14467
rect 4353 14365 4387 14399
rect 6653 14365 6687 14399
rect 6745 14365 6779 14399
rect 8033 14365 8067 14399
rect 9689 14365 9723 14399
rect 12725 14365 12759 14399
rect 5733 14297 5767 14331
rect 6193 14297 6227 14331
rect 12081 14297 12115 14331
rect 7389 14229 7423 14263
rect 11069 14229 11103 14263
rect 14381 14229 14415 14263
rect 2513 14025 2547 14059
rect 3249 14025 3283 14059
rect 7297 14025 7331 14059
rect 10333 14025 10367 14059
rect 1777 13957 1811 13991
rect 4169 13957 4203 13991
rect 5365 13957 5399 13991
rect 9873 13957 9907 13991
rect 15025 13957 15059 13991
rect 4813 13889 4847 13923
rect 5825 13889 5859 13923
rect 5917 13889 5951 13923
rect 7941 13889 7975 13923
rect 10885 13889 10919 13923
rect 12909 13889 12943 13923
rect 13001 13889 13035 13923
rect 14197 13889 14231 13923
rect 1593 13821 1627 13855
rect 2329 13821 2363 13855
rect 3433 13821 3467 13855
rect 7665 13821 7699 13855
rect 8493 13821 8527 13855
rect 14105 13821 14139 13855
rect 14841 13821 14875 13855
rect 4537 13753 4571 13787
rect 4629 13753 4663 13787
rect 5733 13753 5767 13787
rect 8760 13753 8794 13787
rect 12817 13753 12851 13787
rect 14013 13753 14047 13787
rect 3525 13685 3559 13719
rect 7757 13685 7791 13719
rect 10701 13685 10735 13719
rect 10793 13685 10827 13719
rect 11529 13685 11563 13719
rect 12449 13685 12483 13719
rect 13645 13685 13679 13719
rect 8401 13481 8435 13515
rect 12725 13481 12759 13515
rect 14289 13481 14323 13515
rect 5264 13413 5298 13447
rect 8769 13413 8803 13447
rect 8861 13413 8895 13447
rect 14381 13413 14415 13447
rect 1409 13345 1443 13379
rect 2145 13345 2179 13379
rect 2412 13345 2446 13379
rect 7205 13345 7239 13379
rect 7297 13345 7331 13379
rect 8217 13345 8251 13379
rect 10681 13345 10715 13379
rect 12449 13345 12483 13379
rect 13093 13345 13127 13379
rect 13185 13345 13219 13379
rect 4353 13277 4387 13311
rect 4997 13277 5031 13311
rect 7481 13277 7515 13311
rect 8953 13277 8987 13311
rect 9781 13277 9815 13311
rect 10425 13277 10459 13311
rect 13277 13277 13311 13311
rect 14473 13277 14507 13311
rect 11805 13209 11839 13243
rect 1593 13141 1627 13175
rect 3525 13141 3559 13175
rect 6377 13141 6411 13175
rect 6837 13141 6871 13175
rect 8033 13141 8067 13175
rect 12265 13141 12299 13175
rect 13921 13141 13955 13175
rect 3157 12937 3191 12971
rect 8953 12937 8987 12971
rect 13645 12937 13679 12971
rect 5549 12869 5583 12903
rect 10793 12869 10827 12903
rect 12449 12869 12483 12903
rect 15025 12869 15059 12903
rect 2605 12801 2639 12835
rect 3801 12801 3835 12835
rect 4997 12801 5031 12835
rect 6009 12801 6043 12835
rect 6101 12801 6135 12835
rect 8355 12801 8389 12835
rect 9597 12801 9631 12835
rect 11345 12801 11379 12835
rect 13001 12801 13035 12835
rect 14197 12801 14231 12835
rect 2329 12733 2363 12767
rect 3525 12733 3559 12767
rect 6837 12733 6871 12767
rect 8125 12733 8159 12767
rect 11161 12733 11195 12767
rect 12909 12733 12943 12767
rect 14841 12733 14875 12767
rect 3617 12665 3651 12699
rect 4813 12665 4847 12699
rect 7113 12665 7147 12699
rect 9321 12665 9355 12699
rect 14105 12665 14139 12699
rect 1961 12597 1995 12631
rect 2421 12597 2455 12631
rect 4353 12597 4387 12631
rect 4721 12597 4755 12631
rect 5917 12597 5951 12631
rect 7757 12597 7791 12631
rect 8217 12597 8251 12631
rect 9413 12597 9447 12631
rect 10149 12597 10183 12631
rect 11253 12597 11287 12631
rect 12817 12597 12851 12631
rect 14013 12597 14047 12631
rect 1961 12393 1995 12427
rect 3157 12393 3191 12427
rect 3249 12393 3283 12427
rect 7941 12393 7975 12427
rect 11069 12393 11103 12427
rect 12081 12393 12115 12427
rect 12449 12393 12483 12427
rect 4077 12325 4111 12359
rect 6828 12325 6862 12359
rect 8769 12325 8803 12359
rect 2053 12257 2087 12291
rect 4721 12257 4755 12291
rect 4988 12257 5022 12291
rect 9945 12257 9979 12291
rect 11713 12257 11747 12291
rect 13277 12257 13311 12291
rect 14197 12257 14231 12291
rect 2237 12189 2271 12223
rect 3433 12189 3467 12223
rect 6568 12189 6602 12223
rect 8861 12189 8895 12223
rect 9045 12189 9079 12223
rect 9689 12189 9723 12223
rect 12541 12189 12575 12223
rect 12633 12189 12667 12223
rect 13461 12189 13495 12223
rect 14381 12189 14415 12223
rect 1593 12121 1627 12155
rect 8401 12121 8435 12155
rect 11529 12121 11563 12155
rect 2789 12053 2823 12087
rect 6101 12053 6135 12087
rect 1869 11849 1903 11883
rect 11897 11849 11931 11883
rect 6285 11781 6319 11815
rect 8217 11781 8251 11815
rect 2513 11713 2547 11747
rect 3065 11713 3099 11747
rect 9965 11713 9999 11747
rect 10609 11713 10643 11747
rect 11253 11713 11287 11747
rect 13001 11713 13035 11747
rect 2237 11645 2271 11679
rect 4905 11645 4939 11679
rect 6837 11645 6871 11679
rect 7093 11645 7127 11679
rect 8677 11645 8711 11679
rect 9873 11645 9907 11679
rect 12081 11645 12115 11679
rect 13645 11645 13679 11679
rect 14381 11645 14415 11679
rect 2329 11577 2363 11611
rect 3332 11577 3366 11611
rect 5150 11577 5184 11611
rect 12817 11577 12851 11611
rect 4445 11509 4479 11543
rect 8861 11509 8895 11543
rect 9413 11509 9447 11543
rect 9781 11509 9815 11543
rect 12449 11509 12483 11543
rect 12909 11509 12943 11543
rect 13829 11509 13863 11543
rect 14565 11509 14599 11543
rect 1593 11305 1627 11339
rect 1961 11305 1995 11339
rect 2789 11305 2823 11339
rect 4353 11305 4387 11339
rect 4813 11305 4847 11339
rect 6929 11305 6963 11339
rect 9229 11305 9263 11339
rect 9689 11305 9723 11339
rect 11345 11305 11379 11339
rect 12081 11305 12115 11339
rect 13737 11305 13771 11339
rect 2053 11237 2087 11271
rect 3157 11237 3191 11271
rect 7634 11237 7668 11271
rect 10057 11237 10091 11271
rect 12449 11237 12483 11271
rect 12541 11237 12575 11271
rect 4721 11169 4755 11203
rect 5816 11169 5850 11203
rect 7389 11169 7423 11203
rect 9413 11169 9447 11203
rect 9505 11169 9539 11203
rect 10149 11169 10183 11203
rect 11253 11169 11287 11203
rect 13645 11169 13679 11203
rect 14473 11169 14507 11203
rect 2237 11101 2271 11135
rect 3249 11101 3283 11135
rect 3341 11101 3375 11135
rect 4997 11101 5031 11135
rect 5549 11101 5583 11135
rect 10241 11101 10275 11135
rect 11529 11101 11563 11135
rect 12633 11101 12667 11135
rect 13829 11101 13863 11135
rect 8769 11033 8803 11067
rect 9505 11033 9539 11067
rect 10885 11033 10919 11067
rect 13277 11033 13311 11067
rect 14657 10965 14691 10999
rect 6285 10761 6319 10795
rect 8677 10761 8711 10795
rect 9873 10761 9907 10795
rect 12449 10761 12483 10795
rect 2053 10625 2087 10659
rect 2697 10625 2731 10659
rect 2881 10625 2915 10659
rect 3065 10625 3099 10659
rect 4905 10625 4939 10659
rect 9137 10625 9171 10659
rect 9229 10625 9263 10659
rect 10517 10625 10551 10659
rect 11621 10625 11655 10659
rect 13001 10625 13035 10659
rect 14749 10625 14783 10659
rect 1777 10557 1811 10591
rect 6837 10557 6871 10591
rect 7104 10557 7138 10591
rect 10241 10557 10275 10591
rect 10333 10557 10367 10591
rect 11437 10557 11471 10591
rect 13645 10557 13679 10591
rect 14565 10557 14599 10591
rect 2605 10489 2639 10523
rect 3332 10489 3366 10523
rect 5172 10489 5206 10523
rect 9045 10489 9079 10523
rect 12817 10489 12851 10523
rect 13921 10489 13955 10523
rect 1409 10421 1443 10455
rect 1869 10421 1903 10455
rect 2237 10421 2271 10455
rect 4445 10421 4479 10455
rect 8217 10421 8251 10455
rect 11069 10421 11103 10455
rect 11529 10421 11563 10455
rect 12909 10421 12943 10455
rect 1501 10217 1535 10251
rect 2789 10217 2823 10251
rect 7113 10217 7147 10251
rect 8953 10217 8987 10251
rect 11345 10217 11379 10251
rect 12081 10217 12115 10251
rect 12449 10217 12483 10251
rect 13277 10217 13311 10251
rect 1869 10149 1903 10183
rect 4905 10149 4939 10183
rect 5978 10149 6012 10183
rect 7818 10149 7852 10183
rect 10149 10149 10183 10183
rect 13645 10149 13679 10183
rect 2697 10081 2731 10115
rect 3525 10081 3559 10115
rect 10057 10081 10091 10115
rect 11253 10081 11287 10115
rect 14473 10081 14507 10115
rect 1961 10013 1995 10047
rect 2145 10013 2179 10047
rect 2973 10013 3007 10047
rect 3617 10013 3651 10047
rect 3801 10013 3835 10047
rect 4997 10013 5031 10047
rect 5181 10013 5215 10047
rect 5733 10013 5767 10047
rect 7573 10013 7607 10047
rect 10333 10013 10367 10047
rect 11529 10013 11563 10047
rect 12541 10013 12575 10047
rect 12633 10013 12667 10047
rect 13737 10013 13771 10047
rect 13829 10013 13863 10047
rect 4537 9945 4571 9979
rect 10885 9945 10919 9979
rect 14657 9945 14691 9979
rect 2329 9877 2363 9911
rect 3157 9877 3191 9911
rect 9689 9877 9723 9911
rect 8217 9673 8251 9707
rect 2789 9605 2823 9639
rect 6653 9605 6687 9639
rect 9873 9605 9907 9639
rect 15025 9605 15059 9639
rect 2237 9537 2271 9571
rect 3433 9537 3467 9571
rect 3801 9537 3835 9571
rect 5273 9537 5307 9571
rect 9229 9537 9263 9571
rect 10425 9537 10459 9571
rect 11621 9537 11655 9571
rect 12909 9537 12943 9571
rect 13093 9537 13127 9571
rect 14197 9537 14231 9571
rect 2053 9469 2087 9503
rect 4057 9469 4091 9503
rect 6837 9469 6871 9503
rect 9045 9469 9079 9503
rect 9137 9469 9171 9503
rect 14013 9469 14047 9503
rect 14841 9469 14875 9503
rect 1961 9401 1995 9435
rect 3249 9401 3283 9435
rect 5540 9401 5574 9435
rect 7104 9401 7138 9435
rect 10241 9401 10275 9435
rect 1593 9333 1627 9367
rect 3157 9333 3191 9367
rect 5181 9333 5215 9367
rect 8677 9333 8711 9367
rect 10333 9333 10367 9367
rect 11069 9333 11103 9367
rect 11437 9333 11471 9367
rect 11529 9333 11563 9367
rect 12449 9333 12483 9367
rect 12817 9333 12851 9367
rect 13645 9333 13679 9367
rect 14105 9333 14139 9367
rect 2329 9129 2363 9163
rect 4353 9129 4387 9163
rect 4721 9129 4755 9163
rect 10149 9129 10183 9163
rect 11253 9129 11287 9163
rect 12081 9129 12115 9163
rect 1685 9061 1719 9095
rect 3157 9061 3191 9095
rect 3249 9061 3283 9095
rect 7481 9061 7515 9095
rect 10057 9061 10091 9095
rect 12449 9061 12483 9095
rect 12541 9061 12575 9095
rect 1409 8993 1443 9027
rect 5825 8993 5859 9027
rect 7665 8993 7699 9027
rect 7932 8993 7966 9027
rect 11345 8993 11379 9027
rect 13277 8993 13311 9027
rect 14197 8993 14231 9027
rect 2421 8925 2455 8959
rect 2605 8925 2639 8959
rect 3433 8925 3467 8959
rect 4813 8925 4847 8959
rect 4997 8925 5031 8959
rect 10333 8925 10367 8959
rect 11437 8925 11471 8959
rect 12725 8925 12759 8959
rect 13461 8925 13495 8959
rect 14473 8925 14507 8959
rect 9689 8857 9723 8891
rect 10885 8857 10919 8891
rect 1961 8789 1995 8823
rect 2789 8789 2823 8823
rect 9045 8789 9079 8823
rect 1869 8585 1903 8619
rect 2697 8585 2731 8619
rect 4077 8585 4111 8619
rect 6285 8585 6319 8619
rect 10057 8585 10091 8619
rect 12449 8585 12483 8619
rect 8217 8517 8251 8551
rect 10517 8517 10551 8551
rect 13645 8517 13679 8551
rect 2513 8449 2547 8483
rect 3249 8449 3283 8483
rect 3709 8449 3743 8483
rect 4537 8449 4571 8483
rect 4721 8449 4755 8483
rect 6837 8449 6871 8483
rect 11069 8449 11103 8483
rect 11713 8449 11747 8483
rect 12909 8449 12943 8483
rect 13093 8449 13127 8483
rect 14197 8449 14231 8483
rect 2237 8381 2271 8415
rect 3525 8381 3559 8415
rect 4905 8381 4939 8415
rect 7093 8381 7127 8415
rect 8677 8381 8711 8415
rect 10977 8381 11011 8415
rect 14105 8381 14139 8415
rect 14841 8381 14875 8415
rect 3157 8313 3191 8347
rect 4445 8313 4479 8347
rect 5172 8313 5206 8347
rect 8922 8313 8956 8347
rect 10885 8313 10919 8347
rect 14013 8313 14047 8347
rect 2329 8245 2363 8279
rect 3065 8245 3099 8279
rect 12817 8245 12851 8279
rect 15025 8245 15059 8279
rect 2421 8041 2455 8075
rect 2881 8041 2915 8075
rect 4077 8041 4111 8075
rect 8861 8041 8895 8075
rect 11529 8041 11563 8075
rect 11897 8041 11931 8075
rect 13093 8041 13127 8075
rect 14289 8041 14323 8075
rect 7726 7973 7760 8007
rect 11989 7973 12023 8007
rect 1961 7905 1995 7939
rect 2053 7905 2087 7939
rect 2789 7905 2823 7939
rect 3801 7905 3835 7939
rect 4445 7905 4479 7939
rect 5457 7905 5491 7939
rect 5641 7905 5675 7939
rect 5908 7905 5942 7939
rect 7481 7905 7515 7939
rect 9505 7905 9539 7939
rect 9945 7905 9979 7939
rect 2237 7837 2271 7871
rect 3065 7837 3099 7871
rect 4537 7837 4571 7871
rect 4721 7837 4755 7871
rect 9689 7837 9723 7871
rect 12081 7837 12115 7871
rect 13185 7837 13219 7871
rect 13277 7837 13311 7871
rect 14381 7837 14415 7871
rect 14565 7837 14599 7871
rect 9321 7769 9355 7803
rect 1593 7701 1627 7735
rect 3617 7701 3651 7735
rect 5273 7701 5307 7735
rect 7021 7701 7055 7735
rect 11069 7701 11103 7735
rect 12725 7701 12759 7735
rect 13921 7701 13955 7735
rect 6285 7497 6319 7531
rect 10517 7497 10551 7531
rect 12449 7497 12483 7531
rect 13645 7497 13679 7531
rect 2237 7429 2271 7463
rect 4445 7429 4479 7463
rect 8217 7429 8251 7463
rect 15025 7429 15059 7463
rect 1869 7361 1903 7395
rect 2053 7361 2087 7395
rect 2881 7361 2915 7395
rect 4905 7361 4939 7395
rect 6837 7361 6871 7395
rect 11069 7361 11103 7395
rect 13001 7361 13035 7395
rect 14105 7361 14139 7395
rect 14289 7361 14323 7395
rect 3065 7293 3099 7327
rect 8677 7293 8711 7327
rect 10885 7293 10919 7327
rect 12817 7293 12851 7327
rect 14841 7293 14875 7327
rect 2605 7225 2639 7259
rect 3332 7225 3366 7259
rect 5172 7225 5206 7259
rect 7104 7225 7138 7259
rect 8922 7225 8956 7259
rect 11713 7225 11747 7259
rect 1409 7157 1443 7191
rect 1777 7157 1811 7191
rect 2697 7157 2731 7191
rect 10057 7157 10091 7191
rect 10977 7157 11011 7191
rect 12909 7157 12943 7191
rect 14013 7157 14047 7191
rect 4445 6953 4479 6987
rect 11069 6953 11103 6987
rect 8953 6885 8987 6919
rect 9045 6885 9079 6919
rect 11897 6885 11931 6919
rect 13093 6885 13127 6919
rect 1409 6817 1443 6851
rect 2412 6817 2446 6851
rect 5540 6817 5574 6851
rect 7113 6817 7147 6851
rect 7369 6817 7403 6851
rect 9945 6817 9979 6851
rect 14289 6817 14323 6851
rect 2145 6749 2179 6783
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 5273 6749 5307 6783
rect 9137 6749 9171 6783
rect 9689 6749 9723 6783
rect 11989 6749 12023 6783
rect 12081 6749 12115 6783
rect 13185 6749 13219 6783
rect 13277 6749 13311 6783
rect 14381 6749 14415 6783
rect 14473 6749 14507 6783
rect 3525 6681 3559 6715
rect 8585 6681 8619 6715
rect 12725 6681 12759 6715
rect 13921 6681 13955 6715
rect 1593 6613 1627 6647
rect 4077 6613 4111 6647
rect 6653 6613 6687 6647
rect 8493 6613 8527 6647
rect 11529 6613 11563 6647
rect 2789 6409 2823 6443
rect 6929 6409 6963 6443
rect 10517 6409 10551 6443
rect 12449 6409 12483 6443
rect 13645 6409 13679 6443
rect 6285 6341 6319 6375
rect 15025 6341 15059 6375
rect 2145 6273 2179 6307
rect 3065 6273 3099 6307
rect 4905 6273 4939 6307
rect 7481 6273 7515 6307
rect 8033 6273 8067 6307
rect 9505 6273 9539 6307
rect 9873 6273 9907 6307
rect 11069 6273 11103 6307
rect 13001 6273 13035 6307
rect 14197 6273 14231 6307
rect 1961 6205 1995 6239
rect 2973 6205 3007 6239
rect 5172 6205 5206 6239
rect 7389 6205 7423 6239
rect 14013 6205 14047 6239
rect 14841 6205 14875 6239
rect 3332 6137 3366 6171
rect 8300 6137 8334 6171
rect 10885 6137 10919 6171
rect 14105 6137 14139 6171
rect 1593 6069 1627 6103
rect 2053 6069 2087 6103
rect 4445 6069 4479 6103
rect 7297 6069 7331 6103
rect 9413 6069 9447 6103
rect 10977 6069 11011 6103
rect 11713 6069 11747 6103
rect 12817 6069 12851 6103
rect 12909 6069 12943 6103
rect 1961 5865 1995 5899
rect 3525 5865 3559 5899
rect 7665 5865 7699 5899
rect 8769 5865 8803 5899
rect 8861 5865 8895 5899
rect 12725 5865 12759 5899
rect 13921 5865 13955 5899
rect 14381 5865 14415 5899
rect 4712 5797 4746 5831
rect 11897 5797 11931 5831
rect 1409 5729 1443 5763
rect 1777 5729 1811 5763
rect 2145 5729 2179 5763
rect 2412 5729 2446 5763
rect 6541 5729 6575 5763
rect 8285 5729 8319 5763
rect 9956 5729 9990 5763
rect 11989 5729 12023 5763
rect 13093 5729 13127 5763
rect 14289 5729 14323 5763
rect 4445 5661 4479 5695
rect 6285 5661 6319 5695
rect 8953 5661 8987 5695
rect 9689 5661 9723 5695
rect 12081 5661 12115 5695
rect 13185 5661 13219 5695
rect 13369 5661 13403 5695
rect 14565 5661 14599 5695
rect 1593 5593 1627 5627
rect 8125 5593 8159 5627
rect 8401 5593 8435 5627
rect 11529 5593 11563 5627
rect 5825 5525 5859 5559
rect 11069 5525 11103 5559
rect 6837 5321 6871 5355
rect 9229 5321 9263 5355
rect 10517 5321 10551 5355
rect 12449 5321 12483 5355
rect 9321 5253 9355 5287
rect 2237 5185 2271 5219
rect 2697 5185 2731 5219
rect 3065 5185 3099 5219
rect 6469 5185 6503 5219
rect 7389 5185 7423 5219
rect 9965 5185 9999 5219
rect 10977 5185 11011 5219
rect 11069 5185 11103 5219
rect 13093 5185 13127 5219
rect 14105 5185 14139 5219
rect 14197 5185 14231 5219
rect 2421 5117 2455 5151
rect 3332 5117 3366 5151
rect 4905 5117 4939 5151
rect 7849 5117 7883 5151
rect 9781 5117 9815 5151
rect 10149 5117 10183 5151
rect 14013 5117 14047 5151
rect 14841 5117 14875 5151
rect 1961 5049 1995 5083
rect 5150 5049 5184 5083
rect 8094 5049 8128 5083
rect 10885 5049 10919 5083
rect 12817 5049 12851 5083
rect 1593 4981 1627 5015
rect 2053 4981 2087 5015
rect 4445 4981 4479 5015
rect 6285 4981 6319 5015
rect 7205 4981 7239 5015
rect 7297 4981 7331 5015
rect 9689 4981 9723 5015
rect 11713 4981 11747 5015
rect 12909 4981 12943 5015
rect 13645 4981 13679 5015
rect 15025 4981 15059 5015
rect 3341 4777 3375 4811
rect 5457 4777 5491 4811
rect 10885 4777 10919 4811
rect 11253 4777 11287 4811
rect 12449 4777 12483 4811
rect 13737 4777 13771 4811
rect 3249 4709 3283 4743
rect 10149 4709 10183 4743
rect 13645 4709 13679 4743
rect 1676 4641 1710 4675
rect 4344 4641 4378 4675
rect 5917 4641 5951 4675
rect 6184 4641 6218 4675
rect 7389 4641 7423 4675
rect 8024 4641 8058 4675
rect 10057 4641 10091 4675
rect 11345 4641 11379 4675
rect 14473 4641 14507 4675
rect 3525 4573 3559 4607
rect 4077 4573 4111 4607
rect 7757 4573 7791 4607
rect 10241 4573 10275 4607
rect 11437 4573 11471 4607
rect 12541 4573 12575 4607
rect 12633 4573 12667 4607
rect 13829 4573 13863 4607
rect 2789 4505 2823 4539
rect 7573 4505 7607 4539
rect 9137 4505 9171 4539
rect 2881 4437 2915 4471
rect 7297 4437 7331 4471
rect 9689 4437 9723 4471
rect 12081 4437 12115 4471
rect 13277 4437 13311 4471
rect 14657 4437 14691 4471
rect 2789 4233 2823 4267
rect 6285 4233 6319 4267
rect 8309 4233 8343 4267
rect 9873 4233 9907 4267
rect 9781 4165 9815 4199
rect 12449 4165 12483 4199
rect 4905 4097 4939 4131
rect 6837 4097 6871 4131
rect 8861 4097 8895 4131
rect 1409 4029 1443 4063
rect 1676 4029 1710 4063
rect 7093 4029 7127 4063
rect 8677 4029 8711 4063
rect 9689 4029 9723 4063
rect 10425 4097 10459 4131
rect 11621 4097 11655 4131
rect 13001 4097 13035 4131
rect 14197 4097 14231 4131
rect 10241 4029 10275 4063
rect 11437 4029 11471 4063
rect 12817 4029 12851 4063
rect 14013 4029 14047 4063
rect 14841 4029 14875 4063
rect 3148 3961 3182 3995
rect 5172 3961 5206 3995
rect 9781 3961 9815 3995
rect 4261 3893 4295 3927
rect 8217 3893 8251 3927
rect 8769 3893 8803 3927
rect 9505 3893 9539 3927
rect 10333 3893 10367 3927
rect 11069 3893 11103 3927
rect 11529 3893 11563 3927
rect 12909 3893 12943 3927
rect 13645 3893 13679 3927
rect 14105 3893 14139 3927
rect 15025 3893 15059 3927
rect 2881 3689 2915 3723
rect 4445 3689 4479 3723
rect 6837 3689 6871 3723
rect 7389 3689 7423 3723
rect 8953 3689 8987 3723
rect 10885 3689 10919 3723
rect 12081 3689 12115 3723
rect 12909 3689 12943 3723
rect 13277 3689 13311 3723
rect 14749 3689 14783 3723
rect 1676 3621 1710 3655
rect 3341 3621 3375 3655
rect 4537 3621 4571 3655
rect 5713 3621 5747 3655
rect 7297 3621 7331 3655
rect 8217 3621 8251 3655
rect 11253 3621 11287 3655
rect 11345 3621 11379 3655
rect 12541 3621 12575 3655
rect 13369 3621 13403 3655
rect 3249 3553 3283 3587
rect 4905 3553 4939 3587
rect 8125 3553 8159 3587
rect 10057 3553 10091 3587
rect 12449 3553 12483 3587
rect 14105 3553 14139 3587
rect 14565 3553 14599 3587
rect 3525 3485 3559 3519
rect 4629 3485 4663 3519
rect 5089 3485 5123 3519
rect 5457 3485 5491 3519
rect 7481 3485 7515 3519
rect 8401 3485 8435 3519
rect 9045 3485 9079 3519
rect 9229 3485 9263 3519
rect 10149 3485 10183 3519
rect 10333 3485 10367 3519
rect 11437 3485 11471 3519
rect 12725 3485 12759 3519
rect 13461 3485 13495 3519
rect 14197 3485 14231 3519
rect 14289 3485 14323 3519
rect 7757 3417 7791 3451
rect 8585 3417 8619 3451
rect 2789 3349 2823 3383
rect 4077 3349 4111 3383
rect 6929 3349 6963 3383
rect 9689 3349 9723 3383
rect 13737 3349 13771 3383
rect 8217 3145 8251 3179
rect 8309 3145 8343 3179
rect 9505 3145 9539 3179
rect 11069 3145 11103 3179
rect 14473 3145 14507 3179
rect 5733 3077 5767 3111
rect 12265 3077 12299 3111
rect 12449 3077 12483 3111
rect 13645 3077 13679 3111
rect 1409 3009 1443 3043
rect 6377 3009 6411 3043
rect 6837 3009 6871 3043
rect 8861 3009 8895 3043
rect 10425 3009 10459 3043
rect 11621 3009 11655 3043
rect 13093 3009 13127 3043
rect 14105 3009 14139 3043
rect 14197 3009 14231 3043
rect 15025 3009 15059 3043
rect 6285 2941 6319 2975
rect 9689 2941 9723 2975
rect 12265 2941 12299 2975
rect 12817 2941 12851 2975
rect 14933 2941 14967 2975
rect 1676 2873 1710 2907
rect 3148 2873 3182 2907
rect 4620 2873 4654 2907
rect 6193 2873 6227 2907
rect 7104 2873 7138 2907
rect 10241 2873 10275 2907
rect 10333 2873 10367 2907
rect 11529 2873 11563 2907
rect 14013 2873 14047 2907
rect 2789 2805 2823 2839
rect 4261 2805 4295 2839
rect 5825 2805 5859 2839
rect 8677 2805 8711 2839
rect 8769 2805 8803 2839
rect 9873 2805 9907 2839
rect 11437 2805 11471 2839
rect 12909 2805 12943 2839
rect 14841 2805 14875 2839
rect 5549 2601 5583 2635
rect 6009 2601 6043 2635
rect 7297 2601 7331 2635
rect 8585 2601 8619 2635
rect 8953 2601 8987 2635
rect 10241 2601 10275 2635
rect 10977 2601 11011 2635
rect 11437 2601 11471 2635
rect 13829 2601 13863 2635
rect 14289 2601 14323 2635
rect 1685 2533 1719 2567
rect 4344 2533 4378 2567
rect 8125 2533 8159 2567
rect 9045 2533 9079 2567
rect 13001 2533 13035 2567
rect 14197 2533 14231 2567
rect 1409 2465 1443 2499
rect 2412 2465 2446 2499
rect 3617 2465 3651 2499
rect 5917 2465 5951 2499
rect 6377 2465 6411 2499
rect 7389 2465 7423 2499
rect 10149 2465 10183 2499
rect 11345 2465 11379 2499
rect 13093 2465 13127 2499
rect 14841 2465 14875 2499
rect 2145 2397 2179 2431
rect 6101 2397 6135 2431
rect 7481 2397 7515 2431
rect 8217 2397 8251 2431
rect 8309 2397 8343 2431
rect 9137 2397 9171 2431
rect 10333 2397 10367 2431
rect 11621 2397 11655 2431
rect 13185 2397 13219 2431
rect 14473 2397 14507 2431
rect 3801 2329 3835 2363
rect 6561 2329 6595 2363
rect 3525 2261 3559 2295
rect 5457 2261 5491 2295
rect 6929 2261 6963 2295
rect 7757 2261 7791 2295
rect 9781 2261 9815 2295
rect 12633 2261 12667 2295
rect 15025 2261 15059 2295
rect 6101 1853 6135 1887
rect 6101 1445 6135 1479
<< metal1 >>
rect 1394 16464 1400 16516
rect 1452 16504 1458 16516
rect 6638 16504 6644 16516
rect 1452 16476 6644 16504
rect 1452 16464 1458 16476
rect 6638 16464 6644 16476
rect 6696 16464 6702 16516
rect 2406 16396 2412 16448
rect 2464 16436 2470 16448
rect 8202 16436 8208 16448
rect 2464 16408 8208 16436
rect 2464 16396 2470 16408
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 1762 16328 1768 16380
rect 1820 16368 1826 16380
rect 10318 16368 10324 16380
rect 1820 16340 10324 16368
rect 1820 16328 1826 16340
rect 10318 16328 10324 16340
rect 10376 16328 10382 16380
rect 4982 16260 4988 16312
rect 5040 16300 5046 16312
rect 10134 16300 10140 16312
rect 5040 16272 10140 16300
rect 5040 16260 5046 16272
rect 10134 16260 10140 16272
rect 10192 16300 10198 16312
rect 11238 16300 11244 16312
rect 10192 16272 11244 16300
rect 10192 16260 10198 16272
rect 11238 16260 11244 16272
rect 11296 16260 11302 16312
rect 4062 16192 4068 16244
rect 4120 16232 4126 16244
rect 8846 16232 8852 16244
rect 4120 16204 8852 16232
rect 4120 16192 4126 16204
rect 8846 16192 8852 16204
rect 8904 16192 8910 16244
rect 198 16124 204 16176
rect 256 16164 262 16176
rect 13722 16164 13728 16176
rect 256 16136 13728 16164
rect 256 16124 262 16136
rect 13722 16124 13728 16136
rect 13780 16124 13786 16176
rect 6362 16056 6368 16108
rect 6420 16096 6426 16108
rect 12618 16096 12624 16108
rect 6420 16068 12624 16096
rect 6420 16056 6426 16068
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 2774 15988 2780 16040
rect 2832 16028 2838 16040
rect 6086 16028 6092 16040
rect 2832 16000 6092 16028
rect 2832 15988 2838 16000
rect 6086 15988 6092 16000
rect 6144 15988 6150 16040
rect 6914 15988 6920 16040
rect 6972 16028 6978 16040
rect 9398 16028 9404 16040
rect 6972 16000 9404 16028
rect 6972 15988 6978 16000
rect 9398 15988 9404 16000
rect 9456 16028 9462 16040
rect 11330 16028 11336 16040
rect 9456 16000 11336 16028
rect 9456 15988 9462 16000
rect 11330 15988 11336 16000
rect 11388 15988 11394 16040
rect 3050 15920 3056 15972
rect 3108 15960 3114 15972
rect 12894 15960 12900 15972
rect 3108 15932 12900 15960
rect 3108 15920 3114 15932
rect 12894 15920 12900 15932
rect 12952 15920 12958 15972
rect 566 15852 572 15904
rect 624 15892 630 15904
rect 14458 15892 14464 15904
rect 624 15864 14464 15892
rect 624 15852 630 15864
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 1104 15802 15824 15824
rect 1104 15750 5912 15802
rect 5964 15750 5976 15802
rect 6028 15750 6040 15802
rect 6092 15750 6104 15802
rect 6156 15750 10843 15802
rect 10895 15750 10907 15802
rect 10959 15750 10971 15802
rect 11023 15750 11035 15802
rect 11087 15750 15824 15802
rect 1104 15728 15824 15750
rect 1581 15691 1639 15697
rect 1581 15657 1593 15691
rect 1627 15688 1639 15691
rect 2682 15688 2688 15700
rect 1627 15660 2688 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 2682 15648 2688 15660
rect 2740 15648 2746 15700
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 5721 15691 5779 15697
rect 5721 15688 5733 15691
rect 4212 15660 5733 15688
rect 4212 15648 4218 15660
rect 5721 15657 5733 15660
rect 5767 15657 5779 15691
rect 5721 15651 5779 15657
rect 6546 15648 6552 15700
rect 6604 15688 6610 15700
rect 9953 15691 10011 15697
rect 9953 15688 9965 15691
rect 6604 15660 9965 15688
rect 6604 15648 6610 15660
rect 9953 15657 9965 15660
rect 9999 15657 10011 15691
rect 9953 15651 10011 15657
rect 10318 15648 10324 15700
rect 10376 15688 10382 15700
rect 10965 15691 11023 15697
rect 10965 15688 10977 15691
rect 10376 15660 10977 15688
rect 10376 15648 10382 15660
rect 10965 15657 10977 15660
rect 11011 15657 11023 15691
rect 13722 15688 13728 15700
rect 13683 15660 13728 15688
rect 10965 15651 11023 15657
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 14458 15688 14464 15700
rect 14419 15660 14464 15688
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 4801 15623 4859 15629
rect 4801 15589 4813 15623
rect 4847 15620 4859 15623
rect 4982 15620 4988 15632
rect 4847 15592 4988 15620
rect 4847 15589 4859 15592
rect 4801 15583 4859 15589
rect 4982 15580 4988 15592
rect 5040 15580 5046 15632
rect 7285 15623 7343 15629
rect 7285 15589 7297 15623
rect 7331 15620 7343 15623
rect 8294 15620 8300 15632
rect 7331 15592 8300 15620
rect 7331 15589 7343 15592
rect 7285 15583 7343 15589
rect 8294 15580 8300 15592
rect 8352 15580 8358 15632
rect 8481 15623 8539 15629
rect 8481 15620 8493 15623
rect 8404 15592 8493 15620
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 2222 15552 2228 15564
rect 1443 15524 2228 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 2222 15512 2228 15524
rect 2280 15512 2286 15564
rect 2400 15555 2458 15561
rect 2400 15521 2412 15555
rect 2446 15552 2458 15555
rect 2866 15552 2872 15564
rect 2446 15524 2872 15552
rect 2446 15521 2458 15524
rect 2400 15515 2458 15521
rect 2866 15512 2872 15524
rect 2924 15552 2930 15564
rect 4062 15552 4068 15564
rect 2924 15524 4068 15552
rect 2924 15512 2930 15524
rect 4062 15512 4068 15524
rect 4120 15512 4126 15564
rect 4706 15552 4712 15564
rect 4667 15524 4712 15552
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 5537 15555 5595 15561
rect 5537 15521 5549 15555
rect 5583 15552 5595 15555
rect 7190 15552 7196 15564
rect 5583 15524 7196 15552
rect 5583 15521 5595 15524
rect 5537 15515 5595 15521
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 7377 15555 7435 15561
rect 7377 15521 7389 15555
rect 7423 15552 7435 15555
rect 7423 15524 7604 15552
rect 7423 15521 7435 15524
rect 7377 15515 7435 15521
rect 2130 15484 2136 15496
rect 2091 15456 2136 15484
rect 2130 15444 2136 15456
rect 2188 15444 2194 15496
rect 4982 15484 4988 15496
rect 4943 15456 4988 15484
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 6730 15484 6736 15496
rect 5460 15456 6736 15484
rect 4341 15419 4399 15425
rect 4341 15416 4353 15419
rect 3068 15388 4353 15416
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 3068 15348 3096 15388
rect 4341 15385 4353 15388
rect 4387 15385 4399 15419
rect 5460 15416 5488 15456
rect 6730 15444 6736 15456
rect 6788 15484 6794 15496
rect 7469 15487 7527 15493
rect 7469 15484 7481 15487
rect 6788 15456 7481 15484
rect 6788 15444 6794 15456
rect 7469 15453 7481 15456
rect 7515 15453 7527 15487
rect 7576 15484 7604 15524
rect 7650 15512 7656 15564
rect 7708 15552 7714 15564
rect 8404 15552 8432 15592
rect 8481 15589 8493 15592
rect 8527 15589 8539 15623
rect 8481 15583 8539 15589
rect 8662 15580 8668 15632
rect 8720 15620 8726 15632
rect 9582 15620 9588 15632
rect 8720 15592 9588 15620
rect 8720 15580 8726 15592
rect 9582 15580 9588 15592
rect 9640 15580 9646 15632
rect 12158 15580 12164 15632
rect 12216 15620 12222 15632
rect 12894 15620 12900 15632
rect 12216 15592 12756 15620
rect 12855 15592 12900 15620
rect 12216 15580 12222 15592
rect 8573 15555 8631 15561
rect 8573 15552 8585 15555
rect 7708 15524 8432 15552
rect 8496 15524 8585 15552
rect 7708 15512 7714 15524
rect 8386 15484 8392 15496
rect 7576 15456 8392 15484
rect 7469 15447 7527 15453
rect 8386 15444 8392 15456
rect 8444 15444 8450 15496
rect 4341 15379 4399 15385
rect 4448 15388 5488 15416
rect 2832 15320 3096 15348
rect 3513 15351 3571 15357
rect 2832 15308 2838 15320
rect 3513 15317 3525 15351
rect 3559 15348 3571 15351
rect 4448 15348 4476 15388
rect 5534 15376 5540 15428
rect 5592 15416 5598 15428
rect 8496 15416 8524 15524
rect 8573 15521 8585 15524
rect 8619 15521 8631 15555
rect 8573 15515 8631 15521
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 9769 15555 9827 15561
rect 9769 15552 9781 15555
rect 9732 15524 9781 15552
rect 9732 15512 9738 15524
rect 9769 15521 9781 15524
rect 9815 15521 9827 15555
rect 9769 15515 9827 15521
rect 11333 15555 11391 15561
rect 11333 15521 11345 15555
rect 11379 15552 11391 15555
rect 11974 15552 11980 15564
rect 11379 15524 11980 15552
rect 11379 15521 11391 15524
rect 11333 15515 11391 15521
rect 11974 15512 11980 15524
rect 12032 15512 12038 15564
rect 12618 15552 12624 15564
rect 12579 15524 12624 15552
rect 12618 15512 12624 15524
rect 12676 15512 12682 15564
rect 12728 15552 12756 15592
rect 12894 15580 12900 15592
rect 12952 15580 12958 15632
rect 13541 15555 13599 15561
rect 13541 15552 13553 15555
rect 12728 15524 13553 15552
rect 13541 15521 13553 15524
rect 13587 15521 13599 15555
rect 13541 15515 13599 15521
rect 14277 15555 14335 15561
rect 14277 15521 14289 15555
rect 14323 15521 14335 15555
rect 14277 15515 14335 15521
rect 8665 15487 8723 15493
rect 8665 15453 8677 15487
rect 8711 15453 8723 15487
rect 8665 15447 8723 15453
rect 11425 15487 11483 15493
rect 11425 15453 11437 15487
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15484 11667 15487
rect 13722 15484 13728 15496
rect 11655 15456 13728 15484
rect 11655 15453 11667 15456
rect 11609 15447 11667 15453
rect 5592 15388 8524 15416
rect 8680 15416 8708 15447
rect 9306 15416 9312 15428
rect 8680 15388 9312 15416
rect 5592 15376 5598 15388
rect 9306 15376 9312 15388
rect 9364 15376 9370 15428
rect 11440 15416 11468 15447
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 12250 15416 12256 15428
rect 11440 15388 12256 15416
rect 12250 15376 12256 15388
rect 12308 15376 12314 15428
rect 3559 15320 4476 15348
rect 3559 15317 3571 15320
rect 3513 15311 3571 15317
rect 4522 15308 4528 15360
rect 4580 15348 4586 15360
rect 6917 15351 6975 15357
rect 6917 15348 6929 15351
rect 4580 15320 6929 15348
rect 4580 15308 4586 15320
rect 6917 15317 6929 15320
rect 6963 15317 6975 15351
rect 6917 15311 6975 15317
rect 8113 15351 8171 15357
rect 8113 15317 8125 15351
rect 8159 15348 8171 15351
rect 11238 15348 11244 15360
rect 8159 15320 11244 15348
rect 8159 15317 8171 15320
rect 8113 15311 8171 15317
rect 11238 15308 11244 15320
rect 11296 15308 11302 15360
rect 13630 15308 13636 15360
rect 13688 15348 13694 15360
rect 14292 15348 14320 15515
rect 13688 15320 14320 15348
rect 13688 15308 13694 15320
rect 1104 15258 15824 15280
rect 1104 15206 3447 15258
rect 3499 15206 3511 15258
rect 3563 15206 3575 15258
rect 3627 15206 3639 15258
rect 3691 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 13308 15258
rect 13360 15206 13372 15258
rect 13424 15206 13436 15258
rect 13488 15206 13500 15258
rect 13552 15206 15824 15258
rect 1104 15184 15824 15206
rect 1673 15147 1731 15153
rect 1673 15113 1685 15147
rect 1719 15144 1731 15147
rect 2314 15144 2320 15156
rect 1719 15116 2320 15144
rect 1719 15113 1731 15116
rect 1673 15107 1731 15113
rect 2314 15104 2320 15116
rect 2372 15104 2378 15156
rect 4801 15147 4859 15153
rect 4801 15113 4813 15147
rect 4847 15144 4859 15147
rect 5166 15144 5172 15156
rect 4847 15116 5172 15144
rect 4847 15113 4859 15116
rect 4801 15107 4859 15113
rect 5166 15104 5172 15116
rect 5224 15104 5230 15156
rect 5258 15104 5264 15156
rect 5316 15144 5322 15156
rect 6181 15147 6239 15153
rect 6181 15144 6193 15147
rect 5316 15116 6193 15144
rect 5316 15104 5322 15116
rect 6181 15113 6193 15116
rect 6227 15113 6239 15147
rect 6181 15107 6239 15113
rect 7374 15104 7380 15156
rect 7432 15144 7438 15156
rect 8021 15147 8079 15153
rect 8021 15144 8033 15147
rect 7432 15116 8033 15144
rect 7432 15104 7438 15116
rect 8021 15113 8033 15116
rect 8067 15113 8079 15147
rect 8021 15107 8079 15113
rect 8573 15147 8631 15153
rect 8573 15113 8585 15147
rect 8619 15144 8631 15147
rect 8662 15144 8668 15156
rect 8619 15116 8668 15144
rect 8619 15113 8631 15116
rect 8573 15107 8631 15113
rect 8662 15104 8668 15116
rect 8720 15104 8726 15156
rect 9953 15147 10011 15153
rect 9953 15144 9965 15147
rect 8763 15116 9965 15144
rect 1854 15036 1860 15088
rect 1912 15076 1918 15088
rect 2961 15079 3019 15085
rect 2961 15076 2973 15079
rect 1912 15048 2973 15076
rect 1912 15036 1918 15048
rect 2961 15045 2973 15048
rect 3007 15045 3019 15079
rect 2961 15039 3019 15045
rect 5718 15036 5724 15088
rect 5776 15076 5782 15088
rect 8763 15076 8791 15116
rect 9953 15113 9965 15116
rect 9999 15113 10011 15147
rect 9953 15107 10011 15113
rect 11146 15104 11152 15156
rect 11204 15144 11210 15156
rect 15470 15144 15476 15156
rect 11204 15116 15476 15144
rect 11204 15104 11210 15116
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 5776 15048 8791 15076
rect 5776 15036 5782 15048
rect 8938 15036 8944 15088
rect 8996 15076 9002 15088
rect 13538 15076 13544 15088
rect 8996 15048 13544 15076
rect 8996 15036 9002 15048
rect 13538 15036 13544 15048
rect 13596 15036 13602 15088
rect 13817 15079 13875 15085
rect 13817 15076 13829 15079
rect 13740 15048 13829 15076
rect 4062 15008 4068 15020
rect 4023 14980 4068 15008
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 4246 15008 4252 15020
rect 4207 14980 4252 15008
rect 4246 14968 4252 14980
rect 4304 14968 4310 15020
rect 4890 15008 4896 15020
rect 4724 14980 4896 15008
rect 1486 14940 1492 14952
rect 1447 14912 1492 14940
rect 1486 14900 1492 14912
rect 1544 14900 1550 14952
rect 2777 14943 2835 14949
rect 2777 14909 2789 14943
rect 2823 14940 2835 14943
rect 4724 14940 4752 14980
rect 4890 14968 4896 14980
rect 4948 14968 4954 15020
rect 5442 15008 5448 15020
rect 5403 14980 5448 15008
rect 5442 14968 5448 14980
rect 5500 15008 5506 15020
rect 7742 15008 7748 15020
rect 5500 14980 7748 15008
rect 5500 14968 5506 14980
rect 7742 14968 7748 14980
rect 7800 14968 7806 15020
rect 9214 15008 9220 15020
rect 9175 14980 9220 15008
rect 9214 14968 9220 14980
rect 9272 14968 9278 15020
rect 11698 15008 11704 15020
rect 9600 14980 11560 15008
rect 11659 14980 11704 15008
rect 2823 14912 4752 14940
rect 2823 14909 2835 14912
rect 2777 14903 2835 14909
rect 4798 14900 4804 14952
rect 4856 14940 4862 14952
rect 5997 14943 6055 14949
rect 4856 14912 5856 14940
rect 4856 14900 4862 14912
rect 5261 14875 5319 14881
rect 5261 14841 5273 14875
rect 5307 14872 5319 14875
rect 5626 14872 5632 14884
rect 5307 14844 5632 14872
rect 5307 14841 5319 14844
rect 5261 14835 5319 14841
rect 5626 14832 5632 14844
rect 5684 14832 5690 14884
rect 3602 14804 3608 14816
rect 3563 14776 3608 14804
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 3970 14804 3976 14816
rect 3931 14776 3976 14804
rect 3970 14764 3976 14776
rect 4028 14764 4034 14816
rect 5169 14807 5227 14813
rect 5169 14773 5181 14807
rect 5215 14804 5227 14807
rect 5718 14804 5724 14816
rect 5215 14776 5724 14804
rect 5215 14773 5227 14776
rect 5169 14767 5227 14773
rect 5718 14764 5724 14776
rect 5776 14764 5782 14816
rect 5828 14804 5856 14912
rect 5997 14909 6009 14943
rect 6043 14909 6055 14943
rect 5997 14903 6055 14909
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14940 6883 14943
rect 7282 14940 7288 14952
rect 6871 14912 7288 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 6012 14872 6040 14903
rect 7282 14900 7288 14912
rect 7340 14900 7346 14952
rect 7837 14943 7895 14949
rect 7837 14909 7849 14943
rect 7883 14940 7895 14943
rect 9600 14940 9628 14980
rect 7883 14912 9628 14940
rect 9769 14943 9827 14949
rect 7883 14909 7895 14912
rect 7837 14903 7895 14909
rect 9769 14909 9781 14943
rect 9815 14940 9827 14943
rect 10318 14940 10324 14952
rect 9815 14912 10324 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 10318 14900 10324 14912
rect 10376 14900 10382 14952
rect 10502 14900 10508 14952
rect 10560 14940 10566 14952
rect 11425 14943 11483 14949
rect 11425 14940 11437 14943
rect 10560 14912 11437 14940
rect 10560 14900 10566 14912
rect 11425 14909 11437 14912
rect 11471 14909 11483 14943
rect 11532 14940 11560 14980
rect 11698 14968 11704 14980
rect 11756 15008 11762 15020
rect 12894 15008 12900 15020
rect 11756 14980 12900 15008
rect 11756 14968 11762 14980
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 13078 15008 13084 15020
rect 13039 14980 13084 15008
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 12342 14940 12348 14952
rect 11532 14912 12348 14940
rect 11425 14903 11483 14909
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 12986 14900 12992 14952
rect 13044 14940 13050 14952
rect 13633 14943 13691 14949
rect 13633 14940 13645 14943
rect 13044 14912 13645 14940
rect 13044 14900 13050 14912
rect 13633 14909 13645 14912
rect 13679 14909 13691 14943
rect 13633 14903 13691 14909
rect 8754 14872 8760 14884
rect 6012 14844 8760 14872
rect 8754 14832 8760 14844
rect 8812 14832 8818 14884
rect 9033 14875 9091 14881
rect 9033 14841 9045 14875
rect 9079 14872 9091 14875
rect 11146 14872 11152 14884
rect 9079 14844 11152 14872
rect 9079 14841 9091 14844
rect 9033 14835 9091 14841
rect 11146 14832 11152 14844
rect 11204 14832 11210 14884
rect 12066 14832 12072 14884
rect 12124 14872 12130 14884
rect 13740 14872 13768 15048
rect 13817 15045 13829 15048
rect 13863 15045 13875 15079
rect 13817 15039 13875 15045
rect 13998 14900 14004 14952
rect 14056 14940 14062 14952
rect 14369 14943 14427 14949
rect 14369 14940 14381 14943
rect 14056 14912 14381 14940
rect 14056 14900 14062 14912
rect 14369 14909 14381 14912
rect 14415 14909 14427 14943
rect 14369 14903 14427 14909
rect 15102 14872 15108 14884
rect 12124 14844 13768 14872
rect 13924 14844 15108 14872
rect 12124 14832 12130 14844
rect 7009 14807 7067 14813
rect 7009 14804 7021 14807
rect 5828 14776 7021 14804
rect 7009 14773 7021 14776
rect 7055 14773 7067 14807
rect 7009 14767 7067 14773
rect 7374 14764 7380 14816
rect 7432 14804 7438 14816
rect 8941 14807 8999 14813
rect 8941 14804 8953 14807
rect 7432 14776 8953 14804
rect 7432 14764 7438 14776
rect 8941 14773 8953 14776
rect 8987 14773 8999 14807
rect 8941 14767 8999 14773
rect 9214 14764 9220 14816
rect 9272 14804 9278 14816
rect 10686 14804 10692 14816
rect 9272 14776 10692 14804
rect 9272 14764 9278 14776
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 11057 14807 11115 14813
rect 11057 14773 11069 14807
rect 11103 14804 11115 14807
rect 11422 14804 11428 14816
rect 11103 14776 11428 14804
rect 11103 14773 11115 14776
rect 11057 14767 11115 14773
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 11517 14807 11575 14813
rect 11517 14773 11529 14807
rect 11563 14804 11575 14807
rect 11790 14804 11796 14816
rect 11563 14776 11796 14804
rect 11563 14773 11575 14776
rect 11517 14767 11575 14773
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 12434 14804 12440 14816
rect 12395 14776 12440 14804
rect 12434 14764 12440 14776
rect 12492 14764 12498 14816
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 12805 14807 12863 14813
rect 12805 14804 12817 14807
rect 12676 14776 12817 14804
rect 12676 14764 12682 14776
rect 12805 14773 12817 14776
rect 12851 14773 12863 14807
rect 12805 14767 12863 14773
rect 12897 14807 12955 14813
rect 12897 14773 12909 14807
rect 12943 14804 12955 14807
rect 13924 14804 13952 14844
rect 15102 14832 15108 14844
rect 15160 14872 15166 14884
rect 16298 14872 16304 14884
rect 15160 14844 16304 14872
rect 15160 14832 15166 14844
rect 16298 14832 16304 14844
rect 16356 14832 16362 14884
rect 14550 14804 14556 14816
rect 12943 14776 13952 14804
rect 14511 14776 14556 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 1104 14714 15824 14736
rect 1104 14662 5912 14714
rect 5964 14662 5976 14714
rect 6028 14662 6040 14714
rect 6092 14662 6104 14714
rect 6156 14662 10843 14714
rect 10895 14662 10907 14714
rect 10959 14662 10971 14714
rect 11023 14662 11035 14714
rect 11087 14662 15824 14714
rect 1104 14640 15824 14662
rect 1949 14603 2007 14609
rect 1949 14569 1961 14603
rect 1995 14600 2007 14603
rect 3326 14600 3332 14612
rect 1995 14572 3332 14600
rect 1995 14569 2007 14572
rect 1949 14563 2007 14569
rect 3326 14560 3332 14572
rect 3384 14560 3390 14612
rect 3421 14603 3479 14609
rect 3421 14569 3433 14603
rect 3467 14600 3479 14603
rect 3513 14603 3571 14609
rect 3513 14600 3525 14603
rect 3467 14572 3525 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 3513 14569 3525 14572
rect 3559 14569 3571 14603
rect 3513 14563 3571 14569
rect 3602 14560 3608 14612
rect 3660 14600 3666 14612
rect 3660 14572 4568 14600
rect 3660 14560 3666 14572
rect 2130 14492 2136 14544
rect 2188 14532 2194 14544
rect 2777 14535 2835 14541
rect 2188 14504 2728 14532
rect 2188 14492 2194 14504
rect 1765 14467 1823 14473
rect 1765 14433 1777 14467
rect 1811 14433 1823 14467
rect 2498 14464 2504 14476
rect 2459 14436 2504 14464
rect 1765 14427 1823 14433
rect 1780 14396 1808 14427
rect 2498 14424 2504 14436
rect 2556 14424 2562 14476
rect 2700 14464 2728 14504
rect 2777 14501 2789 14535
rect 2823 14532 2835 14535
rect 3878 14532 3884 14544
rect 2823 14504 3884 14532
rect 2823 14501 2835 14504
rect 2777 14495 2835 14501
rect 3878 14492 3884 14504
rect 3936 14492 3942 14544
rect 4540 14532 4568 14572
rect 5166 14560 5172 14612
rect 5224 14600 5230 14612
rect 6362 14600 6368 14612
rect 5224 14572 6368 14600
rect 5224 14560 5230 14572
rect 6362 14560 6368 14572
rect 6420 14560 6426 14612
rect 6549 14603 6607 14609
rect 6549 14569 6561 14603
rect 6595 14600 6607 14603
rect 7466 14600 7472 14612
rect 6595 14572 7472 14600
rect 6595 14569 6607 14572
rect 6549 14563 6607 14569
rect 7466 14560 7472 14572
rect 7524 14560 7530 14612
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 7745 14603 7803 14609
rect 7745 14600 7757 14603
rect 7708 14572 7757 14600
rect 7708 14560 7714 14572
rect 7745 14569 7757 14572
rect 7791 14569 7803 14603
rect 7745 14563 7803 14569
rect 7926 14560 7932 14612
rect 7984 14600 7990 14612
rect 7984 14572 11100 14600
rect 7984 14560 7990 14572
rect 6454 14532 6460 14544
rect 4540 14504 6460 14532
rect 6454 14492 6460 14504
rect 6512 14492 6518 14544
rect 7098 14492 7104 14544
rect 7156 14532 7162 14544
rect 7156 14504 7788 14532
rect 7156 14492 7162 14504
rect 3421 14467 3479 14473
rect 3421 14464 3433 14467
rect 2700 14436 3433 14464
rect 3421 14433 3433 14436
rect 3467 14433 3479 14467
rect 3421 14427 3479 14433
rect 3697 14467 3755 14473
rect 3697 14433 3709 14467
rect 3743 14464 3755 14467
rect 3786 14464 3792 14476
rect 3743 14436 3792 14464
rect 3743 14433 3755 14436
rect 3697 14427 3755 14433
rect 2958 14396 2964 14408
rect 1780 14368 2964 14396
rect 2958 14356 2964 14368
rect 3016 14356 3022 14408
rect 3436 14396 3464 14427
rect 3786 14424 3792 14436
rect 3844 14424 3850 14476
rect 4246 14424 4252 14476
rect 4304 14464 4310 14476
rect 4597 14467 4655 14473
rect 4597 14464 4609 14467
rect 4304 14436 4609 14464
rect 4304 14424 4310 14436
rect 4597 14433 4609 14436
rect 4643 14433 4655 14467
rect 7760 14464 7788 14504
rect 8110 14492 8116 14544
rect 8168 14532 8174 14544
rect 8846 14532 8852 14544
rect 8168 14504 8708 14532
rect 8807 14504 8852 14532
rect 8168 14492 8174 14504
rect 7837 14467 7895 14473
rect 7837 14464 7849 14467
rect 7760 14436 7849 14464
rect 4597 14427 4655 14433
rect 7837 14433 7849 14436
rect 7883 14433 7895 14467
rect 7837 14427 7895 14433
rect 8202 14424 8208 14476
rect 8260 14464 8266 14476
rect 8573 14467 8631 14473
rect 8573 14464 8585 14467
rect 8260 14436 8585 14464
rect 8260 14424 8266 14436
rect 8573 14433 8585 14436
rect 8619 14433 8631 14467
rect 8680 14464 8708 14504
rect 8846 14492 8852 14504
rect 8904 14492 8910 14544
rect 10042 14532 10048 14544
rect 9784 14504 10048 14532
rect 9784 14464 9812 14504
rect 10042 14492 10048 14504
rect 10100 14492 10106 14544
rect 9950 14473 9956 14476
rect 9944 14464 9956 14473
rect 8680 14436 9812 14464
rect 9911 14436 9956 14464
rect 8573 14427 8631 14433
rect 9944 14427 9956 14436
rect 9950 14424 9956 14427
rect 10008 14424 10014 14476
rect 10226 14424 10232 14476
rect 10284 14464 10290 14476
rect 10502 14464 10508 14476
rect 10284 14436 10508 14464
rect 10284 14424 10290 14436
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 11072 14464 11100 14572
rect 11422 14560 11428 14612
rect 11480 14600 11486 14612
rect 12437 14603 12495 14609
rect 12437 14600 12449 14603
rect 11480 14572 12449 14600
rect 11480 14560 11486 14572
rect 12437 14569 12449 14572
rect 12483 14569 12495 14603
rect 12437 14563 12495 14569
rect 12529 14603 12587 14609
rect 12529 14569 12541 14603
rect 12575 14600 12587 14603
rect 13078 14600 13084 14612
rect 12575 14572 13084 14600
rect 12575 14569 12587 14572
rect 12529 14563 12587 14569
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 11790 14492 11796 14544
rect 11848 14532 11854 14544
rect 13538 14532 13544 14544
rect 11848 14504 13400 14532
rect 13499 14504 13544 14532
rect 11848 14492 11854 14504
rect 12066 14464 12072 14476
rect 11072 14436 12072 14464
rect 12066 14424 12072 14436
rect 12124 14424 12130 14476
rect 13262 14464 13268 14476
rect 13223 14436 13268 14464
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 13372 14464 13400 14504
rect 13538 14492 13544 14504
rect 13596 14492 13602 14544
rect 14185 14467 14243 14473
rect 14185 14464 14197 14467
rect 13372 14436 14197 14464
rect 14185 14433 14197 14436
rect 14231 14464 14243 14467
rect 16758 14464 16764 14476
rect 14231 14436 16764 14464
rect 14231 14433 14243 14436
rect 14185 14427 14243 14433
rect 16758 14424 16764 14436
rect 16816 14424 16822 14476
rect 4338 14396 4344 14408
rect 3436 14368 4344 14396
rect 4338 14356 4344 14368
rect 4396 14356 4402 14408
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 6641 14399 6699 14405
rect 6641 14396 6653 14399
rect 5408 14368 6653 14396
rect 5408 14356 5414 14368
rect 6641 14365 6653 14368
rect 6687 14365 6699 14399
rect 6641 14359 6699 14365
rect 6730 14356 6736 14408
rect 6788 14396 6794 14408
rect 8021 14399 8079 14405
rect 6788 14368 6833 14396
rect 6788 14356 6794 14368
rect 8021 14365 8033 14399
rect 8067 14396 8079 14399
rect 8294 14396 8300 14408
rect 8067 14368 8300 14396
rect 8067 14365 8079 14368
rect 8021 14359 8079 14365
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 9674 14396 9680 14408
rect 8536 14368 9680 14396
rect 8536 14356 8542 14368
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 12710 14396 12716 14408
rect 12671 14368 12716 14396
rect 12710 14356 12716 14368
rect 12768 14356 12774 14408
rect 12802 14356 12808 14408
rect 12860 14396 12866 14408
rect 14090 14396 14096 14408
rect 12860 14368 14096 14396
rect 12860 14356 12866 14368
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 5721 14331 5779 14337
rect 5721 14297 5733 14331
rect 5767 14328 5779 14331
rect 6086 14328 6092 14340
rect 5767 14300 6092 14328
rect 5767 14297 5779 14300
rect 5721 14291 5779 14297
rect 6086 14288 6092 14300
rect 6144 14288 6150 14340
rect 6178 14288 6184 14340
rect 6236 14328 6242 14340
rect 9214 14328 9220 14340
rect 6236 14300 6281 14328
rect 6472 14300 7880 14328
rect 6236 14288 6242 14300
rect 3326 14220 3332 14272
rect 3384 14260 3390 14272
rect 6472 14260 6500 14300
rect 3384 14232 6500 14260
rect 3384 14220 3390 14232
rect 6546 14220 6552 14272
rect 6604 14260 6610 14272
rect 7377 14263 7435 14269
rect 7377 14260 7389 14263
rect 6604 14232 7389 14260
rect 6604 14220 6610 14232
rect 7377 14229 7389 14232
rect 7423 14229 7435 14263
rect 7852 14260 7880 14300
rect 8036 14300 9220 14328
rect 8036 14260 8064 14300
rect 9214 14288 9220 14300
rect 9272 14288 9278 14340
rect 11974 14288 11980 14340
rect 12032 14328 12038 14340
rect 12069 14331 12127 14337
rect 12069 14328 12081 14331
rect 12032 14300 12081 14328
rect 12032 14288 12038 14300
rect 12069 14297 12081 14300
rect 12115 14297 12127 14331
rect 12069 14291 12127 14297
rect 7852 14232 8064 14260
rect 7377 14223 7435 14229
rect 10686 14220 10692 14272
rect 10744 14260 10750 14272
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 10744 14232 11069 14260
rect 10744 14220 10750 14232
rect 11057 14229 11069 14232
rect 11103 14260 11115 14263
rect 11330 14260 11336 14272
rect 11103 14232 11336 14260
rect 11103 14229 11115 14232
rect 11057 14223 11115 14229
rect 11330 14220 11336 14232
rect 11388 14220 11394 14272
rect 11422 14220 11428 14272
rect 11480 14260 11486 14272
rect 12802 14260 12808 14272
rect 11480 14232 12808 14260
rect 11480 14220 11486 14232
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 14366 14260 14372 14272
rect 14327 14232 14372 14260
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 1104 14170 15824 14192
rect 1104 14118 3447 14170
rect 3499 14118 3511 14170
rect 3563 14118 3575 14170
rect 3627 14118 3639 14170
rect 3691 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 13308 14170
rect 13360 14118 13372 14170
rect 13424 14118 13436 14170
rect 13488 14118 13500 14170
rect 13552 14118 15824 14170
rect 1104 14096 15824 14118
rect 2406 14016 2412 14068
rect 2464 14056 2470 14068
rect 2501 14059 2559 14065
rect 2501 14056 2513 14059
rect 2464 14028 2513 14056
rect 2464 14016 2470 14028
rect 2501 14025 2513 14028
rect 2547 14025 2559 14059
rect 2501 14019 2559 14025
rect 3237 14059 3295 14065
rect 3237 14025 3249 14059
rect 3283 14056 3295 14059
rect 3786 14056 3792 14068
rect 3283 14028 3792 14056
rect 3283 14025 3295 14028
rect 3237 14019 3295 14025
rect 3786 14016 3792 14028
rect 3844 14056 3850 14068
rect 5626 14056 5632 14068
rect 3844 14028 5632 14056
rect 3844 14016 3850 14028
rect 5626 14016 5632 14028
rect 5684 14016 5690 14068
rect 6362 14016 6368 14068
rect 6420 14056 6426 14068
rect 6914 14056 6920 14068
rect 6420 14028 6920 14056
rect 6420 14016 6426 14028
rect 6914 14016 6920 14028
rect 6972 14016 6978 14068
rect 7285 14059 7343 14065
rect 7285 14025 7297 14059
rect 7331 14056 7343 14059
rect 7558 14056 7564 14068
rect 7331 14028 7564 14056
rect 7331 14025 7343 14028
rect 7285 14019 7343 14025
rect 7558 14016 7564 14028
rect 7616 14016 7622 14068
rect 7650 14016 7656 14068
rect 7708 14056 7714 14068
rect 10321 14059 10379 14065
rect 10321 14056 10333 14059
rect 7708 14028 10333 14056
rect 7708 14016 7714 14028
rect 10321 14025 10333 14028
rect 10367 14025 10379 14059
rect 10321 14019 10379 14025
rect 10502 14016 10508 14068
rect 10560 14056 10566 14068
rect 10560 14028 14872 14056
rect 10560 14016 10566 14028
rect 1765 13991 1823 13997
rect 1765 13957 1777 13991
rect 1811 13988 1823 13991
rect 3050 13988 3056 14000
rect 1811 13960 3056 13988
rect 1811 13957 1823 13960
rect 1765 13951 1823 13957
rect 3050 13948 3056 13960
rect 3108 13948 3114 14000
rect 4157 13991 4215 13997
rect 4157 13957 4169 13991
rect 4203 13988 4215 13991
rect 5166 13988 5172 14000
rect 4203 13960 5172 13988
rect 4203 13957 4215 13960
rect 4157 13951 4215 13957
rect 5166 13948 5172 13960
rect 5224 13948 5230 14000
rect 5353 13991 5411 13997
rect 5353 13957 5365 13991
rect 5399 13988 5411 13991
rect 6822 13988 6828 14000
rect 5399 13960 6828 13988
rect 5399 13957 5411 13960
rect 5353 13951 5411 13957
rect 6822 13948 6828 13960
rect 6880 13948 6886 14000
rect 7466 13948 7472 14000
rect 7524 13988 7530 14000
rect 8018 13988 8024 14000
rect 7524 13960 8024 13988
rect 7524 13948 7530 13960
rect 8018 13948 8024 13960
rect 8076 13988 8082 14000
rect 9858 13988 9864 14000
rect 8076 13960 8432 13988
rect 9819 13960 9864 13988
rect 8076 13948 8082 13960
rect 4614 13920 4620 13932
rect 2332 13892 4620 13920
rect 1581 13855 1639 13861
rect 1581 13821 1593 13855
rect 1627 13852 1639 13855
rect 1670 13852 1676 13864
rect 1627 13824 1676 13852
rect 1627 13821 1639 13824
rect 1581 13815 1639 13821
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 2332 13861 2360 13892
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 4798 13920 4804 13932
rect 4759 13892 4804 13920
rect 4798 13880 4804 13892
rect 4856 13880 4862 13932
rect 5534 13880 5540 13932
rect 5592 13920 5598 13932
rect 5813 13923 5871 13929
rect 5813 13920 5825 13923
rect 5592 13892 5825 13920
rect 5592 13880 5598 13892
rect 5813 13889 5825 13892
rect 5859 13889 5871 13923
rect 5813 13883 5871 13889
rect 5902 13880 5908 13932
rect 5960 13920 5966 13932
rect 5960 13892 6005 13920
rect 5960 13880 5966 13892
rect 7190 13880 7196 13932
rect 7248 13920 7254 13932
rect 7248 13892 7696 13920
rect 7248 13880 7254 13892
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13821 2375 13855
rect 2317 13815 2375 13821
rect 3326 13812 3332 13864
rect 3384 13852 3390 13864
rect 3421 13855 3479 13861
rect 3421 13852 3433 13855
rect 3384 13824 3433 13852
rect 3384 13812 3390 13824
rect 3421 13821 3433 13824
rect 3467 13821 3479 13855
rect 6178 13852 6184 13864
rect 3421 13815 3479 13821
rect 4632 13824 6184 13852
rect 4522 13784 4528 13796
rect 4483 13756 4528 13784
rect 4522 13744 4528 13756
rect 4580 13744 4586 13796
rect 4632 13793 4660 13824
rect 6178 13812 6184 13824
rect 6236 13812 6242 13864
rect 6638 13812 6644 13864
rect 6696 13852 6702 13864
rect 7558 13852 7564 13864
rect 6696 13824 7564 13852
rect 6696 13812 6702 13824
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 7668 13861 7696 13892
rect 7742 13880 7748 13932
rect 7800 13920 7806 13932
rect 7929 13923 7987 13929
rect 7929 13920 7941 13923
rect 7800 13892 7941 13920
rect 7800 13880 7806 13892
rect 7929 13889 7941 13892
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 7653 13855 7711 13861
rect 7653 13821 7665 13855
rect 7699 13852 7711 13855
rect 7834 13852 7840 13864
rect 7699 13824 7840 13852
rect 7699 13821 7711 13824
rect 7653 13815 7711 13821
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 8404 13852 8432 13960
rect 9858 13948 9864 13960
rect 9916 13988 9922 14000
rect 12710 13988 12716 14000
rect 9916 13960 12716 13988
rect 9916 13948 9922 13960
rect 12710 13948 12716 13960
rect 12768 13988 12774 14000
rect 12768 13960 13032 13988
rect 12768 13948 12774 13960
rect 9766 13880 9772 13932
rect 9824 13920 9830 13932
rect 10873 13923 10931 13929
rect 10873 13920 10885 13923
rect 9824 13892 10885 13920
rect 9824 13880 9830 13892
rect 10873 13889 10885 13892
rect 10919 13889 10931 13923
rect 10873 13883 10931 13889
rect 11238 13880 11244 13932
rect 11296 13920 11302 13932
rect 13004 13929 13032 13960
rect 12897 13923 12955 13929
rect 12897 13920 12909 13923
rect 11296 13892 12909 13920
rect 11296 13880 11302 13892
rect 12897 13889 12909 13892
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 12989 13923 13047 13929
rect 12989 13889 13001 13923
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 13170 13880 13176 13932
rect 13228 13920 13234 13932
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 13228 13892 14197 13920
rect 13228 13880 13234 13892
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14844 13861 14872 14028
rect 15010 13988 15016 14000
rect 14971 13960 15016 13988
rect 15010 13948 15016 13960
rect 15068 13948 15074 14000
rect 8481 13855 8539 13861
rect 8481 13852 8493 13855
rect 8404 13824 8493 13852
rect 8481 13821 8493 13824
rect 8527 13821 8539 13855
rect 14093 13855 14151 13861
rect 14093 13852 14105 13855
rect 8481 13815 8539 13821
rect 8588 13824 14105 13852
rect 4617 13787 4675 13793
rect 4617 13753 4629 13787
rect 4663 13753 4675 13787
rect 4617 13747 4675 13753
rect 5721 13787 5779 13793
rect 5721 13753 5733 13787
rect 5767 13784 5779 13787
rect 8202 13784 8208 13796
rect 5767 13756 8208 13784
rect 5767 13753 5779 13756
rect 5721 13747 5779 13753
rect 8202 13744 8208 13756
rect 8260 13744 8266 13796
rect 2866 13676 2872 13728
rect 2924 13716 2930 13728
rect 3418 13716 3424 13728
rect 2924 13688 3424 13716
rect 2924 13676 2930 13688
rect 3418 13676 3424 13688
rect 3476 13676 3482 13728
rect 3513 13719 3571 13725
rect 3513 13685 3525 13719
rect 3559 13716 3571 13719
rect 7558 13716 7564 13728
rect 3559 13688 7564 13716
rect 3559 13685 3571 13688
rect 3513 13679 3571 13685
rect 7558 13676 7564 13688
rect 7616 13676 7622 13728
rect 7742 13716 7748 13728
rect 7703 13688 7748 13716
rect 7742 13676 7748 13688
rect 7800 13676 7806 13728
rect 8294 13676 8300 13728
rect 8352 13716 8358 13728
rect 8588 13716 8616 13824
rect 14093 13821 14105 13824
rect 14139 13821 14151 13855
rect 14093 13815 14151 13821
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13821 14887 13855
rect 14829 13815 14887 13821
rect 8748 13787 8806 13793
rect 8748 13753 8760 13787
rect 8794 13784 8806 13787
rect 8846 13784 8852 13796
rect 8794 13756 8852 13784
rect 8794 13753 8806 13756
rect 8748 13747 8806 13753
rect 8846 13744 8852 13756
rect 8904 13744 8910 13796
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 12805 13787 12863 13793
rect 12805 13784 12817 13787
rect 9180 13756 12817 13784
rect 9180 13744 9186 13756
rect 12805 13753 12817 13756
rect 12851 13753 12863 13787
rect 13998 13784 14004 13796
rect 13959 13756 14004 13784
rect 12805 13747 12863 13753
rect 13998 13744 14004 13756
rect 14056 13744 14062 13796
rect 8352 13688 8616 13716
rect 8352 13676 8358 13688
rect 9030 13676 9036 13728
rect 9088 13716 9094 13728
rect 10689 13719 10747 13725
rect 10689 13716 10701 13719
rect 9088 13688 10701 13716
rect 9088 13676 9094 13688
rect 10689 13685 10701 13688
rect 10735 13685 10747 13719
rect 10689 13679 10747 13685
rect 10781 13719 10839 13725
rect 10781 13685 10793 13719
rect 10827 13716 10839 13719
rect 11238 13716 11244 13728
rect 10827 13688 11244 13716
rect 10827 13685 10839 13688
rect 10781 13679 10839 13685
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 11517 13719 11575 13725
rect 11517 13685 11529 13719
rect 11563 13716 11575 13719
rect 11882 13716 11888 13728
rect 11563 13688 11888 13716
rect 11563 13685 11575 13688
rect 11517 13679 11575 13685
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 12250 13676 12256 13728
rect 12308 13716 12314 13728
rect 12437 13719 12495 13725
rect 12437 13716 12449 13719
rect 12308 13688 12449 13716
rect 12308 13676 12314 13688
rect 12437 13685 12449 13688
rect 12483 13685 12495 13719
rect 12437 13679 12495 13685
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 12768 13688 13645 13716
rect 12768 13676 12774 13688
rect 13633 13685 13645 13688
rect 13679 13685 13691 13719
rect 13633 13679 13691 13685
rect 1104 13626 15824 13648
rect 1104 13574 5912 13626
rect 5964 13574 5976 13626
rect 6028 13574 6040 13626
rect 6092 13574 6104 13626
rect 6156 13574 10843 13626
rect 10895 13574 10907 13626
rect 10959 13574 10971 13626
rect 11023 13574 11035 13626
rect 11087 13574 15824 13626
rect 1104 13552 15824 13574
rect 1578 13472 1584 13524
rect 1636 13512 1642 13524
rect 5534 13512 5540 13524
rect 1636 13484 5540 13512
rect 1636 13472 1642 13484
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 8389 13515 8447 13521
rect 5776 13484 8340 13512
rect 5776 13472 5782 13484
rect 1412 13416 3096 13444
rect 1412 13385 1440 13416
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13345 1455 13379
rect 2130 13376 2136 13388
rect 2091 13348 2136 13376
rect 1397 13339 1455 13345
rect 2130 13336 2136 13348
rect 2188 13336 2194 13388
rect 2400 13379 2458 13385
rect 2400 13345 2412 13379
rect 2446 13376 2458 13379
rect 2866 13376 2872 13388
rect 2446 13348 2872 13376
rect 2446 13345 2458 13348
rect 2400 13339 2458 13345
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 3068 13376 3096 13416
rect 3142 13404 3148 13456
rect 3200 13444 3206 13456
rect 4614 13444 4620 13456
rect 3200 13416 4620 13444
rect 3200 13404 3206 13416
rect 4614 13404 4620 13416
rect 4672 13404 4678 13456
rect 5258 13453 5264 13456
rect 5252 13444 5264 13453
rect 5219 13416 5264 13444
rect 5252 13407 5264 13416
rect 5258 13404 5264 13407
rect 5316 13404 5322 13456
rect 5626 13404 5632 13456
rect 5684 13444 5690 13456
rect 8312 13444 8340 13484
rect 8389 13481 8401 13515
rect 8435 13512 8447 13515
rect 9122 13512 9128 13524
rect 8435 13484 9128 13512
rect 8435 13481 8447 13484
rect 8389 13475 8447 13481
rect 9122 13472 9128 13484
rect 9180 13472 9186 13524
rect 9490 13472 9496 13524
rect 9548 13512 9554 13524
rect 12526 13512 12532 13524
rect 9548 13484 12532 13512
rect 9548 13472 9554 13484
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 12713 13515 12771 13521
rect 12713 13481 12725 13515
rect 12759 13512 12771 13515
rect 13078 13512 13084 13524
rect 12759 13484 13084 13512
rect 12759 13481 12771 13484
rect 12713 13475 12771 13481
rect 13078 13472 13084 13484
rect 13136 13472 13142 13524
rect 14090 13472 14096 13524
rect 14148 13512 14154 13524
rect 14277 13515 14335 13521
rect 14277 13512 14289 13515
rect 14148 13484 14289 13512
rect 14148 13472 14154 13484
rect 14277 13481 14289 13484
rect 14323 13512 14335 13515
rect 14734 13512 14740 13524
rect 14323 13484 14740 13512
rect 14323 13481 14335 13484
rect 14277 13475 14335 13481
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 5684 13416 8248 13444
rect 8312 13416 8616 13444
rect 5684 13404 5690 13416
rect 7006 13376 7012 13388
rect 3068 13348 7012 13376
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 7190 13376 7196 13388
rect 7151 13348 7196 13376
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 7285 13379 7343 13385
rect 7285 13345 7297 13379
rect 7331 13376 7343 13379
rect 7742 13376 7748 13388
rect 7331 13348 7748 13376
rect 7331 13345 7343 13348
rect 7285 13339 7343 13345
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 8220 13385 8248 13416
rect 8205 13379 8263 13385
rect 8205 13345 8217 13379
rect 8251 13345 8263 13379
rect 8588 13376 8616 13416
rect 8662 13404 8668 13456
rect 8720 13444 8726 13456
rect 8757 13447 8815 13453
rect 8757 13444 8769 13447
rect 8720 13416 8769 13444
rect 8720 13404 8726 13416
rect 8757 13413 8769 13416
rect 8803 13413 8815 13447
rect 8757 13407 8815 13413
rect 8849 13447 8907 13453
rect 8849 13413 8861 13447
rect 8895 13444 8907 13447
rect 9030 13444 9036 13456
rect 8895 13416 9036 13444
rect 8895 13413 8907 13416
rect 8849 13407 8907 13413
rect 9030 13404 9036 13416
rect 9088 13404 9094 13456
rect 9674 13404 9680 13456
rect 9732 13444 9738 13456
rect 9858 13444 9864 13456
rect 9732 13416 9864 13444
rect 9732 13404 9738 13416
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 11606 13444 11612 13456
rect 9959 13416 11612 13444
rect 9959 13376 9987 13416
rect 11606 13404 11612 13416
rect 11664 13404 11670 13456
rect 13262 13404 13268 13456
rect 13320 13404 13326 13456
rect 13722 13404 13728 13456
rect 13780 13444 13786 13456
rect 14369 13447 14427 13453
rect 14369 13444 14381 13447
rect 13780 13416 14381 13444
rect 13780 13404 13786 13416
rect 14369 13413 14381 13416
rect 14415 13413 14427 13447
rect 14369 13407 14427 13413
rect 8588 13348 9987 13376
rect 8205 13339 8263 13345
rect 10502 13336 10508 13388
rect 10560 13376 10566 13388
rect 10669 13379 10727 13385
rect 10669 13376 10681 13379
rect 10560 13348 10681 13376
rect 10560 13336 10566 13348
rect 10669 13345 10681 13348
rect 10715 13345 10727 13379
rect 10669 13339 10727 13345
rect 11698 13336 11704 13388
rect 11756 13376 11762 13388
rect 12437 13379 12495 13385
rect 12437 13376 12449 13379
rect 11756 13348 12449 13376
rect 11756 13336 11762 13348
rect 12437 13345 12449 13348
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 13081 13379 13139 13385
rect 13081 13376 13093 13379
rect 12860 13348 13093 13376
rect 12860 13336 12866 13348
rect 13081 13345 13093 13348
rect 13127 13345 13139 13379
rect 13081 13339 13139 13345
rect 13173 13379 13231 13385
rect 13173 13345 13185 13379
rect 13219 13376 13231 13379
rect 13280 13376 13308 13404
rect 14826 13376 14832 13388
rect 13219 13348 14832 13376
rect 13219 13345 13231 13348
rect 13173 13339 13231 13345
rect 14826 13336 14832 13348
rect 14884 13336 14890 13388
rect 4341 13311 4399 13317
rect 4341 13277 4353 13311
rect 4387 13277 4399 13311
rect 4341 13271 4399 13277
rect 4154 13240 4160 13252
rect 3252 13212 4160 13240
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 3252 13172 3280 13212
rect 4154 13200 4160 13212
rect 4212 13200 4218 13252
rect 1627 13144 3280 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 3326 13132 3332 13184
rect 3384 13172 3390 13184
rect 3513 13175 3571 13181
rect 3513 13172 3525 13175
rect 3384 13144 3525 13172
rect 3384 13132 3390 13144
rect 3513 13141 3525 13144
rect 3559 13141 3571 13175
rect 4356 13172 4384 13271
rect 4430 13268 4436 13320
rect 4488 13308 4494 13320
rect 4985 13311 5043 13317
rect 4985 13308 4997 13311
rect 4488 13280 4997 13308
rect 4488 13268 4494 13280
rect 4985 13277 4997 13280
rect 5031 13277 5043 13311
rect 4985 13271 5043 13277
rect 7374 13268 7380 13320
rect 7432 13268 7438 13320
rect 7469 13311 7527 13317
rect 7469 13277 7481 13311
rect 7515 13308 7527 13311
rect 7926 13308 7932 13320
rect 7515 13280 7932 13308
rect 7515 13277 7527 13280
rect 7469 13271 7527 13277
rect 7392 13240 7420 13268
rect 5920 13212 7420 13240
rect 5920 13172 5948 13212
rect 4356 13144 5948 13172
rect 3513 13135 3571 13141
rect 6086 13132 6092 13184
rect 6144 13172 6150 13184
rect 6365 13175 6423 13181
rect 6365 13172 6377 13175
rect 6144 13144 6377 13172
rect 6144 13132 6150 13144
rect 6365 13141 6377 13144
rect 6411 13141 6423 13175
rect 6365 13135 6423 13141
rect 6454 13132 6460 13184
rect 6512 13172 6518 13184
rect 6825 13175 6883 13181
rect 6825 13172 6837 13175
rect 6512 13144 6837 13172
rect 6512 13132 6518 13144
rect 6825 13141 6837 13144
rect 6871 13141 6883 13175
rect 6825 13135 6883 13141
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 7484 13172 7512 13271
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 8386 13268 8392 13320
rect 8444 13308 8450 13320
rect 8846 13308 8852 13320
rect 8444 13280 8852 13308
rect 8444 13268 8450 13280
rect 8846 13268 8852 13280
rect 8904 13308 8910 13320
rect 8941 13311 8999 13317
rect 8941 13308 8953 13311
rect 8904 13280 8953 13308
rect 8904 13268 8910 13280
rect 8941 13277 8953 13280
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13277 9827 13311
rect 9769 13271 9827 13277
rect 7742 13200 7748 13252
rect 7800 13240 7806 13252
rect 7800 13212 8147 13240
rect 7800 13200 7806 13212
rect 8018 13172 8024 13184
rect 7248 13144 7512 13172
rect 7979 13144 8024 13172
rect 7248 13132 7254 13144
rect 8018 13132 8024 13144
rect 8076 13132 8082 13184
rect 8119 13172 8147 13212
rect 8202 13200 8208 13252
rect 8260 13240 8266 13252
rect 9122 13240 9128 13252
rect 8260 13212 9128 13240
rect 8260 13200 8266 13212
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 9784 13240 9812 13271
rect 9858 13268 9864 13320
rect 9916 13308 9922 13320
rect 10413 13311 10471 13317
rect 10413 13308 10425 13311
rect 9916 13280 10425 13308
rect 9916 13268 9922 13280
rect 10413 13277 10425 13280
rect 10459 13277 10471 13311
rect 10413 13271 10471 13277
rect 10226 13240 10232 13252
rect 9784 13212 10232 13240
rect 10226 13200 10232 13212
rect 10284 13200 10290 13252
rect 9858 13172 9864 13184
rect 8119 13144 9864 13172
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 10428 13172 10456 13271
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 12250 13308 12256 13320
rect 11480 13280 12256 13308
rect 11480 13268 11486 13280
rect 12250 13268 12256 13280
rect 12308 13268 12314 13320
rect 13265 13311 13323 13317
rect 13265 13277 13277 13311
rect 13311 13277 13323 13311
rect 14461 13311 14519 13317
rect 14461 13308 14473 13311
rect 13265 13271 13323 13277
rect 13372 13280 14473 13308
rect 11793 13243 11851 13249
rect 11793 13209 11805 13243
rect 11839 13240 11851 13243
rect 11974 13240 11980 13252
rect 11839 13212 11980 13240
rect 11839 13209 11851 13212
rect 11793 13203 11851 13209
rect 11974 13200 11980 13212
rect 12032 13240 12038 13252
rect 12032 13212 12848 13240
rect 12032 13200 12038 13212
rect 12253 13175 12311 13181
rect 12253 13172 12265 13175
rect 10428 13144 12265 13172
rect 12253 13141 12265 13144
rect 12299 13141 12311 13175
rect 12820 13172 12848 13212
rect 12894 13200 12900 13252
rect 12952 13240 12958 13252
rect 13280 13240 13308 13271
rect 12952 13212 13308 13240
rect 12952 13200 12958 13212
rect 13372 13172 13400 13280
rect 14461 13277 14473 13280
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 12820 13144 13400 13172
rect 13909 13175 13967 13181
rect 12253 13135 12311 13141
rect 13909 13141 13921 13175
rect 13955 13172 13967 13175
rect 13998 13172 14004 13184
rect 13955 13144 14004 13172
rect 13955 13141 13967 13144
rect 13909 13135 13967 13141
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 1104 13082 15824 13104
rect 1104 13030 3447 13082
rect 3499 13030 3511 13082
rect 3563 13030 3575 13082
rect 3627 13030 3639 13082
rect 3691 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 13308 13082
rect 13360 13030 13372 13082
rect 13424 13030 13436 13082
rect 13488 13030 13500 13082
rect 13552 13030 15824 13082
rect 1104 13008 15824 13030
rect 3145 12971 3203 12977
rect 3145 12937 3157 12971
rect 3191 12968 3203 12971
rect 5350 12968 5356 12980
rect 3191 12940 5356 12968
rect 3191 12937 3203 12940
rect 3145 12931 3203 12937
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 5442 12928 5448 12980
rect 5500 12968 5506 12980
rect 5500 12940 6868 12968
rect 5500 12928 5506 12940
rect 2130 12860 2136 12912
rect 2188 12900 2194 12912
rect 2314 12900 2320 12912
rect 2188 12872 2320 12900
rect 2188 12860 2194 12872
rect 2314 12860 2320 12872
rect 2372 12860 2378 12912
rect 4798 12860 4804 12912
rect 4856 12900 4862 12912
rect 5258 12900 5264 12912
rect 4856 12872 5264 12900
rect 4856 12860 4862 12872
rect 5258 12860 5264 12872
rect 5316 12860 5322 12912
rect 5537 12903 5595 12909
rect 5537 12869 5549 12903
rect 5583 12900 5595 12903
rect 6730 12900 6736 12912
rect 5583 12872 6736 12900
rect 5583 12869 5595 12872
rect 5537 12863 5595 12869
rect 6730 12860 6736 12872
rect 6788 12860 6794 12912
rect 6840 12900 6868 12940
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 7834 12968 7840 12980
rect 7064 12940 7840 12968
rect 7064 12928 7070 12940
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 7926 12928 7932 12980
rect 7984 12968 7990 12980
rect 8754 12968 8760 12980
rect 7984 12940 8760 12968
rect 7984 12928 7990 12940
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 8941 12971 8999 12977
rect 8941 12937 8953 12971
rect 8987 12968 8999 12971
rect 9030 12968 9036 12980
rect 8987 12940 9036 12968
rect 8987 12937 8999 12940
rect 8941 12931 8999 12937
rect 9030 12928 9036 12940
rect 9088 12928 9094 12980
rect 9950 12928 9956 12980
rect 10008 12968 10014 12980
rect 10008 12940 11468 12968
rect 10008 12928 10014 12940
rect 10781 12903 10839 12909
rect 10781 12900 10793 12903
rect 6840 12872 10793 12900
rect 10781 12869 10793 12872
rect 10827 12869 10839 12903
rect 10781 12863 10839 12869
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12832 2651 12835
rect 3602 12832 3608 12844
rect 2639 12804 3608 12832
rect 2639 12801 2651 12804
rect 2593 12795 2651 12801
rect 3602 12792 3608 12804
rect 3660 12792 3666 12844
rect 3786 12832 3792 12844
rect 3747 12804 3792 12832
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 4430 12792 4436 12844
rect 4488 12832 4494 12844
rect 4614 12832 4620 12844
rect 4488 12804 4620 12832
rect 4488 12792 4494 12804
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12832 5043 12835
rect 5074 12832 5080 12844
rect 5031 12804 5080 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 5902 12792 5908 12844
rect 5960 12832 5966 12844
rect 5997 12835 6055 12841
rect 5997 12832 6009 12835
rect 5960 12804 6009 12832
rect 5960 12792 5966 12804
rect 5997 12801 6009 12804
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6086 12792 6092 12844
rect 6144 12832 6150 12844
rect 7926 12832 7932 12844
rect 6144 12804 6189 12832
rect 6748 12804 7932 12832
rect 6144 12792 6150 12804
rect 2317 12767 2375 12773
rect 2317 12733 2329 12767
rect 2363 12764 2375 12767
rect 2406 12764 2412 12776
rect 2363 12736 2412 12764
rect 2363 12733 2375 12736
rect 2317 12727 2375 12733
rect 2406 12724 2412 12736
rect 2464 12764 2470 12776
rect 2682 12764 2688 12776
rect 2464 12736 2688 12764
rect 2464 12724 2470 12736
rect 2682 12724 2688 12736
rect 2740 12724 2746 12776
rect 3513 12767 3571 12773
rect 3513 12733 3525 12767
rect 3559 12764 3571 12767
rect 6748 12764 6776 12804
rect 7926 12792 7932 12804
rect 7984 12792 7990 12844
rect 8386 12841 8392 12844
rect 8343 12835 8392 12841
rect 8343 12801 8355 12835
rect 8389 12801 8392 12835
rect 8343 12795 8392 12801
rect 8386 12792 8392 12795
rect 8444 12792 8450 12844
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 9306 12832 9312 12844
rect 8904 12804 9312 12832
rect 8904 12792 8910 12804
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 10042 12832 10048 12844
rect 9631 12804 10048 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 11330 12832 11336 12844
rect 11291 12804 11336 12832
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 11440 12832 11468 12940
rect 11606 12928 11612 12980
rect 11664 12968 11670 12980
rect 13633 12971 13691 12977
rect 13633 12968 13645 12971
rect 11664 12940 13645 12968
rect 11664 12928 11670 12940
rect 13633 12937 13645 12940
rect 13679 12937 13691 12971
rect 13633 12931 13691 12937
rect 11514 12860 11520 12912
rect 11572 12900 11578 12912
rect 12437 12903 12495 12909
rect 12437 12900 12449 12903
rect 11572 12872 12449 12900
rect 11572 12860 11578 12872
rect 12437 12869 12449 12872
rect 12483 12869 12495 12903
rect 12437 12863 12495 12869
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 15013 12903 15071 12909
rect 15013 12900 15025 12903
rect 12584 12872 15025 12900
rect 12584 12860 12590 12872
rect 15013 12869 15025 12872
rect 15059 12869 15071 12903
rect 15013 12863 15071 12869
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 11440 12804 13001 12832
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 14182 12832 14188 12844
rect 14143 12804 14188 12832
rect 12989 12795 13047 12801
rect 14182 12792 14188 12804
rect 14240 12792 14246 12844
rect 3559 12736 6776 12764
rect 6825 12767 6883 12773
rect 3559 12733 3571 12736
rect 3513 12727 3571 12733
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 6825 12727 6883 12733
rect 3605 12699 3663 12705
rect 3605 12696 3617 12699
rect 1964 12668 3617 12696
rect 1964 12637 1992 12668
rect 3605 12665 3617 12668
rect 3651 12665 3663 12699
rect 3605 12659 3663 12665
rect 3786 12656 3792 12708
rect 3844 12696 3850 12708
rect 3970 12696 3976 12708
rect 3844 12668 3976 12696
rect 3844 12656 3850 12668
rect 3970 12656 3976 12668
rect 4028 12656 4034 12708
rect 4154 12656 4160 12708
rect 4212 12696 4218 12708
rect 4801 12699 4859 12705
rect 4801 12696 4813 12699
rect 4212 12668 4813 12696
rect 4212 12656 4218 12668
rect 4801 12665 4813 12668
rect 4847 12665 4859 12699
rect 4801 12659 4859 12665
rect 5442 12656 5448 12708
rect 5500 12696 5506 12708
rect 6840 12696 6868 12727
rect 7282 12724 7288 12776
rect 7340 12764 7346 12776
rect 8110 12764 8116 12776
rect 7340 12736 8116 12764
rect 7340 12724 7346 12736
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 8812 12736 9628 12764
rect 8812 12724 8818 12736
rect 5500 12668 6868 12696
rect 5500 12656 5506 12668
rect 7006 12656 7012 12708
rect 7064 12696 7070 12708
rect 7101 12699 7159 12705
rect 7101 12696 7113 12699
rect 7064 12668 7113 12696
rect 7064 12656 7070 12668
rect 7101 12665 7113 12668
rect 7147 12665 7159 12699
rect 7101 12659 7159 12665
rect 7558 12656 7564 12708
rect 7616 12696 7622 12708
rect 9030 12696 9036 12708
rect 7616 12668 9036 12696
rect 7616 12656 7622 12668
rect 9030 12656 9036 12668
rect 9088 12656 9094 12708
rect 9309 12699 9367 12705
rect 9309 12665 9321 12699
rect 9355 12696 9367 12699
rect 9490 12696 9496 12708
rect 9355 12668 9496 12696
rect 9355 12665 9367 12668
rect 9309 12659 9367 12665
rect 9490 12656 9496 12668
rect 9548 12656 9554 12708
rect 9600 12696 9628 12736
rect 10502 12724 10508 12776
rect 10560 12764 10566 12776
rect 11149 12767 11207 12773
rect 11149 12764 11161 12767
rect 10560 12736 11161 12764
rect 10560 12724 10566 12736
rect 11149 12733 11161 12736
rect 11195 12733 11207 12767
rect 11149 12727 11207 12733
rect 11238 12724 11244 12776
rect 11296 12764 11302 12776
rect 12526 12764 12532 12776
rect 11296 12736 12532 12764
rect 11296 12724 11302 12736
rect 12526 12724 12532 12736
rect 12584 12724 12590 12776
rect 12897 12767 12955 12773
rect 12897 12733 12909 12767
rect 12943 12764 12955 12767
rect 13906 12764 13912 12776
rect 12943 12736 13912 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 13906 12724 13912 12736
rect 13964 12724 13970 12776
rect 14826 12764 14832 12776
rect 14739 12736 14832 12764
rect 14826 12724 14832 12736
rect 14884 12764 14890 12776
rect 15102 12764 15108 12776
rect 14884 12736 15108 12764
rect 14884 12724 14890 12736
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 11514 12696 11520 12708
rect 9600 12668 11520 12696
rect 11514 12656 11520 12668
rect 11572 12656 11578 12708
rect 13630 12656 13636 12708
rect 13688 12696 13694 12708
rect 14093 12699 14151 12705
rect 14093 12696 14105 12699
rect 13688 12668 14105 12696
rect 13688 12656 13694 12668
rect 14093 12665 14105 12668
rect 14139 12665 14151 12699
rect 14093 12659 14151 12665
rect 1949 12631 2007 12637
rect 1949 12597 1961 12631
rect 1995 12597 2007 12631
rect 2406 12628 2412 12640
rect 2319 12600 2412 12628
rect 1949 12591 2007 12597
rect 2406 12588 2412 12600
rect 2464 12628 2470 12640
rect 3050 12628 3056 12640
rect 2464 12600 3056 12628
rect 2464 12588 2470 12600
rect 3050 12588 3056 12600
rect 3108 12588 3114 12640
rect 4338 12628 4344 12640
rect 4299 12600 4344 12628
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 4430 12588 4436 12640
rect 4488 12628 4494 12640
rect 4709 12631 4767 12637
rect 4709 12628 4721 12631
rect 4488 12600 4721 12628
rect 4488 12588 4494 12600
rect 4709 12597 4721 12600
rect 4755 12597 4767 12631
rect 4709 12591 4767 12597
rect 5810 12588 5816 12640
rect 5868 12628 5874 12640
rect 5905 12631 5963 12637
rect 5905 12628 5917 12631
rect 5868 12600 5917 12628
rect 5868 12588 5874 12600
rect 5905 12597 5917 12600
rect 5951 12597 5963 12631
rect 7742 12628 7748 12640
rect 7703 12600 7748 12628
rect 5905 12591 5963 12597
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 7926 12588 7932 12640
rect 7984 12628 7990 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 7984 12600 8217 12628
rect 7984 12588 7990 12600
rect 8205 12597 8217 12600
rect 8251 12597 8263 12631
rect 8205 12591 8263 12597
rect 8938 12588 8944 12640
rect 8996 12628 9002 12640
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 8996 12600 9413 12628
rect 8996 12588 9002 12600
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 9401 12591 9459 12597
rect 10042 12588 10048 12640
rect 10100 12628 10106 12640
rect 10137 12631 10195 12637
rect 10137 12628 10149 12631
rect 10100 12600 10149 12628
rect 10100 12588 10106 12600
rect 10137 12597 10149 12600
rect 10183 12597 10195 12631
rect 10137 12591 10195 12597
rect 10410 12588 10416 12640
rect 10468 12628 10474 12640
rect 11241 12631 11299 12637
rect 11241 12628 11253 12631
rect 10468 12600 11253 12628
rect 10468 12588 10474 12600
rect 11241 12597 11253 12600
rect 11287 12628 11299 12631
rect 12158 12628 12164 12640
rect 11287 12600 12164 12628
rect 11287 12597 11299 12600
rect 11241 12591 11299 12597
rect 12158 12588 12164 12600
rect 12216 12628 12222 12640
rect 12805 12631 12863 12637
rect 12805 12628 12817 12631
rect 12216 12600 12817 12628
rect 12216 12588 12222 12600
rect 12805 12597 12817 12600
rect 12851 12597 12863 12631
rect 12805 12591 12863 12597
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14001 12631 14059 12637
rect 14001 12628 14013 12631
rect 13964 12600 14013 12628
rect 13964 12588 13970 12600
rect 14001 12597 14013 12600
rect 14047 12597 14059 12631
rect 14001 12591 14059 12597
rect 1104 12538 15824 12560
rect 1104 12486 5912 12538
rect 5964 12486 5976 12538
rect 6028 12486 6040 12538
rect 6092 12486 6104 12538
rect 6156 12486 10843 12538
rect 10895 12486 10907 12538
rect 10959 12486 10971 12538
rect 11023 12486 11035 12538
rect 11087 12486 15824 12538
rect 1104 12464 15824 12486
rect 1949 12427 2007 12433
rect 1949 12393 1961 12427
rect 1995 12424 2007 12427
rect 2038 12424 2044 12436
rect 1995 12396 2044 12424
rect 1995 12393 2007 12396
rect 1949 12387 2007 12393
rect 2038 12384 2044 12396
rect 2096 12384 2102 12436
rect 3142 12424 3148 12436
rect 3103 12396 3148 12424
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 3234 12384 3240 12436
rect 3292 12424 3298 12436
rect 7466 12424 7472 12436
rect 3292 12396 3337 12424
rect 6831 12396 7472 12424
rect 3292 12384 3298 12396
rect 4065 12359 4123 12365
rect 4065 12325 4077 12359
rect 4111 12356 4123 12359
rect 6638 12356 6644 12368
rect 4111 12328 5948 12356
rect 4111 12325 4123 12328
rect 4065 12319 4123 12325
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12288 2099 12291
rect 2774 12288 2780 12300
rect 2087 12260 2780 12288
rect 2087 12257 2099 12260
rect 2041 12251 2099 12257
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 3050 12248 3056 12300
rect 3108 12288 3114 12300
rect 4430 12288 4436 12300
rect 3108 12260 4436 12288
rect 3108 12248 3114 12260
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 4706 12288 4712 12300
rect 4667 12260 4712 12288
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 4976 12291 5034 12297
rect 4976 12257 4988 12291
rect 5022 12288 5034 12291
rect 5258 12288 5264 12300
rect 5022 12260 5264 12288
rect 5022 12257 5034 12260
rect 4976 12251 5034 12257
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 5920 12288 5948 12328
rect 6104 12328 6644 12356
rect 6104 12288 6132 12328
rect 6638 12316 6644 12328
rect 6696 12316 6702 12368
rect 6831 12365 6859 12396
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 7558 12384 7564 12436
rect 7616 12424 7622 12436
rect 7929 12427 7987 12433
rect 7929 12424 7941 12427
rect 7616 12396 7941 12424
rect 7616 12384 7622 12396
rect 7929 12393 7941 12396
rect 7975 12393 7987 12427
rect 7929 12387 7987 12393
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 11057 12427 11115 12433
rect 11057 12424 11069 12427
rect 8076 12396 11069 12424
rect 8076 12384 8082 12396
rect 6816 12359 6874 12365
rect 6816 12325 6828 12359
rect 6862 12325 6874 12359
rect 6816 12319 6874 12325
rect 6914 12316 6920 12368
rect 6972 12356 6978 12368
rect 8757 12359 8815 12365
rect 8757 12356 8769 12359
rect 6972 12328 8769 12356
rect 6972 12316 6978 12328
rect 8757 12325 8769 12328
rect 8803 12325 8815 12359
rect 8757 12319 8815 12325
rect 8386 12288 8392 12300
rect 5920 12260 6132 12288
rect 6187 12260 8392 12288
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12220 2283 12223
rect 3421 12223 3479 12229
rect 3421 12220 3433 12223
rect 2271 12192 3433 12220
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 3421 12189 3433 12192
rect 3467 12220 3479 12223
rect 3467 12192 4752 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 4724 12164 4752 12192
rect 5994 12180 6000 12232
rect 6052 12220 6058 12232
rect 6187 12220 6215 12260
rect 8386 12248 8392 12260
rect 8444 12248 8450 12300
rect 6556 12223 6614 12229
rect 6556 12220 6568 12223
rect 6052 12192 6215 12220
rect 6052 12180 6058 12192
rect 6544 12189 6568 12220
rect 6602 12189 6614 12223
rect 6544 12183 6614 12189
rect 1581 12155 1639 12161
rect 1581 12121 1593 12155
rect 1627 12152 1639 12155
rect 3050 12152 3056 12164
rect 1627 12124 3056 12152
rect 1627 12121 1639 12124
rect 1581 12115 1639 12121
rect 3050 12112 3056 12124
rect 3108 12112 3114 12164
rect 3234 12112 3240 12164
rect 3292 12152 3298 12164
rect 4338 12152 4344 12164
rect 3292 12124 4344 12152
rect 3292 12112 3298 12124
rect 4338 12112 4344 12124
rect 4396 12112 4402 12164
rect 4706 12112 4712 12164
rect 4764 12112 4770 12164
rect 5718 12112 5724 12164
rect 5776 12152 5782 12164
rect 6178 12152 6184 12164
rect 5776 12124 6184 12152
rect 5776 12112 5782 12124
rect 6178 12112 6184 12124
rect 6236 12112 6242 12164
rect 2777 12087 2835 12093
rect 2777 12053 2789 12087
rect 2823 12084 2835 12087
rect 4154 12084 4160 12096
rect 2823 12056 4160 12084
rect 2823 12053 2835 12056
rect 2777 12047 2835 12053
rect 4154 12044 4160 12056
rect 4212 12044 4218 12096
rect 4614 12044 4620 12096
rect 4672 12084 4678 12096
rect 5442 12084 5448 12096
rect 4672 12056 5448 12084
rect 4672 12044 4678 12056
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 6086 12084 6092 12096
rect 6047 12056 6092 12084
rect 6086 12044 6092 12056
rect 6144 12044 6150 12096
rect 6544 12084 6572 12183
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 8754 12220 8760 12232
rect 7616 12192 8760 12220
rect 7616 12180 7622 12192
rect 8754 12180 8760 12192
rect 8812 12180 8818 12232
rect 9048 12229 9076 12396
rect 11057 12393 11069 12396
rect 11103 12424 11115 12427
rect 11330 12424 11336 12436
rect 11103 12396 11336 12424
rect 11103 12393 11115 12396
rect 11057 12387 11115 12393
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 11422 12384 11428 12436
rect 11480 12424 11486 12436
rect 12069 12427 12127 12433
rect 12069 12424 12081 12427
rect 11480 12396 12081 12424
rect 11480 12384 11486 12396
rect 12069 12393 12081 12396
rect 12115 12393 12127 12427
rect 12434 12424 12440 12436
rect 12395 12396 12440 12424
rect 12069 12387 12127 12393
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 14642 12356 14648 12368
rect 9140 12328 14648 12356
rect 8849 12223 8907 12229
rect 8849 12189 8861 12223
rect 8895 12189 8907 12223
rect 8849 12183 8907 12189
rect 9033 12223 9091 12229
rect 9033 12189 9045 12223
rect 9079 12189 9091 12223
rect 9033 12183 9091 12189
rect 8386 12152 8392 12164
rect 8347 12124 8392 12152
rect 8386 12112 8392 12124
rect 8444 12112 8450 12164
rect 8662 12112 8668 12164
rect 8720 12152 8726 12164
rect 8864 12152 8892 12183
rect 9140 12152 9168 12328
rect 14642 12316 14648 12328
rect 14700 12316 14706 12368
rect 9766 12288 9772 12300
rect 8720 12124 9168 12152
rect 9232 12260 9772 12288
rect 8720 12112 8726 12124
rect 7282 12084 7288 12096
rect 6544 12056 7288 12084
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 8846 12044 8852 12096
rect 8904 12084 8910 12096
rect 9232 12084 9260 12260
rect 9766 12248 9772 12260
rect 9824 12288 9830 12300
rect 9933 12291 9991 12297
rect 9933 12288 9945 12291
rect 9824 12260 9945 12288
rect 9824 12248 9830 12260
rect 9933 12257 9945 12260
rect 9979 12257 9991 12291
rect 9933 12251 9991 12257
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12257 11759 12291
rect 11701 12251 11759 12257
rect 9674 12220 9680 12232
rect 9635 12192 9680 12220
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 11020 12192 11560 12220
rect 11020 12180 11026 12192
rect 11238 12152 11244 12164
rect 10796 12124 11244 12152
rect 8904 12056 9260 12084
rect 8904 12044 8910 12056
rect 9306 12044 9312 12096
rect 9364 12084 9370 12096
rect 9674 12084 9680 12096
rect 9364 12056 9680 12084
rect 9364 12044 9370 12056
rect 9674 12044 9680 12056
rect 9732 12044 9738 12096
rect 10686 12044 10692 12096
rect 10744 12084 10750 12096
rect 10796 12084 10824 12124
rect 11238 12112 11244 12124
rect 11296 12112 11302 12164
rect 11532 12161 11560 12192
rect 11606 12180 11612 12232
rect 11664 12220 11670 12232
rect 11716 12220 11744 12251
rect 12250 12248 12256 12300
rect 12308 12288 12314 12300
rect 13262 12288 13268 12300
rect 12308 12260 12664 12288
rect 13223 12260 13268 12288
rect 12308 12248 12314 12260
rect 12526 12220 12532 12232
rect 11664 12192 11744 12220
rect 12487 12192 12532 12220
rect 11664 12180 11670 12192
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 12636 12229 12664 12260
rect 13262 12248 13268 12260
rect 13320 12248 13326 12300
rect 14182 12288 14188 12300
rect 14143 12260 14188 12288
rect 14182 12248 14188 12260
rect 14240 12248 14246 12300
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 13446 12220 13452 12232
rect 13407 12192 13452 12220
rect 12621 12183 12679 12189
rect 13446 12180 13452 12192
rect 13504 12180 13510 12232
rect 13538 12180 13544 12232
rect 13596 12220 13602 12232
rect 14369 12223 14427 12229
rect 14369 12220 14381 12223
rect 13596 12192 14381 12220
rect 13596 12180 13602 12192
rect 14369 12189 14381 12192
rect 14415 12189 14427 12223
rect 14369 12183 14427 12189
rect 11517 12155 11575 12161
rect 11517 12121 11529 12155
rect 11563 12121 11575 12155
rect 11517 12115 11575 12121
rect 10744 12056 10824 12084
rect 10744 12044 10750 12056
rect 10870 12044 10876 12096
rect 10928 12084 10934 12096
rect 12066 12084 12072 12096
rect 10928 12056 12072 12084
rect 10928 12044 10934 12056
rect 12066 12044 12072 12056
rect 12124 12084 12130 12096
rect 13078 12084 13084 12096
rect 12124 12056 13084 12084
rect 12124 12044 12130 12056
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 1104 11994 15824 12016
rect 1104 11942 3447 11994
rect 3499 11942 3511 11994
rect 3563 11942 3575 11994
rect 3627 11942 3639 11994
rect 3691 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 13308 11994
rect 13360 11942 13372 11994
rect 13424 11942 13436 11994
rect 13488 11942 13500 11994
rect 13552 11942 15824 11994
rect 1104 11920 15824 11942
rect 1854 11880 1860 11892
rect 1815 11852 1860 11880
rect 1854 11840 1860 11852
rect 1912 11840 1918 11892
rect 2038 11840 2044 11892
rect 2096 11880 2102 11892
rect 5994 11880 6000 11892
rect 2096 11852 6000 11880
rect 2096 11840 2102 11852
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 6086 11840 6092 11892
rect 6144 11880 6150 11892
rect 8938 11880 8944 11892
rect 6144 11852 8944 11880
rect 6144 11840 6150 11852
rect 8938 11840 8944 11852
rect 8996 11840 9002 11892
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 10318 11880 10324 11892
rect 9272 11852 10324 11880
rect 9272 11840 9278 11852
rect 10318 11840 10324 11852
rect 10376 11840 10382 11892
rect 11606 11840 11612 11892
rect 11664 11880 11670 11892
rect 11885 11883 11943 11889
rect 11885 11880 11897 11883
rect 11664 11852 11897 11880
rect 11664 11840 11670 11852
rect 11885 11849 11897 11852
rect 11931 11849 11943 11883
rect 11885 11843 11943 11849
rect 2314 11772 2320 11824
rect 2372 11812 2378 11824
rect 2372 11784 3096 11812
rect 2372 11772 2378 11784
rect 3068 11753 3096 11784
rect 6178 11772 6184 11824
rect 6236 11812 6242 11824
rect 6273 11815 6331 11821
rect 6273 11812 6285 11815
rect 6236 11784 6285 11812
rect 6236 11772 6242 11784
rect 6273 11781 6285 11784
rect 6319 11812 6331 11815
rect 6822 11812 6828 11824
rect 6319 11784 6828 11812
rect 6319 11781 6331 11784
rect 6273 11775 6331 11781
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 8205 11815 8263 11821
rect 8205 11781 8217 11815
rect 8251 11812 8263 11815
rect 10870 11812 10876 11824
rect 8251 11784 10876 11812
rect 8251 11781 8263 11784
rect 8205 11775 8263 11781
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11744 2559 11747
rect 3053 11747 3111 11753
rect 2547 11716 3004 11744
rect 2547 11713 2559 11716
rect 2501 11707 2559 11713
rect 2222 11676 2228 11688
rect 2135 11648 2228 11676
rect 2222 11636 2228 11648
rect 2280 11676 2286 11688
rect 2682 11676 2688 11688
rect 2280 11648 2688 11676
rect 2280 11636 2286 11648
rect 2682 11636 2688 11648
rect 2740 11636 2746 11688
rect 2976 11676 3004 11716
rect 3053 11713 3065 11747
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 4724 11716 5028 11744
rect 4724 11676 4752 11716
rect 4890 11676 4896 11688
rect 2976 11648 4752 11676
rect 4851 11648 4896 11676
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 5000 11676 5028 11716
rect 5902 11704 5908 11756
rect 5960 11744 5966 11756
rect 6638 11744 6644 11756
rect 5960 11716 6644 11744
rect 5960 11704 5966 11716
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 6748 11716 6960 11744
rect 6270 11676 6276 11688
rect 5000 11648 6276 11676
rect 6270 11636 6276 11648
rect 6328 11676 6334 11688
rect 6748 11676 6776 11716
rect 6328 11648 6776 11676
rect 6825 11679 6883 11685
rect 6328 11636 6334 11648
rect 6825 11645 6837 11679
rect 6871 11645 6883 11679
rect 6932 11676 6960 11716
rect 7081 11679 7139 11685
rect 7081 11676 7093 11679
rect 6932 11648 7093 11676
rect 6825 11639 6883 11645
rect 7081 11645 7093 11648
rect 7127 11645 7139 11679
rect 7081 11639 7139 11645
rect 2317 11611 2375 11617
rect 2317 11577 2329 11611
rect 2363 11608 2375 11611
rect 2406 11608 2412 11620
rect 2363 11580 2412 11608
rect 2363 11577 2375 11580
rect 2317 11571 2375 11577
rect 2406 11568 2412 11580
rect 2464 11608 2470 11620
rect 3142 11608 3148 11620
rect 2464 11580 3148 11608
rect 2464 11568 2470 11580
rect 3142 11568 3148 11580
rect 3200 11568 3206 11620
rect 3320 11611 3378 11617
rect 3320 11577 3332 11611
rect 3366 11577 3378 11611
rect 3320 11571 3378 11577
rect 3344 11540 3372 11571
rect 3418 11568 3424 11620
rect 3476 11608 3482 11620
rect 5138 11611 5196 11617
rect 5138 11608 5150 11611
rect 3476 11580 5150 11608
rect 3476 11568 3482 11580
rect 5138 11577 5150 11580
rect 5184 11577 5196 11611
rect 5138 11571 5196 11577
rect 5258 11568 5264 11620
rect 5316 11608 5322 11620
rect 6730 11608 6736 11620
rect 5316 11580 6736 11608
rect 5316 11568 5322 11580
rect 6730 11568 6736 11580
rect 6788 11568 6794 11620
rect 6840 11608 6868 11639
rect 7466 11636 7472 11688
rect 7524 11676 7530 11688
rect 8220 11676 8248 11775
rect 10870 11772 10876 11784
rect 10928 11772 10934 11824
rect 11146 11772 11152 11824
rect 11204 11812 11210 11824
rect 11514 11812 11520 11824
rect 11204 11784 11520 11812
rect 11204 11772 11210 11784
rect 11514 11772 11520 11784
rect 11572 11772 11578 11824
rect 13814 11812 13820 11824
rect 11624 11784 13820 11812
rect 11624 11756 11652 11784
rect 13814 11772 13820 11784
rect 13872 11772 13878 11824
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8536 11716 8984 11744
rect 8536 11704 8542 11716
rect 8662 11676 8668 11688
rect 7524 11648 8248 11676
rect 8623 11648 8668 11676
rect 7524 11636 7530 11648
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 8846 11636 8852 11688
rect 8904 11636 8910 11688
rect 6914 11608 6920 11620
rect 6840 11580 6920 11608
rect 6914 11568 6920 11580
rect 6972 11568 6978 11620
rect 8864 11608 8892 11636
rect 8119 11580 8892 11608
rect 8956 11608 8984 11716
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 9953 11747 10011 11753
rect 9953 11744 9965 11747
rect 9364 11716 9965 11744
rect 9364 11704 9370 11716
rect 9953 11713 9965 11716
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11744 10655 11747
rect 11054 11744 11060 11756
rect 10643 11716 11060 11744
rect 10643 11713 10655 11716
rect 10597 11707 10655 11713
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 11241 11747 11299 11753
rect 11241 11744 11253 11747
rect 11164 11716 11253 11744
rect 11164 11688 11192 11716
rect 11241 11713 11253 11716
rect 11287 11713 11299 11747
rect 11241 11707 11299 11713
rect 11606 11704 11612 11756
rect 11664 11704 11670 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12176 11716 13001 11744
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 9861 11679 9919 11685
rect 9861 11676 9873 11679
rect 9732 11648 9873 11676
rect 9732 11636 9738 11648
rect 9861 11645 9873 11648
rect 9907 11645 9919 11679
rect 10962 11676 10968 11688
rect 9861 11639 9919 11645
rect 9948 11648 10968 11676
rect 9948 11608 9976 11648
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11146 11636 11152 11688
rect 11204 11636 11210 11688
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11256 11648 12081 11676
rect 8956 11580 9976 11608
rect 3786 11540 3792 11552
rect 3344 11512 3792 11540
rect 3786 11500 3792 11512
rect 3844 11500 3850 11552
rect 4433 11543 4491 11549
rect 4433 11509 4445 11543
rect 4479 11540 4491 11543
rect 8119 11540 8147 11580
rect 10318 11568 10324 11620
rect 10376 11608 10382 11620
rect 11256 11608 11284 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 10376 11580 11284 11608
rect 10376 11568 10382 11580
rect 11330 11568 11336 11620
rect 11388 11608 11394 11620
rect 12176 11608 12204 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 13170 11636 13176 11688
rect 13228 11676 13234 11688
rect 13633 11679 13691 11685
rect 13633 11676 13645 11679
rect 13228 11648 13645 11676
rect 13228 11636 13234 11648
rect 13633 11645 13645 11648
rect 13679 11645 13691 11679
rect 13633 11639 13691 11645
rect 14369 11679 14427 11685
rect 14369 11645 14381 11679
rect 14415 11676 14427 11679
rect 14458 11676 14464 11688
rect 14415 11648 14464 11676
rect 14415 11645 14427 11648
rect 14369 11639 14427 11645
rect 14458 11636 14464 11648
rect 14516 11676 14522 11688
rect 15930 11676 15936 11688
rect 14516 11648 15936 11676
rect 14516 11636 14522 11648
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 12526 11608 12532 11620
rect 11388 11580 12204 11608
rect 12268 11580 12532 11608
rect 11388 11568 11394 11580
rect 4479 11512 8147 11540
rect 4479 11509 4491 11512
rect 4433 11503 4491 11509
rect 8202 11500 8208 11552
rect 8260 11540 8266 11552
rect 8849 11543 8907 11549
rect 8849 11540 8861 11543
rect 8260 11512 8861 11540
rect 8260 11500 8266 11512
rect 8849 11509 8861 11512
rect 8895 11509 8907 11543
rect 8849 11503 8907 11509
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 9401 11543 9459 11549
rect 9401 11540 9413 11543
rect 8996 11512 9413 11540
rect 8996 11500 9002 11512
rect 9401 11509 9413 11512
rect 9447 11509 9459 11543
rect 9401 11503 9459 11509
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 9769 11543 9827 11549
rect 9769 11540 9781 11543
rect 9732 11512 9781 11540
rect 9732 11500 9738 11512
rect 9769 11509 9781 11512
rect 9815 11509 9827 11543
rect 9769 11503 9827 11509
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 12268 11540 12296 11580
rect 12526 11568 12532 11580
rect 12584 11568 12590 11620
rect 12710 11568 12716 11620
rect 12768 11608 12774 11620
rect 12805 11611 12863 11617
rect 12805 11608 12817 11611
rect 12768 11580 12817 11608
rect 12768 11568 12774 11580
rect 12805 11577 12817 11580
rect 12851 11577 12863 11611
rect 12805 11571 12863 11577
rect 13262 11568 13268 11620
rect 13320 11608 13326 11620
rect 13320 11580 14596 11608
rect 13320 11568 13326 11580
rect 10008 11512 12296 11540
rect 10008 11500 10014 11512
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12894 11540 12900 11552
rect 12492 11512 12537 11540
rect 12855 11512 12900 11540
rect 12492 11500 12498 11512
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 13538 11500 13544 11552
rect 13596 11540 13602 11552
rect 14568 11549 14596 11580
rect 13817 11543 13875 11549
rect 13817 11540 13829 11543
rect 13596 11512 13829 11540
rect 13596 11500 13602 11512
rect 13817 11509 13829 11512
rect 13863 11509 13875 11543
rect 13817 11503 13875 11509
rect 14553 11543 14611 11549
rect 14553 11509 14565 11543
rect 14599 11509 14611 11543
rect 14553 11503 14611 11509
rect 1104 11450 15824 11472
rect 1104 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 6104 11450
rect 6156 11398 10843 11450
rect 10895 11398 10907 11450
rect 10959 11398 10971 11450
rect 11023 11398 11035 11450
rect 11087 11398 15824 11450
rect 1104 11376 15824 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2682 11336 2688 11348
rect 1995 11308 2688 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 2823 11308 2912 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 2038 11268 2044 11280
rect 1999 11240 2044 11268
rect 2038 11228 2044 11240
rect 2096 11228 2102 11280
rect 2884 11268 2912 11308
rect 3050 11296 3056 11348
rect 3108 11336 3114 11348
rect 4062 11336 4068 11348
rect 3108 11308 4068 11336
rect 3108 11296 3114 11308
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4338 11336 4344 11348
rect 4299 11308 4344 11336
rect 4338 11296 4344 11308
rect 4396 11296 4402 11348
rect 4801 11339 4859 11345
rect 4801 11305 4813 11339
rect 4847 11336 4859 11339
rect 6546 11336 6552 11348
rect 4847 11308 6552 11336
rect 4847 11305 4859 11308
rect 4801 11299 4859 11305
rect 6546 11296 6552 11308
rect 6604 11296 6610 11348
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 6917 11339 6975 11345
rect 6917 11336 6929 11339
rect 6788 11308 6929 11336
rect 6788 11296 6794 11308
rect 6917 11305 6929 11308
rect 6963 11305 6975 11339
rect 6917 11299 6975 11305
rect 7024 11308 7788 11336
rect 3145 11271 3203 11277
rect 2884 11240 3096 11268
rect 3068 11200 3096 11240
rect 3145 11237 3157 11271
rect 3191 11268 3203 11271
rect 7024 11268 7052 11308
rect 7650 11277 7656 11280
rect 3191 11240 7052 11268
rect 7622 11271 7656 11277
rect 3191 11237 3203 11240
rect 3145 11231 3203 11237
rect 7622 11237 7634 11271
rect 7622 11231 7656 11237
rect 7650 11228 7656 11231
rect 7708 11228 7714 11280
rect 7760 11268 7788 11308
rect 8110 11296 8116 11348
rect 8168 11336 8174 11348
rect 9214 11336 9220 11348
rect 8168 11308 8791 11336
rect 9175 11308 9220 11336
rect 8168 11296 8174 11308
rect 8570 11268 8576 11280
rect 7760 11240 8576 11268
rect 8570 11228 8576 11240
rect 8628 11228 8634 11280
rect 8763 11268 8791 11308
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 9674 11336 9680 11348
rect 9635 11308 9680 11336
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 11333 11339 11391 11345
rect 11333 11305 11345 11339
rect 11379 11336 11391 11339
rect 11606 11336 11612 11348
rect 11379 11308 11612 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 12069 11339 12127 11345
rect 12069 11305 12081 11339
rect 12115 11336 12127 11339
rect 12710 11336 12716 11348
rect 12115 11308 12716 11336
rect 12115 11305 12127 11308
rect 12069 11299 12127 11305
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 13630 11296 13636 11348
rect 13688 11336 13694 11348
rect 13725 11339 13783 11345
rect 13725 11336 13737 11339
rect 13688 11308 13737 11336
rect 13688 11296 13694 11308
rect 13725 11305 13737 11308
rect 13771 11305 13783 11339
rect 13725 11299 13783 11305
rect 9306 11268 9312 11280
rect 8763 11240 9312 11268
rect 9306 11228 9312 11240
rect 9364 11228 9370 11280
rect 10042 11268 10048 11280
rect 10003 11240 10048 11268
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 11514 11228 11520 11280
rect 11572 11268 11578 11280
rect 12437 11271 12495 11277
rect 12437 11268 12449 11271
rect 11572 11240 12449 11268
rect 11572 11228 11578 11240
rect 12437 11237 12449 11240
rect 12483 11237 12495 11271
rect 12437 11231 12495 11237
rect 12529 11271 12587 11277
rect 12529 11237 12541 11271
rect 12575 11268 12587 11271
rect 14274 11268 14280 11280
rect 12575 11240 14280 11268
rect 12575 11237 12587 11240
rect 12529 11231 12587 11237
rect 14274 11228 14280 11240
rect 14332 11228 14338 11280
rect 3068 11172 4016 11200
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 3050 11132 3056 11144
rect 2271 11104 3056 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 3234 11132 3240 11144
rect 3195 11104 3240 11132
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 3326 11092 3332 11144
rect 3384 11132 3390 11144
rect 3988 11132 4016 11172
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4709 11203 4767 11209
rect 4709 11200 4721 11203
rect 4212 11172 4721 11200
rect 4212 11160 4218 11172
rect 4709 11169 4721 11172
rect 4755 11169 4767 11203
rect 5442 11200 5448 11212
rect 4709 11163 4767 11169
rect 4816 11172 5448 11200
rect 4816 11132 4844 11172
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 5804 11203 5862 11209
rect 5804 11169 5816 11203
rect 5850 11200 5862 11203
rect 6546 11200 6552 11212
rect 5850 11172 6552 11200
rect 5850 11169 5862 11172
rect 5804 11163 5862 11169
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 7377 11203 7435 11209
rect 7377 11200 7389 11203
rect 6972 11172 7389 11200
rect 6972 11160 6978 11172
rect 7377 11169 7389 11172
rect 7423 11200 7435 11203
rect 8478 11200 8484 11212
rect 7423 11172 8484 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 9401 11203 9459 11209
rect 9401 11200 9413 11203
rect 8680 11172 9413 11200
rect 8680 11144 8708 11172
rect 9401 11169 9413 11172
rect 9447 11169 9459 11203
rect 9401 11163 9459 11169
rect 9493 11203 9551 11209
rect 9493 11169 9505 11203
rect 9539 11200 9551 11203
rect 9858 11200 9864 11212
rect 9539 11172 9864 11200
rect 9539 11169 9551 11172
rect 9493 11163 9551 11169
rect 9858 11160 9864 11172
rect 9916 11160 9922 11212
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11200 10195 11203
rect 11241 11203 11299 11209
rect 10183 11172 11192 11200
rect 10183 11169 10195 11172
rect 10137 11163 10195 11169
rect 4982 11132 4988 11144
rect 3384 11104 3429 11132
rect 3988 11104 4844 11132
rect 4943 11104 4988 11132
rect 3384 11092 3390 11104
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5350 11092 5356 11144
rect 5408 11132 5414 11144
rect 5537 11135 5595 11141
rect 5537 11132 5549 11135
rect 5408 11104 5549 11132
rect 5408 11092 5414 11104
rect 5537 11101 5549 11104
rect 5583 11101 5595 11135
rect 5537 11095 5595 11101
rect 8662 11092 8668 11144
rect 8720 11092 8726 11144
rect 10229 11135 10287 11141
rect 10229 11132 10241 11135
rect 8772 11104 10241 11132
rect 1670 11024 1676 11076
rect 1728 11064 1734 11076
rect 5074 11064 5080 11076
rect 1728 11036 5080 11064
rect 1728 11024 1734 11036
rect 5074 11024 5080 11036
rect 5132 11024 5138 11076
rect 6546 11024 6552 11076
rect 6604 11064 6610 11076
rect 7098 11064 7104 11076
rect 6604 11036 7104 11064
rect 6604 11024 6610 11036
rect 7098 11024 7104 11036
rect 7156 11024 7162 11076
rect 8386 11024 8392 11076
rect 8444 11064 8450 11076
rect 8772 11073 8800 11104
rect 10229 11101 10241 11104
rect 10275 11101 10287 11135
rect 11164 11132 11192 11172
rect 11241 11169 11253 11203
rect 11287 11200 11299 11203
rect 11330 11200 11336 11212
rect 11287 11172 11336 11200
rect 11287 11169 11299 11172
rect 11241 11163 11299 11169
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 12250 11200 12256 11212
rect 11532 11172 12256 11200
rect 11532 11141 11560 11172
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 12802 11160 12808 11212
rect 12860 11200 12866 11212
rect 13262 11200 13268 11212
rect 12860 11172 13268 11200
rect 12860 11160 12866 11172
rect 13262 11160 13268 11172
rect 13320 11160 13326 11212
rect 13630 11200 13636 11212
rect 13591 11172 13636 11200
rect 13630 11160 13636 11172
rect 13688 11200 13694 11212
rect 13906 11200 13912 11212
rect 13688 11172 13912 11200
rect 13688 11160 13694 11172
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11200 14519 11203
rect 15470 11200 15476 11212
rect 14507 11172 15476 11200
rect 14507 11169 14519 11172
rect 14461 11163 14519 11169
rect 11517 11135 11575 11141
rect 11164 11104 11284 11132
rect 10229 11095 10287 11101
rect 11256 11076 11284 11104
rect 11517 11101 11529 11135
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 12342 11132 12348 11144
rect 12032 11104 12348 11132
rect 12032 11092 12038 11104
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12618 11132 12624 11144
rect 12579 11104 12624 11132
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 13817 11135 13875 11141
rect 13817 11132 13829 11135
rect 12728 11104 13829 11132
rect 8757 11067 8815 11073
rect 8757 11064 8769 11067
rect 8444 11036 8769 11064
rect 8444 11024 8450 11036
rect 8757 11033 8769 11036
rect 8803 11033 8815 11067
rect 9493 11067 9551 11073
rect 9493 11064 9505 11067
rect 8757 11027 8815 11033
rect 9048 11036 9505 11064
rect 3050 10956 3056 11008
rect 3108 10996 3114 11008
rect 4890 10996 4896 11008
rect 3108 10968 4896 10996
rect 3108 10956 3114 10968
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 5718 10956 5724 11008
rect 5776 10996 5782 11008
rect 6730 10996 6736 11008
rect 5776 10968 6736 10996
rect 5776 10956 5782 10968
rect 6730 10956 6736 10968
rect 6788 10956 6794 11008
rect 6822 10956 6828 11008
rect 6880 10996 6886 11008
rect 9048 10996 9076 11036
rect 9493 11033 9505 11036
rect 9539 11033 9551 11067
rect 9493 11027 9551 11033
rect 9766 11024 9772 11076
rect 9824 11064 9830 11076
rect 10873 11067 10931 11073
rect 10873 11064 10885 11067
rect 9824 11036 10885 11064
rect 9824 11024 9830 11036
rect 10873 11033 10885 11036
rect 10919 11033 10931 11067
rect 10873 11027 10931 11033
rect 11238 11024 11244 11076
rect 11296 11024 11302 11076
rect 6880 10968 9076 10996
rect 6880 10956 6886 10968
rect 9214 10956 9220 11008
rect 9272 10996 9278 11008
rect 12728 10996 12756 11104
rect 13817 11101 13829 11104
rect 13863 11101 13875 11135
rect 13817 11095 13875 11101
rect 13262 11064 13268 11076
rect 13223 11036 13268 11064
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 13906 11024 13912 11076
rect 13964 11064 13970 11076
rect 14476 11064 14504 11163
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 13964 11036 14504 11064
rect 13964 11024 13970 11036
rect 9272 10968 12756 10996
rect 9272 10956 9278 10968
rect 13078 10956 13084 11008
rect 13136 10996 13142 11008
rect 14645 10999 14703 11005
rect 14645 10996 14657 10999
rect 13136 10968 14657 10996
rect 13136 10956 13142 10968
rect 14645 10965 14657 10968
rect 14691 10965 14703 10999
rect 14645 10959 14703 10965
rect 1104 10906 15824 10928
rect 1104 10854 3447 10906
rect 3499 10854 3511 10906
rect 3563 10854 3575 10906
rect 3627 10854 3639 10906
rect 3691 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 13308 10906
rect 13360 10854 13372 10906
rect 13424 10854 13436 10906
rect 13488 10854 13500 10906
rect 13552 10854 15824 10906
rect 1104 10832 15824 10854
rect 2682 10752 2688 10804
rect 2740 10752 2746 10804
rect 3786 10792 3792 10804
rect 2976 10764 3792 10792
rect 2700 10724 2728 10752
rect 1964 10696 2728 10724
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10588 1823 10591
rect 1964 10588 1992 10696
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10625 2099 10659
rect 2682 10656 2688 10668
rect 2643 10628 2688 10656
rect 2041 10619 2099 10625
rect 1811 10560 1992 10588
rect 2056 10588 2084 10619
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 2866 10656 2872 10668
rect 2827 10628 2872 10656
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 2976 10588 3004 10764
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 4632 10764 5856 10792
rect 3050 10616 3056 10668
rect 3108 10656 3114 10668
rect 3108 10628 3153 10656
rect 3108 10616 3114 10628
rect 3602 10588 3608 10600
rect 2056 10560 3004 10588
rect 3252 10560 3608 10588
rect 1811 10557 1823 10560
rect 1765 10551 1823 10557
rect 2406 10520 2412 10532
rect 1412 10492 2412 10520
rect 1412 10461 1440 10492
rect 2406 10480 2412 10492
rect 2464 10480 2470 10532
rect 2593 10523 2651 10529
rect 2593 10489 2605 10523
rect 2639 10520 2651 10523
rect 3252 10520 3280 10560
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 2639 10492 3280 10520
rect 3320 10523 3378 10529
rect 2639 10489 2651 10492
rect 2593 10483 2651 10489
rect 3320 10489 3332 10523
rect 3366 10520 3378 10523
rect 4632 10520 4660 10764
rect 5828 10724 5856 10764
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 6273 10795 6331 10801
rect 6273 10792 6285 10795
rect 5960 10764 6285 10792
rect 5960 10752 5966 10764
rect 6273 10761 6285 10764
rect 6319 10761 6331 10795
rect 6273 10755 6331 10761
rect 6454 10752 6460 10804
rect 6512 10792 6518 10804
rect 7558 10792 7564 10804
rect 6512 10764 7564 10792
rect 6512 10752 6518 10764
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 8018 10752 8024 10804
rect 8076 10792 8082 10804
rect 8665 10795 8723 10801
rect 8665 10792 8677 10795
rect 8076 10764 8677 10792
rect 8076 10752 8082 10764
rect 8665 10761 8677 10764
rect 8711 10761 8723 10795
rect 8665 10755 8723 10761
rect 9861 10795 9919 10801
rect 9861 10761 9873 10795
rect 9907 10792 9919 10795
rect 9950 10792 9956 10804
rect 9907 10764 9956 10792
rect 9907 10761 9919 10764
rect 9861 10755 9919 10761
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 10226 10752 10232 10804
rect 10284 10792 10290 10804
rect 10686 10792 10692 10804
rect 10284 10764 10692 10792
rect 10284 10752 10290 10764
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 12437 10795 12495 10801
rect 12437 10792 12449 10795
rect 10796 10764 12449 10792
rect 5828 10696 6776 10724
rect 4890 10656 4896 10668
rect 4851 10628 4896 10656
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5718 10548 5724 10600
rect 5776 10588 5782 10600
rect 6454 10588 6460 10600
rect 5776 10560 6460 10588
rect 5776 10548 5782 10560
rect 6454 10548 6460 10560
rect 6512 10548 6518 10600
rect 3366 10492 4660 10520
rect 3366 10489 3378 10492
rect 3320 10483 3378 10489
rect 4706 10480 4712 10532
rect 4764 10520 4770 10532
rect 5160 10523 5218 10529
rect 5160 10520 5172 10523
rect 4764 10492 5172 10520
rect 4764 10480 4770 10492
rect 5160 10489 5172 10492
rect 5206 10520 5218 10523
rect 6748 10520 6776 10696
rect 9140 10696 9628 10724
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 9140 10665 9168 10696
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 8168 10628 9137 10656
rect 8168 10616 8174 10628
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10588 6883 10591
rect 6914 10588 6920 10600
rect 6871 10560 6920 10588
rect 6871 10557 6883 10560
rect 6825 10551 6883 10557
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 7098 10597 7104 10600
rect 7092 10588 7104 10597
rect 7059 10560 7104 10588
rect 7092 10551 7104 10560
rect 7098 10548 7104 10551
rect 7156 10548 7162 10600
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 9232 10588 9260 10619
rect 7708 10560 9260 10588
rect 9600 10588 9628 10696
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 10796 10724 10824 10764
rect 12437 10761 12449 10764
rect 12483 10761 12495 10795
rect 12437 10755 12495 10761
rect 12986 10752 12992 10804
rect 13044 10792 13050 10804
rect 13044 10764 13124 10792
rect 13044 10752 13050 10764
rect 9732 10696 10824 10724
rect 9732 10684 9738 10696
rect 11146 10684 11152 10736
rect 11204 10724 11210 10736
rect 12066 10724 12072 10736
rect 11204 10696 12072 10724
rect 11204 10684 11210 10696
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 10505 10659 10563 10665
rect 10505 10656 10517 10659
rect 9916 10628 10517 10656
rect 9916 10616 9922 10628
rect 10505 10625 10517 10628
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 10778 10616 10784 10668
rect 10836 10656 10842 10668
rect 11514 10656 11520 10668
rect 10836 10628 11520 10656
rect 10836 10616 10842 10628
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 11624 10665 11652 10696
rect 12066 10684 12072 10696
rect 12124 10684 12130 10736
rect 11609 10659 11667 10665
rect 11609 10625 11621 10659
rect 11655 10625 11667 10659
rect 11609 10619 11667 10625
rect 12618 10616 12624 10668
rect 12676 10656 12682 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12676 10628 13001 10656
rect 12676 10616 12682 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 9600 10560 10088 10588
rect 7708 10548 7714 10560
rect 7834 10520 7840 10532
rect 5206 10492 6408 10520
rect 6748 10492 7840 10520
rect 5206 10489 5218 10492
rect 5160 10483 5218 10489
rect 1397 10455 1455 10461
rect 1397 10421 1409 10455
rect 1443 10421 1455 10455
rect 1397 10415 1455 10421
rect 1857 10455 1915 10461
rect 1857 10421 1869 10455
rect 1903 10452 1915 10455
rect 2225 10455 2283 10461
rect 2225 10452 2237 10455
rect 1903 10424 2237 10452
rect 1903 10421 1915 10424
rect 1857 10415 1915 10421
rect 2225 10421 2237 10424
rect 2271 10421 2283 10455
rect 2225 10415 2283 10421
rect 3050 10412 3056 10464
rect 3108 10452 3114 10464
rect 4433 10455 4491 10461
rect 4433 10452 4445 10455
rect 3108 10424 4445 10452
rect 3108 10412 3114 10424
rect 4433 10421 4445 10424
rect 4479 10452 4491 10455
rect 6270 10452 6276 10464
rect 4479 10424 6276 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 6380 10452 6408 10492
rect 7834 10480 7840 10492
rect 7892 10480 7898 10532
rect 8018 10480 8024 10532
rect 8076 10520 8082 10532
rect 8662 10520 8668 10532
rect 8076 10492 8668 10520
rect 8076 10480 8082 10492
rect 8662 10480 8668 10492
rect 8720 10480 8726 10532
rect 9033 10523 9091 10529
rect 9033 10489 9045 10523
rect 9079 10520 9091 10523
rect 9674 10520 9680 10532
rect 9079 10492 9680 10520
rect 9079 10489 9091 10492
rect 9033 10483 9091 10489
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 10060 10520 10088 10560
rect 10134 10548 10140 10600
rect 10192 10588 10198 10600
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 10192 10560 10241 10588
rect 10192 10548 10198 10560
rect 10229 10557 10241 10560
rect 10275 10557 10287 10591
rect 10229 10551 10287 10557
rect 10321 10591 10379 10597
rect 10321 10557 10333 10591
rect 10367 10588 10379 10591
rect 10410 10588 10416 10600
rect 10367 10560 10416 10588
rect 10367 10557 10379 10560
rect 10321 10551 10379 10557
rect 10410 10548 10416 10560
rect 10468 10548 10474 10600
rect 11425 10591 11483 10597
rect 10704 10560 10916 10588
rect 10704 10520 10732 10560
rect 10060 10492 10732 10520
rect 10778 10480 10784 10532
rect 10836 10480 10842 10532
rect 10888 10520 10916 10560
rect 11425 10557 11437 10591
rect 11471 10588 11483 10591
rect 13096 10588 13124 10764
rect 14734 10656 14740 10668
rect 14695 10628 14740 10656
rect 14734 10616 14740 10628
rect 14792 10616 14798 10668
rect 13262 10588 13268 10600
rect 11471 10560 13268 10588
rect 11471 10557 11483 10560
rect 11425 10551 11483 10557
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 13633 10591 13691 10597
rect 13633 10557 13645 10591
rect 13679 10557 13691 10591
rect 13633 10551 13691 10557
rect 12066 10520 12072 10532
rect 10888 10492 12072 10520
rect 12066 10480 12072 10492
rect 12124 10520 12130 10532
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 12124 10492 12817 10520
rect 12124 10480 12130 10492
rect 12805 10489 12817 10492
rect 12851 10489 12863 10523
rect 12805 10483 12863 10489
rect 12986 10480 12992 10532
rect 13044 10520 13050 10532
rect 13648 10520 13676 10551
rect 13722 10548 13728 10600
rect 13780 10588 13786 10600
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 13780 10560 14565 10588
rect 13780 10548 13786 10560
rect 14553 10557 14565 10560
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 13906 10520 13912 10532
rect 13044 10492 13676 10520
rect 13867 10492 13912 10520
rect 13044 10480 13050 10492
rect 13906 10480 13912 10492
rect 13964 10480 13970 10532
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 6380 10424 8217 10452
rect 8205 10421 8217 10424
rect 8251 10421 8263 10455
rect 8205 10415 8263 10421
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 10796 10452 10824 10480
rect 8352 10424 10824 10452
rect 11057 10455 11115 10461
rect 8352 10412 8358 10424
rect 11057 10421 11069 10455
rect 11103 10452 11115 10455
rect 11422 10452 11428 10464
rect 11103 10424 11428 10452
rect 11103 10421 11115 10424
rect 11057 10415 11115 10421
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 11517 10455 11575 10461
rect 11517 10421 11529 10455
rect 11563 10452 11575 10455
rect 11974 10452 11980 10464
rect 11563 10424 11980 10452
rect 11563 10421 11575 10424
rect 11517 10415 11575 10421
rect 11974 10412 11980 10424
rect 12032 10452 12038 10464
rect 12250 10452 12256 10464
rect 12032 10424 12256 10452
rect 12032 10412 12038 10424
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 12342 10412 12348 10464
rect 12400 10452 12406 10464
rect 12897 10455 12955 10461
rect 12897 10452 12909 10455
rect 12400 10424 12909 10452
rect 12400 10412 12406 10424
rect 12897 10421 12909 10424
rect 12943 10452 12955 10455
rect 15194 10452 15200 10464
rect 12943 10424 15200 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 1104 10362 15824 10384
rect 1104 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 6104 10362
rect 6156 10310 10843 10362
rect 10895 10310 10907 10362
rect 10959 10310 10971 10362
rect 11023 10310 11035 10362
rect 11087 10310 15824 10362
rect 1104 10288 15824 10310
rect 1489 10251 1547 10257
rect 1489 10217 1501 10251
rect 1535 10248 1547 10251
rect 2682 10248 2688 10260
rect 1535 10220 2688 10248
rect 1535 10217 1547 10220
rect 1489 10211 1547 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 7101 10251 7159 10257
rect 2823 10220 6224 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 1857 10183 1915 10189
rect 1857 10149 1869 10183
rect 1903 10180 1915 10183
rect 4522 10180 4528 10192
rect 1903 10152 4528 10180
rect 1903 10149 1915 10152
rect 1857 10143 1915 10149
rect 4522 10140 4528 10152
rect 4580 10180 4586 10192
rect 4893 10183 4951 10189
rect 4893 10180 4905 10183
rect 4580 10152 4905 10180
rect 4580 10140 4586 10152
rect 4893 10149 4905 10152
rect 4939 10180 4951 10183
rect 5718 10180 5724 10192
rect 4939 10152 5724 10180
rect 4939 10149 4951 10152
rect 4893 10143 4951 10149
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 5810 10140 5816 10192
rect 5868 10180 5874 10192
rect 5966 10183 6024 10189
rect 5966 10180 5978 10183
rect 5868 10152 5978 10180
rect 5868 10140 5874 10152
rect 5966 10149 5978 10152
rect 6012 10149 6024 10183
rect 5966 10143 6024 10149
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 2774 10112 2780 10124
rect 2731 10084 2780 10112
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 3050 10112 3056 10124
rect 2976 10084 3056 10112
rect 1854 10004 1860 10056
rect 1912 10044 1918 10056
rect 2976 10053 3004 10084
rect 3050 10072 3056 10084
rect 3108 10072 3114 10124
rect 3418 10072 3424 10124
rect 3476 10112 3482 10124
rect 3513 10115 3571 10121
rect 3513 10112 3525 10115
rect 3476 10084 3525 10112
rect 3476 10072 3482 10084
rect 3513 10081 3525 10084
rect 3559 10081 3571 10115
rect 5534 10112 5540 10124
rect 3513 10075 3571 10081
rect 3712 10084 5540 10112
rect 1949 10047 2007 10053
rect 1949 10044 1961 10047
rect 1912 10016 1961 10044
rect 1912 10004 1918 10016
rect 1949 10013 1961 10016
rect 1995 10013 2007 10047
rect 1949 10007 2007 10013
rect 2133 10047 2191 10053
rect 2133 10013 2145 10047
rect 2179 10013 2191 10047
rect 2133 10007 2191 10013
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 2148 9976 2176 10007
rect 3142 10004 3148 10056
rect 3200 10044 3206 10056
rect 3605 10047 3663 10053
rect 3605 10044 3617 10047
rect 3200 10016 3617 10044
rect 3200 10004 3206 10016
rect 3605 10013 3617 10016
rect 3651 10013 3663 10047
rect 3605 10007 3663 10013
rect 3712 9976 3740 10084
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 6196 10112 6224 10220
rect 7101 10217 7113 10251
rect 7147 10248 7159 10251
rect 7190 10248 7196 10260
rect 7147 10220 7196 10248
rect 7147 10217 7159 10220
rect 7101 10211 7159 10217
rect 7190 10208 7196 10220
rect 7248 10248 7254 10260
rect 7650 10248 7656 10260
rect 7248 10220 7656 10248
rect 7248 10208 7254 10220
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 7926 10208 7932 10260
rect 7984 10248 7990 10260
rect 8386 10248 8392 10260
rect 7984 10220 8392 10248
rect 7984 10208 7990 10220
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 8662 10208 8668 10260
rect 8720 10248 8726 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8720 10220 8953 10248
rect 8720 10208 8726 10220
rect 8941 10217 8953 10220
rect 8987 10248 8999 10251
rect 9214 10248 9220 10260
rect 8987 10220 9220 10248
rect 8987 10217 8999 10220
rect 8941 10211 8999 10217
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 9324 10220 10456 10248
rect 6270 10140 6276 10192
rect 6328 10180 6334 10192
rect 7806 10183 7864 10189
rect 7806 10180 7818 10183
rect 6328 10152 7818 10180
rect 6328 10140 6334 10152
rect 7806 10149 7818 10152
rect 7852 10149 7864 10183
rect 9324 10180 9352 10220
rect 7806 10143 7864 10149
rect 7935 10152 9352 10180
rect 7935 10112 7963 10152
rect 9766 10140 9772 10192
rect 9824 10180 9830 10192
rect 10137 10183 10195 10189
rect 10137 10180 10149 10183
rect 9824 10152 10149 10180
rect 9824 10140 9830 10152
rect 10137 10149 10149 10152
rect 10183 10180 10195 10183
rect 10318 10180 10324 10192
rect 10183 10152 10324 10180
rect 10183 10149 10195 10152
rect 10137 10143 10195 10149
rect 10318 10140 10324 10152
rect 10376 10140 10382 10192
rect 10428 10180 10456 10220
rect 10502 10208 10508 10260
rect 10560 10248 10566 10260
rect 11333 10251 11391 10257
rect 11333 10248 11345 10251
rect 10560 10220 11345 10248
rect 10560 10208 10566 10220
rect 11333 10217 11345 10220
rect 11379 10248 11391 10251
rect 11974 10248 11980 10260
rect 11379 10220 11980 10248
rect 11379 10217 11391 10220
rect 11333 10211 11391 10217
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12069 10251 12127 10257
rect 12069 10217 12081 10251
rect 12115 10217 12127 10251
rect 12069 10211 12127 10217
rect 12437 10251 12495 10257
rect 12437 10217 12449 10251
rect 12483 10248 12495 10251
rect 13265 10251 13323 10257
rect 13265 10248 13277 10251
rect 12483 10220 13277 10248
rect 12483 10217 12495 10220
rect 12437 10211 12495 10217
rect 13265 10217 13277 10220
rect 13311 10217 13323 10251
rect 13265 10211 13323 10217
rect 12084 10180 12112 10211
rect 10428 10152 12112 10180
rect 12618 10140 12624 10192
rect 12676 10140 12682 10192
rect 12802 10140 12808 10192
rect 12860 10180 12866 10192
rect 12860 10152 13032 10180
rect 12860 10140 12866 10152
rect 6196 10084 7963 10112
rect 8110 10072 8116 10124
rect 8168 10112 8174 10124
rect 8294 10112 8300 10124
rect 8168 10084 8300 10112
rect 8168 10072 8174 10084
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 10042 10112 10048 10124
rect 8444 10084 10048 10112
rect 8444 10072 8450 10084
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 10502 10112 10508 10124
rect 10152 10084 10508 10112
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 2148 9948 3740 9976
rect 2314 9908 2320 9920
rect 2275 9880 2320 9908
rect 2314 9868 2320 9880
rect 2372 9868 2378 9920
rect 2406 9868 2412 9920
rect 2464 9908 2470 9920
rect 2958 9908 2964 9920
rect 2464 9880 2964 9908
rect 2464 9868 2470 9880
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 3142 9908 3148 9920
rect 3103 9880 3148 9908
rect 3142 9868 3148 9880
rect 3200 9868 3206 9920
rect 3804 9908 3832 10007
rect 4430 10004 4436 10056
rect 4488 10044 4494 10056
rect 4985 10047 5043 10053
rect 4985 10044 4997 10047
rect 4488 10016 4997 10044
rect 4488 10004 4494 10016
rect 4985 10013 4997 10016
rect 5031 10013 5043 10047
rect 5166 10044 5172 10056
rect 5127 10016 5172 10044
rect 4985 10007 5043 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 5442 10004 5448 10056
rect 5500 10044 5506 10056
rect 5721 10047 5779 10053
rect 5721 10044 5733 10047
rect 5500 10016 5733 10044
rect 5500 10004 5506 10016
rect 5721 10013 5733 10016
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 6914 10004 6920 10056
rect 6972 10044 6978 10056
rect 7558 10044 7564 10056
rect 6972 10016 7564 10044
rect 6972 10004 6978 10016
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 10152 10044 10180 10084
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 10744 10084 11253 10112
rect 10744 10072 10750 10084
rect 11241 10081 11253 10084
rect 11287 10081 11299 10115
rect 12636 10112 12664 10140
rect 11241 10075 11299 10081
rect 11532 10084 12664 10112
rect 9732 10016 10180 10044
rect 10321 10047 10379 10053
rect 9732 10004 9738 10016
rect 10321 10013 10333 10047
rect 10367 10044 10379 10047
rect 11146 10044 11152 10056
rect 10367 10016 11152 10044
rect 10367 10013 10379 10016
rect 10321 10007 10379 10013
rect 11146 10004 11152 10016
rect 11204 10004 11210 10056
rect 11422 10004 11428 10056
rect 11480 10044 11486 10056
rect 11532 10053 11560 10084
rect 12894 10072 12900 10124
rect 12952 10072 12958 10124
rect 13004 10112 13032 10152
rect 13170 10140 13176 10192
rect 13228 10180 13234 10192
rect 13633 10183 13691 10189
rect 13633 10180 13645 10183
rect 13228 10152 13645 10180
rect 13228 10140 13234 10152
rect 13633 10149 13645 10152
rect 13679 10149 13691 10183
rect 13633 10143 13691 10149
rect 13538 10112 13544 10124
rect 13004 10084 13544 10112
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 14274 10072 14280 10124
rect 14332 10112 14338 10124
rect 14461 10115 14519 10121
rect 14461 10112 14473 10115
rect 14332 10084 14473 10112
rect 14332 10072 14338 10084
rect 14461 10081 14473 10084
rect 14507 10112 14519 10115
rect 14734 10112 14740 10124
rect 14507 10084 14740 10112
rect 14507 10081 14519 10084
rect 14461 10075 14519 10081
rect 14734 10072 14740 10084
rect 14792 10072 14798 10124
rect 11517 10047 11575 10053
rect 11517 10044 11529 10047
rect 11480 10016 11529 10044
rect 11480 10004 11486 10016
rect 11517 10013 11529 10016
rect 11563 10013 11575 10047
rect 12526 10044 12532 10056
rect 12487 10016 12532 10044
rect 11517 10007 11575 10013
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 12676 10016 12721 10044
rect 12676 10004 12682 10016
rect 4525 9979 4583 9985
rect 4525 9945 4537 9979
rect 4571 9976 4583 9979
rect 5626 9976 5632 9988
rect 4571 9948 5632 9976
rect 4571 9945 4583 9948
rect 4525 9939 4583 9945
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 8938 9936 8944 9988
rect 8996 9976 9002 9988
rect 10594 9976 10600 9988
rect 8996 9948 10600 9976
rect 8996 9936 9002 9948
rect 10594 9936 10600 9948
rect 10652 9936 10658 9988
rect 10873 9979 10931 9985
rect 10873 9945 10885 9979
rect 10919 9976 10931 9979
rect 12912 9976 12940 10072
rect 13722 10044 13728 10056
rect 13683 10016 13728 10044
rect 13722 10004 13728 10016
rect 13780 10004 13786 10056
rect 13817 10047 13875 10053
rect 13817 10013 13829 10047
rect 13863 10013 13875 10047
rect 13817 10007 13875 10013
rect 10919 9948 12940 9976
rect 10919 9945 10931 9948
rect 10873 9939 10931 9945
rect 13078 9936 13084 9988
rect 13136 9976 13142 9988
rect 13832 9976 13860 10007
rect 14642 9976 14648 9988
rect 13136 9948 13860 9976
rect 14603 9948 14648 9976
rect 13136 9936 13142 9948
rect 14642 9936 14648 9948
rect 14700 9936 14706 9988
rect 6086 9908 6092 9920
rect 3804 9880 6092 9908
rect 6086 9868 6092 9880
rect 6144 9868 6150 9920
rect 6730 9868 6736 9920
rect 6788 9908 6794 9920
rect 9677 9911 9735 9917
rect 9677 9908 9689 9911
rect 6788 9880 9689 9908
rect 6788 9868 6794 9880
rect 9677 9877 9689 9880
rect 9723 9877 9735 9911
rect 9677 9871 9735 9877
rect 10042 9868 10048 9920
rect 10100 9908 10106 9920
rect 12894 9908 12900 9920
rect 10100 9880 12900 9908
rect 10100 9868 10106 9880
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 1104 9818 15824 9840
rect 1104 9766 3447 9818
rect 3499 9766 3511 9818
rect 3563 9766 3575 9818
rect 3627 9766 3639 9818
rect 3691 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 13308 9818
rect 13360 9766 13372 9818
rect 13424 9766 13436 9818
rect 13488 9766 13500 9818
rect 13552 9766 15824 9818
rect 1104 9744 15824 9766
rect 1486 9664 1492 9716
rect 1544 9704 1550 9716
rect 3050 9704 3056 9716
rect 1544 9676 3056 9704
rect 1544 9664 1550 9676
rect 3050 9664 3056 9676
rect 3108 9664 3114 9716
rect 5442 9704 5448 9716
rect 3804 9676 5448 9704
rect 2777 9639 2835 9645
rect 2777 9605 2789 9639
rect 2823 9636 2835 9639
rect 3602 9636 3608 9648
rect 2823 9608 3608 9636
rect 2823 9605 2835 9608
rect 2777 9599 2835 9605
rect 3602 9596 3608 9608
rect 3660 9596 3666 9648
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 3421 9571 3479 9577
rect 2271 9540 3372 9568
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 2041 9503 2099 9509
rect 2041 9469 2053 9503
rect 2087 9500 2099 9503
rect 3142 9500 3148 9512
rect 2087 9472 3148 9500
rect 2087 9469 2099 9472
rect 2041 9463 2099 9469
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 1946 9432 1952 9444
rect 1907 9404 1952 9432
rect 1946 9392 1952 9404
rect 2004 9392 2010 9444
rect 2682 9392 2688 9444
rect 2740 9432 2746 9444
rect 3237 9435 3295 9441
rect 3237 9432 3249 9435
rect 2740 9404 3249 9432
rect 2740 9392 2746 9404
rect 3237 9401 3249 9404
rect 3283 9401 3295 9435
rect 3344 9432 3372 9540
rect 3421 9537 3433 9571
rect 3467 9568 3479 9571
rect 3694 9568 3700 9580
rect 3467 9540 3700 9568
rect 3467 9537 3479 9540
rect 3421 9531 3479 9537
rect 3694 9528 3700 9540
rect 3752 9528 3758 9580
rect 3804 9577 3832 9676
rect 5276 9577 5304 9676
rect 5442 9664 5448 9676
rect 5500 9664 5506 9716
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 5592 9676 8217 9704
rect 5592 9664 5598 9676
rect 8205 9673 8217 9676
rect 8251 9704 8263 9707
rect 11422 9704 11428 9716
rect 8251 9676 11428 9704
rect 8251 9673 8263 9676
rect 8205 9667 8263 9673
rect 11422 9664 11428 9676
rect 11480 9664 11486 9716
rect 14642 9704 14648 9716
rect 13648 9676 14648 9704
rect 13648 9648 13676 9676
rect 14642 9664 14648 9676
rect 14700 9664 14706 9716
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6641 9639 6699 9645
rect 6641 9636 6653 9639
rect 6604 9608 6653 9636
rect 6604 9596 6610 9608
rect 6641 9605 6653 9608
rect 6687 9605 6699 9639
rect 6641 9599 6699 9605
rect 7926 9596 7932 9648
rect 7984 9636 7990 9648
rect 8294 9636 8300 9648
rect 7984 9608 8300 9636
rect 7984 9596 7990 9608
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 8570 9596 8576 9648
rect 8628 9636 8634 9648
rect 9674 9636 9680 9648
rect 8628 9608 9680 9636
rect 8628 9596 8634 9608
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 9861 9639 9919 9645
rect 9861 9605 9873 9639
rect 9907 9636 9919 9639
rect 11146 9636 11152 9648
rect 9907 9608 11152 9636
rect 9907 9605 9919 9608
rect 9861 9599 9919 9605
rect 11146 9596 11152 9608
rect 11204 9596 11210 9648
rect 12802 9636 12808 9648
rect 11256 9608 12808 9636
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 9217 9571 9275 9577
rect 9217 9568 9229 9571
rect 7892 9540 9229 9568
rect 7892 9528 7898 9540
rect 9217 9537 9229 9540
rect 9263 9537 9275 9571
rect 9217 9531 9275 9537
rect 10226 9528 10232 9580
rect 10284 9568 10290 9580
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 10284 9540 10425 9568
rect 10284 9528 10290 9540
rect 10413 9537 10425 9540
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10594 9528 10600 9580
rect 10652 9568 10658 9580
rect 11256 9568 11284 9608
rect 12802 9596 12808 9608
rect 12860 9596 12866 9648
rect 13630 9636 13636 9648
rect 12912 9608 13636 9636
rect 10652 9540 11284 9568
rect 11609 9571 11667 9577
rect 10652 9528 10658 9540
rect 11609 9537 11621 9571
rect 11655 9568 11667 9571
rect 12618 9568 12624 9580
rect 11655 9540 12624 9568
rect 11655 9537 11667 9540
rect 11609 9531 11667 9537
rect 4053 9509 4059 9512
rect 4045 9503 4059 9509
rect 4045 9469 4057 9503
rect 4111 9500 4117 9512
rect 4111 9472 4145 9500
rect 4045 9463 4059 9469
rect 4053 9460 4059 9463
rect 4111 9460 4117 9472
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 6825 9503 6883 9509
rect 5132 9472 5764 9500
rect 5132 9460 5138 9472
rect 5534 9441 5540 9444
rect 3344 9404 5488 9432
rect 3237 9395 3295 9401
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 3142 9364 3148 9376
rect 3103 9336 3148 9364
rect 3142 9324 3148 9336
rect 3200 9324 3206 9376
rect 3786 9324 3792 9376
rect 3844 9364 3850 9376
rect 5169 9367 5227 9373
rect 5169 9364 5181 9367
rect 3844 9336 5181 9364
rect 3844 9324 3850 9336
rect 5169 9333 5181 9336
rect 5215 9333 5227 9367
rect 5460 9364 5488 9404
rect 5528 9395 5540 9441
rect 5592 9432 5598 9444
rect 5736 9432 5764 9472
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 6914 9500 6920 9512
rect 6871 9472 6920 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 8570 9500 8576 9512
rect 7024 9472 8576 9500
rect 7024 9432 7052 9472
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 8662 9460 8668 9512
rect 8720 9460 8726 9512
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9500 9183 9503
rect 10042 9500 10048 9512
rect 9171 9472 10048 9500
rect 9171 9469 9183 9472
rect 9125 9463 9183 9469
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 11624 9500 11652 9531
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 12912 9577 12940 9608
rect 13630 9596 13636 9608
rect 13688 9596 13694 9648
rect 14274 9596 14280 9648
rect 14332 9636 14338 9648
rect 14826 9636 14832 9648
rect 14332 9608 14832 9636
rect 14332 9596 14338 9608
rect 14826 9596 14832 9608
rect 14884 9596 14890 9648
rect 15010 9636 15016 9648
rect 14971 9608 15016 9636
rect 15010 9596 15016 9608
rect 15068 9596 15074 9648
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9537 12955 9571
rect 13078 9568 13084 9580
rect 13039 9540 13084 9568
rect 12897 9531 12955 9537
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 13354 9528 13360 9580
rect 13412 9568 13418 9580
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 13412 9540 14197 9568
rect 13412 9528 13418 9540
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 10152 9472 11652 9500
rect 5592 9404 5628 9432
rect 5736 9404 7052 9432
rect 7092 9435 7150 9441
rect 5534 9392 5540 9395
rect 5592 9392 5598 9404
rect 7092 9401 7104 9435
rect 7138 9432 7150 9435
rect 8680 9432 8708 9460
rect 7138 9404 8708 9432
rect 7138 9401 7150 9404
rect 7092 9395 7150 9401
rect 9766 9392 9772 9444
rect 9824 9432 9830 9444
rect 10152 9432 10180 9472
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 13906 9500 13912 9512
rect 12216 9472 13912 9500
rect 12216 9460 12222 9472
rect 13906 9460 13912 9472
rect 13964 9500 13970 9512
rect 14001 9503 14059 9509
rect 14001 9500 14013 9503
rect 13964 9472 14013 9500
rect 13964 9460 13970 9472
rect 14001 9469 14013 9472
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 14642 9460 14648 9512
rect 14700 9500 14706 9512
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 14700 9472 14841 9500
rect 14700 9460 14706 9472
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 9824 9404 10180 9432
rect 10229 9435 10287 9441
rect 9824 9392 9830 9404
rect 10229 9401 10241 9435
rect 10275 9432 10287 9435
rect 11882 9432 11888 9444
rect 10275 9404 11888 9432
rect 10275 9401 10287 9404
rect 10229 9395 10287 9401
rect 11882 9392 11888 9404
rect 11940 9392 11946 9444
rect 6730 9364 6736 9376
rect 5460 9336 6736 9364
rect 5169 9327 5227 9333
rect 6730 9324 6736 9336
rect 6788 9324 6794 9376
rect 7834 9324 7840 9376
rect 7892 9364 7898 9376
rect 8665 9367 8723 9373
rect 8665 9364 8677 9367
rect 7892 9336 8677 9364
rect 7892 9324 7898 9336
rect 8665 9333 8677 9336
rect 8711 9333 8723 9367
rect 8665 9327 8723 9333
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 10321 9367 10379 9373
rect 10321 9364 10333 9367
rect 9732 9336 10333 9364
rect 9732 9324 9738 9336
rect 10321 9333 10333 9336
rect 10367 9364 10379 9367
rect 10410 9364 10416 9376
rect 10367 9336 10416 9364
rect 10367 9333 10379 9336
rect 10321 9327 10379 9333
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 10594 9324 10600 9376
rect 10652 9364 10658 9376
rect 11057 9367 11115 9373
rect 11057 9364 11069 9367
rect 10652 9336 11069 9364
rect 10652 9324 10658 9336
rect 11057 9333 11069 9336
rect 11103 9333 11115 9367
rect 11422 9364 11428 9376
rect 11383 9336 11428 9364
rect 11057 9327 11115 9333
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 11517 9367 11575 9373
rect 11517 9333 11529 9367
rect 11563 9364 11575 9367
rect 12437 9367 12495 9373
rect 12437 9364 12449 9367
rect 11563 9336 12449 9364
rect 11563 9333 11575 9336
rect 11517 9327 11575 9333
rect 12437 9333 12449 9336
rect 12483 9333 12495 9367
rect 12437 9327 12495 9333
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9364 12863 9367
rect 13262 9364 13268 9376
rect 12851 9336 13268 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 13630 9364 13636 9376
rect 13591 9336 13636 9364
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 14090 9324 14096 9376
rect 14148 9364 14154 9376
rect 14148 9336 14193 9364
rect 14148 9324 14154 9336
rect 1104 9274 15824 9296
rect 1104 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 6104 9274
rect 6156 9222 10843 9274
rect 10895 9222 10907 9274
rect 10959 9222 10971 9274
rect 11023 9222 11035 9274
rect 11087 9222 15824 9274
rect 1104 9200 15824 9222
rect 2317 9163 2375 9169
rect 2317 9129 2329 9163
rect 2363 9160 2375 9163
rect 4341 9163 4399 9169
rect 4341 9160 4353 9163
rect 2363 9132 4353 9160
rect 2363 9129 2375 9132
rect 2317 9123 2375 9129
rect 4341 9129 4353 9132
rect 4387 9129 4399 9163
rect 4341 9123 4399 9129
rect 4709 9163 4767 9169
rect 4709 9129 4721 9163
rect 4755 9160 4767 9163
rect 4890 9160 4896 9172
rect 4755 9132 4896 9160
rect 4755 9129 4767 9132
rect 4709 9123 4767 9129
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 5074 9120 5080 9172
rect 5132 9160 5138 9172
rect 10137 9163 10195 9169
rect 10137 9160 10149 9163
rect 5132 9132 10149 9160
rect 5132 9120 5138 9132
rect 10137 9129 10149 9132
rect 10183 9129 10195 9163
rect 10137 9123 10195 9129
rect 11241 9163 11299 9169
rect 11241 9129 11253 9163
rect 11287 9160 11299 9163
rect 11606 9160 11612 9172
rect 11287 9132 11612 9160
rect 11287 9129 11299 9132
rect 11241 9123 11299 9129
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 12069 9163 12127 9169
rect 12069 9129 12081 9163
rect 12115 9160 12127 9163
rect 13722 9160 13728 9172
rect 12115 9132 13728 9160
rect 12115 9129 12127 9132
rect 12069 9123 12127 9129
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 1670 9092 1676 9104
rect 1631 9064 1676 9092
rect 1670 9052 1676 9064
rect 1728 9052 1734 9104
rect 3050 9052 3056 9104
rect 3108 9092 3114 9104
rect 3145 9095 3203 9101
rect 3145 9092 3157 9095
rect 3108 9064 3157 9092
rect 3108 9052 3114 9064
rect 3145 9061 3157 9064
rect 3191 9061 3203 9095
rect 3145 9055 3203 9061
rect 3237 9095 3295 9101
rect 3237 9061 3249 9095
rect 3283 9092 3295 9095
rect 6914 9092 6920 9104
rect 3283 9064 6920 9092
rect 3283 9061 3295 9064
rect 3237 9055 3295 9061
rect 6914 9052 6920 9064
rect 6972 9052 6978 9104
rect 7006 9052 7012 9104
rect 7064 9092 7070 9104
rect 7469 9095 7527 9101
rect 7469 9092 7481 9095
rect 7064 9064 7481 9092
rect 7064 9052 7070 9064
rect 7469 9061 7481 9064
rect 7515 9092 7527 9095
rect 8018 9092 8024 9104
rect 7515 9064 8024 9092
rect 7515 9061 7527 9064
rect 7469 9055 7527 9061
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 8294 9052 8300 9104
rect 8352 9092 8358 9104
rect 9766 9092 9772 9104
rect 8352 9064 9772 9092
rect 8352 9052 8358 9064
rect 9766 9052 9772 9064
rect 9824 9052 9830 9104
rect 10045 9095 10103 9101
rect 10045 9061 10057 9095
rect 10091 9092 10103 9095
rect 10091 9064 11192 9092
rect 10091 9061 10103 9064
rect 10045 9055 10103 9061
rect 11164 9036 11192 9064
rect 11256 9064 11560 9092
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2314 9024 2320 9036
rect 1443 8996 2320 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 5626 9024 5632 9036
rect 2792 8996 5632 9024
rect 2406 8956 2412 8968
rect 2367 8928 2412 8956
rect 2406 8916 2412 8928
rect 2464 8916 2470 8968
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8925 2651 8959
rect 2593 8919 2651 8925
rect 2608 8888 2636 8919
rect 2792 8888 2820 8996
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 5810 9024 5816 9036
rect 5771 8996 5816 9024
rect 5810 8984 5816 8996
rect 5868 8984 5874 9036
rect 6270 8984 6276 9036
rect 6328 9024 6334 9036
rect 6328 8996 7052 9024
rect 6328 8984 6334 8996
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 4430 8956 4436 8968
rect 3467 8928 4436 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 7024 8956 7052 8996
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 7558 9024 7564 9036
rect 7156 8996 7564 9024
rect 7156 8984 7162 8996
rect 7558 8984 7564 8996
rect 7616 9024 7622 9036
rect 7653 9027 7711 9033
rect 7653 9024 7665 9027
rect 7616 8996 7665 9024
rect 7616 8984 7622 8996
rect 7653 8993 7665 8996
rect 7699 8993 7711 9027
rect 7920 9027 7978 9033
rect 7920 9024 7932 9027
rect 7653 8987 7711 8993
rect 7760 8996 7932 9024
rect 7760 8956 7788 8996
rect 7920 8993 7932 8996
rect 7966 9024 7978 9027
rect 7966 8996 10456 9024
rect 7966 8993 7978 8996
rect 7920 8987 7978 8993
rect 5031 8928 6960 8956
rect 7024 8928 7788 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 2608 8860 2820 8888
rect 3050 8848 3056 8900
rect 3108 8888 3114 8900
rect 4154 8888 4160 8900
rect 3108 8860 4160 8888
rect 3108 8848 3114 8860
rect 4154 8848 4160 8860
rect 4212 8848 4218 8900
rect 1946 8820 1952 8832
rect 1907 8792 1952 8820
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 2832 8792 2877 8820
rect 2832 8780 2838 8792
rect 3786 8780 3792 8832
rect 3844 8820 3850 8832
rect 4062 8820 4068 8832
rect 3844 8792 4068 8820
rect 3844 8780 3850 8792
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 4816 8820 4844 8919
rect 4890 8848 4896 8900
rect 4948 8888 4954 8900
rect 6178 8888 6184 8900
rect 4948 8860 6184 8888
rect 4948 8848 4954 8860
rect 6178 8848 6184 8860
rect 6236 8848 6242 8900
rect 6932 8888 6960 8928
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 10321 8959 10379 8965
rect 8812 8928 8953 8956
rect 8812 8916 8818 8928
rect 7558 8888 7564 8900
rect 6932 8860 7564 8888
rect 7558 8848 7564 8860
rect 7616 8848 7622 8900
rect 8925 8888 8953 8928
rect 10321 8925 10333 8959
rect 10367 8925 10379 8959
rect 10428 8956 10456 8996
rect 10502 8984 10508 9036
rect 10560 9024 10566 9036
rect 11054 9024 11060 9036
rect 10560 8996 11060 9024
rect 10560 8984 10566 8996
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 11146 8984 11152 9036
rect 11204 8984 11210 9036
rect 11256 8956 11284 9064
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11388 8996 11433 9024
rect 11388 8984 11394 8996
rect 10428 8928 11284 8956
rect 11425 8959 11483 8965
rect 10321 8919 10379 8925
rect 11425 8925 11437 8959
rect 11471 8925 11483 8959
rect 11532 8956 11560 9064
rect 11698 9052 11704 9104
rect 11756 9092 11762 9104
rect 12434 9092 12440 9104
rect 11756 9064 12440 9092
rect 11756 9052 11762 9064
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 12529 9095 12587 9101
rect 12529 9061 12541 9095
rect 12575 9061 12587 9095
rect 13354 9092 13360 9104
rect 12529 9055 12587 9061
rect 12728 9064 13360 9092
rect 12066 8984 12072 9036
rect 12124 9024 12130 9036
rect 12250 9024 12256 9036
rect 12124 8996 12256 9024
rect 12124 8984 12130 8996
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 12342 8984 12348 9036
rect 12400 9024 12406 9036
rect 12544 9024 12572 9055
rect 12400 8996 12572 9024
rect 12400 8984 12406 8996
rect 12728 8965 12756 9064
rect 13354 9052 13360 9064
rect 13412 9052 13418 9104
rect 12802 8984 12808 9036
rect 12860 9024 12866 9036
rect 13265 9027 13323 9033
rect 13265 9024 13277 9027
rect 12860 8996 13277 9024
rect 12860 8984 12866 8996
rect 13265 8993 13277 8996
rect 13311 8993 13323 9027
rect 14182 9024 14188 9036
rect 14143 8996 14188 9024
rect 13265 8987 13323 8993
rect 14182 8984 14188 8996
rect 14240 8984 14246 9036
rect 12713 8959 12771 8965
rect 12713 8956 12725 8959
rect 11532 8928 12725 8956
rect 11425 8919 11483 8925
rect 12713 8925 12725 8928
rect 12759 8925 12771 8959
rect 12713 8919 12771 8925
rect 9677 8891 9735 8897
rect 9677 8888 9689 8891
rect 8925 8860 9689 8888
rect 9677 8857 9689 8860
rect 9723 8857 9735 8891
rect 10336 8888 10364 8919
rect 10410 8888 10416 8900
rect 10336 8860 10416 8888
rect 9677 8851 9735 8857
rect 10410 8848 10416 8860
rect 10468 8848 10474 8900
rect 10873 8891 10931 8897
rect 10873 8857 10885 8891
rect 10919 8888 10931 8891
rect 11330 8888 11336 8900
rect 10919 8860 11336 8888
rect 10919 8857 10931 8860
rect 10873 8851 10931 8857
rect 11330 8848 11336 8860
rect 11388 8848 11394 8900
rect 11440 8888 11468 8919
rect 12986 8916 12992 8968
rect 13044 8956 13050 8968
rect 13449 8959 13507 8965
rect 13449 8956 13461 8959
rect 13044 8928 13461 8956
rect 13044 8916 13050 8928
rect 13449 8925 13461 8928
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8956 14519 8959
rect 15102 8956 15108 8968
rect 14507 8928 15108 8956
rect 14507 8925 14519 8928
rect 14461 8919 14519 8925
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 13078 8888 13084 8900
rect 11440 8860 13084 8888
rect 6822 8820 6828 8832
rect 4816 8792 6828 8820
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 8018 8820 8024 8832
rect 6972 8792 8024 8820
rect 6972 8780 6978 8792
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 9033 8823 9091 8829
rect 9033 8820 9045 8823
rect 8812 8792 9045 8820
rect 8812 8780 8818 8792
rect 9033 8789 9045 8792
rect 9079 8820 9091 8823
rect 11440 8820 11468 8860
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 15286 8888 15292 8900
rect 13320 8860 15292 8888
rect 13320 8848 13326 8860
rect 15286 8848 15292 8860
rect 15344 8848 15350 8900
rect 9079 8792 11468 8820
rect 9079 8789 9091 8792
rect 9033 8783 9091 8789
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 13170 8820 13176 8832
rect 12492 8792 13176 8820
rect 12492 8780 12498 8792
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 1104 8730 15824 8752
rect 1104 8678 3447 8730
rect 3499 8678 3511 8730
rect 3563 8678 3575 8730
rect 3627 8678 3639 8730
rect 3691 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 13308 8730
rect 13360 8678 13372 8730
rect 13424 8678 13436 8730
rect 13488 8678 13500 8730
rect 13552 8678 15824 8730
rect 1104 8656 15824 8678
rect 1857 8619 1915 8625
rect 1857 8585 1869 8619
rect 1903 8616 1915 8619
rect 2498 8616 2504 8628
rect 1903 8588 2504 8616
rect 1903 8585 1915 8588
rect 1857 8579 1915 8585
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 2682 8616 2688 8628
rect 2643 8588 2688 8616
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 3142 8576 3148 8628
rect 3200 8616 3206 8628
rect 4065 8619 4123 8625
rect 4065 8616 4077 8619
rect 3200 8588 4077 8616
rect 3200 8576 3206 8588
rect 4065 8585 4077 8588
rect 4111 8585 4123 8619
rect 4065 8579 4123 8585
rect 4430 8576 4436 8628
rect 4488 8616 4494 8628
rect 6270 8616 6276 8628
rect 4488 8588 5847 8616
rect 6231 8588 6276 8616
rect 4488 8576 4494 8588
rect 5819 8548 5847 8588
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 7098 8616 7104 8628
rect 6840 8588 7104 8616
rect 3252 8520 4752 8548
rect 5819 8520 6408 8548
rect 2498 8480 2504 8492
rect 2459 8452 2504 8480
rect 2498 8440 2504 8452
rect 2556 8440 2562 8492
rect 3252 8489 3280 8520
rect 4724 8492 4752 8520
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 3697 8483 3755 8489
rect 3697 8480 3709 8483
rect 3384 8452 3709 8480
rect 3384 8440 3390 8452
rect 3697 8449 3709 8452
rect 3743 8449 3755 8483
rect 4522 8480 4528 8492
rect 4483 8452 4528 8480
rect 3697 8443 3755 8449
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 4706 8480 4712 8492
rect 4667 8452 4712 8480
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8412 2283 8415
rect 2314 8412 2320 8424
rect 2271 8384 2320 8412
rect 2271 8381 2283 8384
rect 2225 8375 2283 8381
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 2958 8372 2964 8424
rect 3016 8412 3022 8424
rect 3513 8415 3571 8421
rect 3513 8412 3525 8415
rect 3016 8384 3525 8412
rect 3016 8372 3022 8384
rect 3513 8381 3525 8384
rect 3559 8381 3571 8415
rect 4890 8412 4896 8424
rect 4851 8384 4896 8412
rect 3513 8375 3571 8381
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 5534 8412 5540 8424
rect 5092 8384 5540 8412
rect 3145 8347 3203 8353
rect 3145 8313 3157 8347
rect 3191 8344 3203 8347
rect 4338 8344 4344 8356
rect 3191 8316 4344 8344
rect 3191 8313 3203 8316
rect 3145 8307 3203 8313
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 4433 8347 4491 8353
rect 4433 8313 4445 8347
rect 4479 8344 4491 8347
rect 5092 8344 5120 8384
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 6380 8412 6408 8520
rect 6840 8489 6868 8588
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 7616 8588 10057 8616
rect 7616 8576 7622 8588
rect 10045 8585 10057 8588
rect 10091 8616 10103 8619
rect 10410 8616 10416 8628
rect 10091 8588 10416 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 11422 8616 11428 8628
rect 10652 8588 11428 8616
rect 10652 8576 10658 8588
rect 11422 8576 11428 8588
rect 11480 8576 11486 8628
rect 12434 8616 12440 8628
rect 12395 8588 12440 8616
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 14458 8616 14464 8628
rect 12912 8588 14464 8616
rect 8205 8551 8263 8557
rect 8205 8517 8217 8551
rect 8251 8548 8263 8551
rect 8294 8548 8300 8560
rect 8251 8520 8300 8548
rect 8251 8517 8263 8520
rect 8205 8511 8263 8517
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 10505 8551 10563 8557
rect 10505 8548 10517 8551
rect 9692 8520 10517 8548
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 6825 8443 6883 8449
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 7984 8452 8791 8480
rect 7984 8440 7990 8452
rect 6380 8384 6859 8412
rect 4479 8316 5120 8344
rect 5160 8347 5218 8353
rect 4479 8313 4491 8316
rect 4433 8307 4491 8313
rect 5160 8313 5172 8347
rect 5206 8344 5218 8347
rect 5626 8344 5632 8356
rect 5206 8316 5632 8344
rect 5206 8313 5218 8316
rect 5160 8307 5218 8313
rect 5626 8304 5632 8316
rect 5684 8344 5690 8356
rect 6730 8344 6736 8356
rect 5684 8316 6736 8344
rect 5684 8304 5690 8316
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 6831 8344 6859 8384
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 7081 8415 7139 8421
rect 7081 8412 7093 8415
rect 6972 8384 7093 8412
rect 6972 8372 6978 8384
rect 7081 8381 7093 8384
rect 7127 8412 7139 8415
rect 8478 8412 8484 8424
rect 7127 8384 8484 8412
rect 7127 8381 7139 8384
rect 7081 8375 7139 8381
rect 8478 8372 8484 8384
rect 8536 8372 8542 8424
rect 8662 8412 8668 8424
rect 8623 8384 8668 8412
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 8763 8412 8791 8452
rect 9692 8412 9720 8520
rect 10505 8517 10517 8520
rect 10551 8517 10563 8551
rect 10505 8511 10563 8517
rect 10962 8508 10968 8560
rect 11020 8548 11026 8560
rect 11974 8548 11980 8560
rect 11020 8520 11980 8548
rect 11020 8508 11026 8520
rect 11974 8508 11980 8520
rect 12032 8508 12038 8560
rect 10778 8440 10784 8492
rect 10836 8480 10842 8492
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10836 8452 11069 8480
rect 10836 8440 10842 8452
rect 11057 8449 11069 8452
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 12912 8489 12940 8588
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 13633 8551 13691 8557
rect 13633 8517 13645 8551
rect 13679 8548 13691 8551
rect 14274 8548 14280 8560
rect 13679 8520 14280 8548
rect 13679 8517 13691 8520
rect 13633 8511 13691 8517
rect 14274 8508 14280 8520
rect 14332 8508 14338 8560
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11664 8452 11713 8480
rect 11664 8440 11670 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8480 13139 8483
rect 13446 8480 13452 8492
rect 13127 8452 13452 8480
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 8763 8384 9720 8412
rect 10042 8372 10048 8424
rect 10100 8412 10106 8424
rect 10965 8415 11023 8421
rect 10965 8412 10977 8415
rect 10100 8384 10977 8412
rect 10100 8372 10106 8384
rect 10965 8381 10977 8384
rect 11011 8412 11023 8415
rect 12912 8412 12940 8443
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 14185 8483 14243 8489
rect 14185 8480 14197 8483
rect 13780 8452 14197 8480
rect 13780 8440 13786 8452
rect 14185 8449 14197 8452
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 11011 8384 12940 8412
rect 14093 8415 14151 8421
rect 11011 8381 11023 8384
rect 10965 8375 11023 8381
rect 14093 8381 14105 8415
rect 14139 8412 14151 8415
rect 14366 8412 14372 8424
rect 14139 8384 14372 8412
rect 14139 8381 14151 8384
rect 14093 8375 14151 8381
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 14734 8372 14740 8424
rect 14792 8412 14798 8424
rect 14829 8415 14887 8421
rect 14829 8412 14841 8415
rect 14792 8384 14841 8412
rect 14792 8372 14798 8384
rect 14829 8381 14841 8384
rect 14875 8381 14887 8415
rect 14829 8375 14887 8381
rect 6831 8316 8156 8344
rect 2314 8236 2320 8288
rect 2372 8276 2378 8288
rect 2372 8248 2417 8276
rect 2372 8236 2378 8248
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3053 8279 3111 8285
rect 3053 8276 3065 8279
rect 3016 8248 3065 8276
rect 3016 8236 3022 8248
rect 3053 8245 3065 8248
rect 3099 8245 3111 8279
rect 3053 8239 3111 8245
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 4614 8276 4620 8288
rect 3476 8248 4620 8276
rect 3476 8236 3482 8248
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 7834 8276 7840 8288
rect 4948 8248 7840 8276
rect 4948 8236 4954 8248
rect 7834 8236 7840 8248
rect 7892 8236 7898 8288
rect 8128 8276 8156 8316
rect 8202 8304 8208 8356
rect 8260 8344 8266 8356
rect 8910 8347 8968 8353
rect 8910 8344 8922 8347
rect 8260 8316 8922 8344
rect 8260 8304 8266 8316
rect 8910 8313 8922 8316
rect 8956 8344 8968 8347
rect 8956 8316 10364 8344
rect 8956 8313 8968 8316
rect 8910 8307 8968 8313
rect 9582 8276 9588 8288
rect 8128 8248 9588 8276
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 10336 8276 10364 8316
rect 10410 8304 10416 8356
rect 10468 8344 10474 8356
rect 10873 8347 10931 8353
rect 10873 8344 10885 8347
rect 10468 8316 10885 8344
rect 10468 8304 10474 8316
rect 10873 8313 10885 8316
rect 10919 8313 10931 8347
rect 10873 8307 10931 8313
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 14001 8347 14059 8353
rect 14001 8344 14013 8347
rect 11112 8316 14013 8344
rect 11112 8304 11118 8316
rect 14001 8313 14013 8316
rect 14047 8313 14059 8347
rect 14001 8307 14059 8313
rect 10686 8276 10692 8288
rect 10336 8248 10692 8276
rect 10686 8236 10692 8248
rect 10744 8236 10750 8288
rect 12802 8276 12808 8288
rect 12763 8248 12808 8276
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 14458 8276 14464 8288
rect 13504 8248 14464 8276
rect 13504 8236 13510 8248
rect 14458 8236 14464 8248
rect 14516 8236 14522 8288
rect 14642 8236 14648 8288
rect 14700 8276 14706 8288
rect 15013 8279 15071 8285
rect 15013 8276 15025 8279
rect 14700 8248 15025 8276
rect 14700 8236 14706 8248
rect 15013 8245 15025 8248
rect 15059 8245 15071 8279
rect 15013 8239 15071 8245
rect 1104 8186 15824 8208
rect 1104 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 6104 8186
rect 6156 8134 10843 8186
rect 10895 8134 10907 8186
rect 10959 8134 10971 8186
rect 11023 8134 11035 8186
rect 11087 8134 15824 8186
rect 1104 8112 15824 8134
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 2409 8075 2467 8081
rect 2409 8072 2421 8075
rect 2372 8044 2421 8072
rect 2372 8032 2378 8044
rect 2409 8041 2421 8044
rect 2455 8041 2467 8075
rect 2409 8035 2467 8041
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 2869 8075 2927 8081
rect 2869 8072 2881 8075
rect 2832 8044 2881 8072
rect 2832 8032 2838 8044
rect 2869 8041 2881 8044
rect 2915 8041 2927 8075
rect 2869 8035 2927 8041
rect 4065 8075 4123 8081
rect 4065 8041 4077 8075
rect 4111 8072 4123 8075
rect 6546 8072 6552 8084
rect 4111 8044 6552 8072
rect 4111 8041 4123 8044
rect 4065 8035 4123 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 8849 8075 8907 8081
rect 8849 8072 8861 8075
rect 6788 8044 8861 8072
rect 6788 8032 6794 8044
rect 8849 8041 8861 8044
rect 8895 8041 8907 8075
rect 8849 8035 8907 8041
rect 9766 8032 9772 8084
rect 9824 8072 9830 8084
rect 10226 8072 10232 8084
rect 9824 8044 10232 8072
rect 9824 8032 9830 8044
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 10652 8044 11100 8072
rect 10652 8032 10658 8044
rect 2498 7964 2504 8016
rect 2556 8004 2562 8016
rect 7006 8004 7012 8016
rect 2556 7976 3648 8004
rect 2556 7964 2562 7976
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7905 2007 7939
rect 1949 7899 2007 7905
rect 1964 7800 1992 7899
rect 2038 7896 2044 7948
rect 2096 7936 2102 7948
rect 2096 7908 2141 7936
rect 2096 7896 2102 7908
rect 2774 7896 2780 7948
rect 2832 7936 2838 7948
rect 2832 7908 2877 7936
rect 2832 7896 2838 7908
rect 2958 7896 2964 7948
rect 3016 7936 3022 7948
rect 3418 7936 3424 7948
rect 3016 7908 3424 7936
rect 3016 7896 3022 7908
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7868 2283 7871
rect 2682 7868 2688 7880
rect 2271 7840 2688 7868
rect 2271 7837 2283 7840
rect 2225 7831 2283 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3142 7868 3148 7880
rect 3099 7840 3148 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3620 7868 3648 7976
rect 3804 7976 5396 8004
rect 3804 7948 3832 7976
rect 3786 7936 3792 7948
rect 3699 7908 3792 7936
rect 3786 7896 3792 7908
rect 3844 7896 3850 7948
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 5074 7936 5080 7948
rect 4479 7908 5080 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 4338 7868 4344 7880
rect 3620 7840 4344 7868
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4522 7868 4528 7880
rect 4483 7840 4528 7868
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7868 4767 7871
rect 5258 7868 5264 7880
rect 4755 7840 5264 7868
rect 4755 7837 4767 7840
rect 4709 7831 4767 7837
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5368 7868 5396 7976
rect 5460 7976 7012 8004
rect 5460 7945 5488 7976
rect 7006 7964 7012 7976
rect 7064 7964 7070 8016
rect 7282 7964 7288 8016
rect 7340 7964 7346 8016
rect 7558 7964 7564 8016
rect 7616 8004 7622 8016
rect 7714 8007 7772 8013
rect 7714 8004 7726 8007
rect 7616 7976 7726 8004
rect 7616 7964 7622 7976
rect 7714 7973 7726 7976
rect 7760 7973 7772 8007
rect 7714 7967 7772 7973
rect 7834 7964 7840 8016
rect 7892 8004 7898 8016
rect 8570 8004 8576 8016
rect 7892 7976 8576 8004
rect 7892 7964 7898 7976
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 5445 7939 5503 7945
rect 5445 7905 5457 7939
rect 5491 7905 5503 7939
rect 5626 7936 5632 7948
rect 5587 7908 5632 7936
rect 5445 7899 5503 7905
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 5896 7939 5954 7945
rect 5896 7905 5908 7939
rect 5942 7936 5954 7939
rect 7300 7936 7328 7964
rect 7469 7939 7527 7945
rect 7469 7936 7481 7939
rect 5942 7908 7328 7936
rect 7372 7908 7481 7936
rect 5942 7905 5954 7908
rect 5896 7899 5954 7905
rect 5368 7840 5571 7868
rect 5442 7800 5448 7812
rect 1964 7772 5448 7800
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 3326 7732 3332 7744
rect 1627 7704 3332 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 3326 7692 3332 7704
rect 3384 7692 3390 7744
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 3970 7732 3976 7744
rect 3651 7704 3976 7732
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 3970 7692 3976 7704
rect 4028 7692 4034 7744
rect 5258 7732 5264 7744
rect 5219 7704 5264 7732
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 5543 7732 5571 7840
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 7372 7868 7400 7908
rect 7469 7905 7481 7908
rect 7515 7905 7527 7939
rect 9493 7939 9551 7945
rect 9493 7936 9505 7939
rect 7469 7899 7527 7905
rect 7576 7908 9505 7936
rect 7576 7868 7604 7908
rect 9493 7905 9505 7908
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 9582 7896 9588 7948
rect 9640 7936 9646 7948
rect 9933 7939 9991 7945
rect 9933 7936 9945 7939
rect 9640 7908 9945 7936
rect 9640 7896 9646 7908
rect 9933 7905 9945 7908
rect 9979 7936 9991 7939
rect 10502 7936 10508 7948
rect 9979 7908 10508 7936
rect 9979 7905 9991 7908
rect 9933 7899 9991 7905
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 11072 7936 11100 8044
rect 11146 8032 11152 8084
rect 11204 8072 11210 8084
rect 11517 8075 11575 8081
rect 11517 8072 11529 8075
rect 11204 8044 11529 8072
rect 11204 8032 11210 8044
rect 11517 8041 11529 8044
rect 11563 8041 11575 8075
rect 11517 8035 11575 8041
rect 11606 8032 11612 8084
rect 11664 8072 11670 8084
rect 11885 8075 11943 8081
rect 11885 8072 11897 8075
rect 11664 8044 11897 8072
rect 11664 8032 11670 8044
rect 11885 8041 11897 8044
rect 11931 8072 11943 8075
rect 12342 8072 12348 8084
rect 11931 8044 12348 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 13081 8075 13139 8081
rect 13081 8041 13093 8075
rect 13127 8072 13139 8075
rect 13170 8072 13176 8084
rect 13127 8044 13176 8072
rect 13127 8041 13139 8044
rect 13081 8035 13139 8041
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 14274 8072 14280 8084
rect 14235 8044 14280 8072
rect 14274 8032 14280 8044
rect 14332 8032 14338 8084
rect 11974 8004 11980 8016
rect 11935 7976 11980 8004
rect 11974 7964 11980 7976
rect 12032 7964 12038 8016
rect 11882 7936 11888 7948
rect 11072 7908 11888 7936
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 12526 7896 12532 7948
rect 12584 7936 12590 7948
rect 12584 7908 13308 7936
rect 12584 7896 12590 7908
rect 6788 7840 7400 7868
rect 7484 7840 7604 7868
rect 6788 7828 6794 7840
rect 7484 7800 7512 7840
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 9677 7871 9735 7877
rect 8628 7840 9352 7868
rect 8628 7828 8634 7840
rect 9324 7809 9352 7840
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 9309 7803 9367 7809
rect 6564 7772 7512 7800
rect 8680 7772 9076 7800
rect 6564 7732 6592 7772
rect 5543 7704 6592 7732
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7009 7735 7067 7741
rect 7009 7732 7021 7735
rect 6972 7704 7021 7732
rect 6972 7692 6978 7704
rect 7009 7701 7021 7704
rect 7055 7732 7067 7735
rect 8680 7732 8708 7772
rect 7055 7704 8708 7732
rect 7055 7701 7067 7704
rect 7009 7695 7067 7701
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 8938 7732 8944 7744
rect 8812 7704 8944 7732
rect 8812 7692 8818 7704
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 9048 7732 9076 7772
rect 9309 7769 9321 7803
rect 9355 7769 9367 7803
rect 9309 7763 9367 7769
rect 9490 7760 9496 7812
rect 9548 7800 9554 7812
rect 9692 7800 9720 7831
rect 10686 7828 10692 7880
rect 10744 7868 10750 7880
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 10744 7840 12081 7868
rect 10744 7828 10750 7840
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 13170 7868 13176 7880
rect 13131 7840 13176 7868
rect 12069 7831 12127 7837
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 13280 7877 13308 7908
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7837 13323 7871
rect 13265 7831 13323 7837
rect 13630 7828 13636 7880
rect 13688 7868 13694 7880
rect 14369 7871 14427 7877
rect 14369 7868 14381 7871
rect 13688 7840 14381 7868
rect 13688 7828 13694 7840
rect 14369 7837 14381 7840
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 15378 7868 15384 7880
rect 14599 7840 15384 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 14568 7800 14596 7831
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 9548 7772 9720 7800
rect 10612 7772 14596 7800
rect 9548 7760 9554 7772
rect 10612 7732 10640 7772
rect 9048 7704 10640 7732
rect 11057 7735 11115 7741
rect 11057 7701 11069 7735
rect 11103 7732 11115 7735
rect 11146 7732 11152 7744
rect 11103 7704 11152 7732
rect 11103 7701 11115 7704
rect 11057 7695 11115 7701
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 11606 7692 11612 7744
rect 11664 7732 11670 7744
rect 12713 7735 12771 7741
rect 12713 7732 12725 7735
rect 11664 7704 12725 7732
rect 11664 7692 11670 7704
rect 12713 7701 12725 7704
rect 12759 7701 12771 7735
rect 13906 7732 13912 7744
rect 13867 7704 13912 7732
rect 12713 7695 12771 7701
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 13998 7692 14004 7744
rect 14056 7732 14062 7744
rect 14366 7732 14372 7744
rect 14056 7704 14372 7732
rect 14056 7692 14062 7704
rect 14366 7692 14372 7704
rect 14424 7692 14430 7744
rect 1104 7642 15824 7664
rect 1104 7590 3447 7642
rect 3499 7590 3511 7642
rect 3563 7590 3575 7642
rect 3627 7590 3639 7642
rect 3691 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 13308 7642
rect 13360 7590 13372 7642
rect 13424 7590 13436 7642
rect 13488 7590 13500 7642
rect 13552 7590 15824 7642
rect 1104 7568 15824 7590
rect 5994 7528 6000 7540
rect 3068 7500 6000 7528
rect 2225 7463 2283 7469
rect 2225 7429 2237 7463
rect 2271 7460 2283 7463
rect 2958 7460 2964 7472
rect 2271 7432 2964 7460
rect 2271 7429 2283 7432
rect 2225 7423 2283 7429
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 1486 7352 1492 7404
rect 1544 7392 1550 7404
rect 1670 7392 1676 7404
rect 1544 7364 1676 7392
rect 1544 7352 1550 7364
rect 1670 7352 1676 7364
rect 1728 7392 1734 7404
rect 1857 7395 1915 7401
rect 1857 7392 1869 7395
rect 1728 7364 1869 7392
rect 1728 7352 1734 7364
rect 1857 7361 1869 7364
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7392 2099 7395
rect 2498 7392 2504 7404
rect 2087 7364 2504 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7392 2927 7395
rect 3068 7392 3096 7500
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 6270 7528 6276 7540
rect 6231 7500 6276 7528
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 10505 7531 10563 7537
rect 10505 7528 10517 7531
rect 6880 7500 8432 7528
rect 6880 7488 6886 7500
rect 4338 7420 4344 7472
rect 4396 7460 4402 7472
rect 4433 7463 4491 7469
rect 4433 7460 4445 7463
rect 4396 7432 4445 7460
rect 4396 7420 4402 7432
rect 4433 7429 4445 7432
rect 4479 7429 4491 7463
rect 4433 7423 4491 7429
rect 5902 7420 5908 7472
rect 5960 7460 5966 7472
rect 6178 7460 6184 7472
rect 5960 7432 6184 7460
rect 5960 7420 5966 7432
rect 6178 7420 6184 7432
rect 6236 7420 6242 7472
rect 8205 7463 8263 7469
rect 8205 7460 8217 7463
rect 7944 7432 8217 7460
rect 4890 7392 4896 7404
rect 2915 7364 3096 7392
rect 4851 7364 4896 7392
rect 2915 7361 2927 7364
rect 2869 7355 2927 7361
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 6822 7392 6828 7404
rect 5911 7364 6572 7392
rect 6783 7364 6828 7392
rect 1762 7284 1768 7336
rect 1820 7324 1826 7336
rect 2222 7324 2228 7336
rect 1820 7296 2228 7324
rect 1820 7284 1826 7296
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 2406 7284 2412 7336
rect 2464 7324 2470 7336
rect 3053 7327 3111 7333
rect 3053 7324 3065 7327
rect 2464 7296 3065 7324
rect 2464 7284 2470 7296
rect 3053 7293 3065 7296
rect 3099 7324 3111 7327
rect 4908 7324 4936 7352
rect 5911 7324 5939 7364
rect 3099 7296 4936 7324
rect 5000 7296 5939 7324
rect 3099 7293 3111 7296
rect 3053 7287 3111 7293
rect 2593 7259 2651 7265
rect 2593 7225 2605 7259
rect 2639 7256 2651 7259
rect 2774 7256 2780 7268
rect 2639 7228 2780 7256
rect 2639 7225 2651 7228
rect 2593 7219 2651 7225
rect 2774 7216 2780 7228
rect 2832 7216 2838 7268
rect 3142 7216 3148 7268
rect 3200 7256 3206 7268
rect 3320 7259 3378 7265
rect 3320 7256 3332 7259
rect 3200 7228 3332 7256
rect 3200 7216 3206 7228
rect 3320 7225 3332 7228
rect 3366 7256 3378 7259
rect 5000 7256 5028 7296
rect 5994 7284 6000 7336
rect 6052 7324 6058 7336
rect 6544 7324 6572 7364
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 7944 7336 7972 7432
rect 8205 7429 8217 7432
rect 8251 7429 8263 7463
rect 8404 7460 8432 7500
rect 8588 7500 10517 7528
rect 8588 7460 8616 7500
rect 10505 7497 10517 7500
rect 10551 7497 10563 7531
rect 10505 7491 10563 7497
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 12437 7531 12495 7537
rect 12437 7528 12449 7531
rect 11112 7500 12449 7528
rect 11112 7488 11118 7500
rect 12437 7497 12449 7500
rect 12483 7497 12495 7531
rect 12437 7491 12495 7497
rect 12986 7488 12992 7540
rect 13044 7488 13050 7540
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 13633 7531 13691 7537
rect 13633 7528 13645 7531
rect 13228 7500 13645 7528
rect 13228 7488 13234 7500
rect 13633 7497 13645 7500
rect 13679 7497 13691 7531
rect 13633 7491 13691 7497
rect 14734 7488 14740 7540
rect 14792 7528 14798 7540
rect 14918 7528 14924 7540
rect 14792 7500 14924 7528
rect 14792 7488 14798 7500
rect 14918 7488 14924 7500
rect 14976 7488 14982 7540
rect 8404 7432 8616 7460
rect 8205 7423 8263 7429
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 13004 7460 13032 7488
rect 9732 7432 13032 7460
rect 9732 7420 9738 7432
rect 13262 7420 13268 7472
rect 13320 7460 13326 7472
rect 15013 7463 15071 7469
rect 15013 7460 15025 7463
rect 13320 7432 15025 7460
rect 13320 7420 13326 7432
rect 15013 7429 15025 7432
rect 15059 7429 15071 7463
rect 15013 7423 15071 7429
rect 10226 7352 10232 7404
rect 10284 7392 10290 7404
rect 10502 7392 10508 7404
rect 10284 7364 10508 7392
rect 10284 7352 10290 7364
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 10686 7352 10692 7404
rect 10744 7392 10750 7404
rect 11057 7395 11115 7401
rect 11057 7392 11069 7395
rect 10744 7364 11069 7392
rect 10744 7352 10750 7364
rect 11057 7361 11069 7364
rect 11103 7361 11115 7395
rect 11057 7355 11115 7361
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12434 7392 12440 7404
rect 12124 7364 12440 7392
rect 12124 7352 12130 7364
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12676 7364 13001 7392
rect 12676 7352 12682 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13354 7352 13360 7404
rect 13412 7392 13418 7404
rect 14093 7395 14151 7401
rect 14093 7392 14105 7395
rect 13412 7364 14105 7392
rect 13412 7352 13418 7364
rect 14093 7361 14105 7364
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7392 14335 7395
rect 14458 7392 14464 7404
rect 14323 7364 14464 7392
rect 14323 7361 14335 7364
rect 14277 7355 14335 7361
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 14550 7352 14556 7404
rect 14608 7392 14614 7404
rect 14608 7364 14964 7392
rect 14608 7352 14614 7364
rect 7466 7324 7472 7336
rect 6052 7296 6500 7324
rect 6544 7296 7472 7324
rect 6052 7284 6058 7296
rect 5166 7265 5172 7268
rect 5160 7256 5172 7265
rect 3366 7228 5028 7256
rect 5127 7228 5172 7256
rect 3366 7225 3378 7228
rect 3320 7219 3378 7225
rect 5160 7219 5172 7228
rect 5166 7216 5172 7219
rect 5224 7216 5230 7268
rect 5442 7216 5448 7268
rect 5500 7256 5506 7268
rect 6472 7256 6500 7296
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 7926 7284 7932 7336
rect 7984 7284 7990 7336
rect 8018 7284 8024 7336
rect 8076 7324 8082 7336
rect 8662 7324 8668 7336
rect 8076 7296 8668 7324
rect 8076 7284 8082 7296
rect 8662 7284 8668 7296
rect 8720 7324 8726 7336
rect 9490 7324 9496 7336
rect 8720 7296 9496 7324
rect 8720 7284 8726 7296
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 10042 7284 10048 7336
rect 10100 7324 10106 7336
rect 10410 7324 10416 7336
rect 10100 7296 10416 7324
rect 10100 7284 10106 7296
rect 10410 7284 10416 7296
rect 10468 7284 10474 7336
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 11606 7324 11612 7336
rect 10919 7296 11612 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 11606 7284 11612 7296
rect 11664 7284 11670 7336
rect 12710 7324 12716 7336
rect 12268 7296 12716 7324
rect 7098 7265 7104 7268
rect 7092 7256 7104 7265
rect 5500 7228 6408 7256
rect 6472 7228 7104 7256
rect 5500 7216 5506 7228
rect 1397 7191 1455 7197
rect 1397 7157 1409 7191
rect 1443 7188 1455 7191
rect 1578 7188 1584 7200
rect 1443 7160 1584 7188
rect 1443 7157 1455 7160
rect 1397 7151 1455 7157
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 1762 7188 1768 7200
rect 1723 7160 1768 7188
rect 1762 7148 1768 7160
rect 1820 7148 1826 7200
rect 2685 7191 2743 7197
rect 2685 7157 2697 7191
rect 2731 7188 2743 7191
rect 4062 7188 4068 7200
rect 2731 7160 4068 7188
rect 2731 7157 2743 7160
rect 2685 7151 2743 7157
rect 4062 7148 4068 7160
rect 4120 7148 4126 7200
rect 4706 7148 4712 7200
rect 4764 7188 4770 7200
rect 5175 7188 5203 7216
rect 4764 7160 5203 7188
rect 4764 7148 4770 7160
rect 5350 7148 5356 7200
rect 5408 7188 5414 7200
rect 6270 7188 6276 7200
rect 5408 7160 6276 7188
rect 5408 7148 5414 7160
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 6380 7188 6408 7228
rect 7092 7219 7104 7228
rect 7098 7216 7104 7219
rect 7156 7216 7162 7268
rect 8910 7259 8968 7265
rect 8910 7256 8922 7259
rect 7208 7228 8922 7256
rect 7208 7188 7236 7228
rect 8910 7225 8922 7228
rect 8956 7225 8968 7259
rect 11146 7256 11152 7268
rect 8910 7219 8968 7225
rect 9048 7228 11152 7256
rect 6380 7160 7236 7188
rect 7282 7148 7288 7200
rect 7340 7188 7346 7200
rect 7466 7188 7472 7200
rect 7340 7160 7472 7188
rect 7340 7148 7346 7160
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 8110 7148 8116 7200
rect 8168 7188 8174 7200
rect 9048 7188 9076 7228
rect 11146 7216 11152 7228
rect 11204 7216 11210 7268
rect 11701 7259 11759 7265
rect 11701 7225 11713 7259
rect 11747 7256 11759 7259
rect 12268 7256 12296 7296
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 12894 7324 12900 7336
rect 12851 7296 12900 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 13170 7284 13176 7336
rect 13228 7324 13234 7336
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 13228 7296 14841 7324
rect 13228 7284 13234 7296
rect 14829 7293 14841 7296
rect 14875 7293 14887 7327
rect 14829 7287 14887 7293
rect 14090 7256 14096 7268
rect 11747 7228 12296 7256
rect 12912 7228 14096 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 8168 7160 9076 7188
rect 8168 7148 8174 7160
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 10045 7191 10103 7197
rect 10045 7188 10057 7191
rect 9824 7160 10057 7188
rect 9824 7148 9830 7160
rect 10045 7157 10057 7160
rect 10091 7157 10103 7191
rect 10045 7151 10103 7157
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10410 7188 10416 7200
rect 10192 7160 10416 7188
rect 10192 7148 10198 7160
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 12250 7188 12256 7200
rect 11011 7160 12256 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 12912 7197 12940 7228
rect 14090 7216 14096 7228
rect 14148 7256 14154 7268
rect 14550 7256 14556 7268
rect 14148 7228 14556 7256
rect 14148 7216 14154 7228
rect 14550 7216 14556 7228
rect 14608 7216 14614 7268
rect 12897 7191 12955 7197
rect 12897 7157 12909 7191
rect 12943 7157 12955 7191
rect 12897 7151 12955 7157
rect 13262 7148 13268 7200
rect 13320 7188 13326 7200
rect 14001 7191 14059 7197
rect 14001 7188 14013 7191
rect 13320 7160 14013 7188
rect 13320 7148 13326 7160
rect 14001 7157 14013 7160
rect 14047 7188 14059 7191
rect 14936 7188 14964 7364
rect 15930 7188 15936 7200
rect 14047 7160 15936 7188
rect 14047 7157 14059 7160
rect 14001 7151 14059 7157
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 1104 7098 15824 7120
rect 1104 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 6104 7098
rect 6156 7046 10843 7098
rect 10895 7046 10907 7098
rect 10959 7046 10971 7098
rect 11023 7046 11035 7098
rect 11087 7046 15824 7098
rect 1104 7024 15824 7046
rect 1762 6944 1768 6996
rect 1820 6984 1826 6996
rect 2314 6984 2320 6996
rect 1820 6956 2320 6984
rect 1820 6944 1826 6956
rect 2314 6944 2320 6956
rect 2372 6984 2378 6996
rect 3050 6984 3056 6996
rect 2372 6956 3056 6984
rect 2372 6944 2378 6956
rect 3050 6944 3056 6956
rect 3108 6944 3114 6996
rect 4430 6984 4436 6996
rect 4391 6956 4436 6984
rect 4430 6944 4436 6956
rect 4488 6944 4494 6996
rect 5166 6944 5172 6996
rect 5224 6984 5230 6996
rect 9766 6984 9772 6996
rect 5224 6956 9772 6984
rect 5224 6944 5230 6956
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 10594 6944 10600 6996
rect 10652 6984 10658 6996
rect 11057 6987 11115 6993
rect 11057 6984 11069 6987
rect 10652 6956 11069 6984
rect 10652 6944 10658 6956
rect 11057 6953 11069 6956
rect 11103 6984 11115 6987
rect 12618 6984 12624 6996
rect 11103 6956 12624 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 12618 6944 12624 6956
rect 12676 6944 12682 6996
rect 1578 6876 1584 6928
rect 1636 6916 1642 6928
rect 4614 6916 4620 6928
rect 1636 6888 4620 6916
rect 1636 6876 1642 6888
rect 4614 6876 4620 6888
rect 4672 6876 4678 6928
rect 5350 6916 5356 6928
rect 4724 6888 5356 6916
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 2400 6851 2458 6857
rect 2400 6817 2412 6851
rect 2446 6848 2458 6851
rect 2682 6848 2688 6860
rect 2446 6820 2688 6848
rect 2446 6817 2458 6820
rect 2400 6811 2458 6817
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 4430 6740 4436 6792
rect 4488 6780 4494 6792
rect 4724 6789 4752 6888
rect 5350 6876 5356 6888
rect 5408 6876 5414 6928
rect 6822 6876 6828 6928
rect 6880 6916 6886 6928
rect 7650 6916 7656 6928
rect 6880 6888 7656 6916
rect 6880 6876 6886 6888
rect 5528 6851 5586 6857
rect 5528 6817 5540 6851
rect 5574 6848 5586 6851
rect 6086 6848 6092 6860
rect 5574 6820 6092 6848
rect 5574 6817 5586 6820
rect 5528 6811 5586 6817
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 7107 6857 7135 6888
rect 7650 6876 7656 6888
rect 7708 6876 7714 6928
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 8938 6916 8944 6928
rect 8352 6888 8944 6916
rect 8352 6876 8358 6888
rect 8938 6876 8944 6888
rect 8996 6876 9002 6928
rect 9030 6876 9036 6928
rect 9088 6916 9094 6928
rect 11885 6919 11943 6925
rect 9088 6888 9133 6916
rect 9088 6876 9094 6888
rect 11885 6885 11897 6919
rect 11931 6916 11943 6919
rect 12434 6916 12440 6928
rect 11931 6888 12440 6916
rect 11931 6885 11943 6888
rect 11885 6879 11943 6885
rect 12434 6876 12440 6888
rect 12492 6876 12498 6928
rect 12802 6916 12808 6928
rect 12544 6888 12808 6916
rect 7101 6851 7159 6857
rect 7101 6817 7113 6851
rect 7147 6817 7159 6851
rect 7357 6851 7415 6857
rect 7357 6848 7369 6851
rect 7101 6811 7159 6817
rect 7208 6820 7369 6848
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 4488 6752 4537 6780
rect 4488 6740 4494 6752
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6749 4767 6783
rect 4709 6743 4767 6749
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5166 6780 5172 6792
rect 4948 6752 5172 6780
rect 4948 6740 4954 6752
rect 5166 6740 5172 6752
rect 5224 6780 5230 6792
rect 5261 6783 5319 6789
rect 5261 6780 5273 6783
rect 5224 6752 5273 6780
rect 5224 6740 5230 6752
rect 5261 6749 5273 6752
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 6270 6740 6276 6792
rect 6328 6780 6334 6792
rect 7208 6780 7236 6820
rect 7357 6817 7369 6820
rect 7403 6848 7415 6851
rect 7926 6848 7932 6860
rect 7403 6820 7932 6848
rect 7403 6817 7415 6820
rect 7357 6811 7415 6817
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 9766 6848 9772 6860
rect 8303 6820 9772 6848
rect 8303 6780 8331 6820
rect 9766 6808 9772 6820
rect 9824 6848 9830 6860
rect 9933 6851 9991 6857
rect 9933 6848 9945 6851
rect 9824 6820 9945 6848
rect 9824 6808 9830 6820
rect 9933 6817 9945 6820
rect 9979 6817 9991 6851
rect 9933 6811 9991 6817
rect 10410 6808 10416 6860
rect 10468 6848 10474 6860
rect 11054 6848 11060 6860
rect 10468 6820 11060 6848
rect 10468 6808 10474 6820
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 11204 6820 12112 6848
rect 11204 6808 11210 6820
rect 6328 6752 7236 6780
rect 8128 6752 8331 6780
rect 6328 6740 6334 6752
rect 3513 6715 3571 6721
rect 3513 6681 3525 6715
rect 3559 6712 3571 6715
rect 8128 6712 8156 6752
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8444 6752 9137 6780
rect 8444 6740 8450 6752
rect 9125 6749 9137 6752
rect 9171 6780 9183 6783
rect 9214 6780 9220 6792
rect 9171 6752 9220 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9548 6752 9689 6780
rect 9548 6740 9554 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 12084 6789 12112 6820
rect 12250 6808 12256 6860
rect 12308 6848 12314 6860
rect 12544 6848 12572 6888
rect 12802 6876 12808 6888
rect 12860 6876 12866 6928
rect 13081 6919 13139 6925
rect 13081 6885 13093 6919
rect 13127 6916 13139 6919
rect 15286 6916 15292 6928
rect 13127 6888 15292 6916
rect 13127 6885 13139 6888
rect 13081 6879 13139 6885
rect 15286 6876 15292 6888
rect 15344 6916 15350 6928
rect 16298 6916 16304 6928
rect 15344 6888 16304 6916
rect 15344 6876 15350 6888
rect 16298 6876 16304 6888
rect 16356 6876 16362 6928
rect 12308 6820 12572 6848
rect 12308 6808 12314 6820
rect 12618 6808 12624 6860
rect 12676 6848 12682 6860
rect 14274 6848 14280 6860
rect 12676 6820 13308 6848
rect 14235 6820 14280 6848
rect 12676 6808 12682 6820
rect 13004 6792 13032 6820
rect 11977 6783 12035 6789
rect 10744 6752 11836 6780
rect 10744 6740 10750 6752
rect 3559 6684 5304 6712
rect 3559 6681 3571 6684
rect 3513 6675 3571 6681
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 2498 6644 2504 6656
rect 1627 6616 2504 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 4065 6647 4123 6653
rect 4065 6613 4077 6647
rect 4111 6644 4123 6647
rect 4522 6644 4528 6656
rect 4111 6616 4528 6644
rect 4111 6613 4123 6616
rect 4065 6607 4123 6613
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 5276 6644 5304 6684
rect 6564 6684 7144 6712
rect 6564 6644 6592 6684
rect 5276 6616 6592 6644
rect 6641 6647 6699 6653
rect 6641 6613 6653 6647
rect 6687 6644 6699 6647
rect 6730 6644 6736 6656
rect 6687 6616 6736 6644
rect 6687 6613 6699 6616
rect 6641 6607 6699 6613
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 7116 6644 7144 6684
rect 8027 6684 8156 6712
rect 8573 6715 8631 6721
rect 8027 6644 8055 6684
rect 8573 6681 8585 6715
rect 8619 6712 8631 6715
rect 11698 6712 11704 6724
rect 8619 6684 9727 6712
rect 8619 6681 8631 6684
rect 8573 6675 8631 6681
rect 7116 6616 8055 6644
rect 8481 6647 8539 6653
rect 8481 6613 8493 6647
rect 8527 6644 8539 6647
rect 9582 6644 9588 6656
rect 8527 6616 9588 6644
rect 8527 6613 8539 6616
rect 8481 6607 8539 6613
rect 9582 6604 9588 6616
rect 9640 6604 9646 6656
rect 9699 6644 9727 6684
rect 11348 6684 11704 6712
rect 11348 6644 11376 6684
rect 11698 6672 11704 6684
rect 11756 6672 11762 6724
rect 9699 6616 11376 6644
rect 11422 6604 11428 6656
rect 11480 6644 11486 6656
rect 11517 6647 11575 6653
rect 11517 6644 11529 6647
rect 11480 6616 11529 6644
rect 11480 6604 11486 6616
rect 11517 6613 11529 6616
rect 11563 6613 11575 6647
rect 11808 6644 11836 6752
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 11992 6712 12020 6743
rect 12158 6740 12164 6792
rect 12216 6780 12222 6792
rect 12216 6752 12940 6780
rect 12216 6740 12222 6752
rect 12713 6715 12771 6721
rect 12713 6712 12725 6715
rect 11992 6684 12725 6712
rect 12713 6681 12725 6684
rect 12759 6681 12771 6715
rect 12912 6712 12940 6752
rect 12986 6740 12992 6792
rect 13044 6740 13050 6792
rect 13170 6780 13176 6792
rect 13083 6752 13176 6780
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 13280 6789 13308 6820
rect 14274 6808 14280 6820
rect 14332 6808 14338 6860
rect 13265 6783 13323 6789
rect 13265 6749 13277 6783
rect 13311 6749 13323 6783
rect 14366 6780 14372 6792
rect 14327 6752 14372 6780
rect 13265 6743 13323 6749
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 13188 6712 13216 6740
rect 12912 6684 13216 6712
rect 12713 6675 12771 6681
rect 13814 6672 13820 6724
rect 13872 6712 13878 6724
rect 13909 6715 13967 6721
rect 13909 6712 13921 6715
rect 13872 6684 13921 6712
rect 13872 6672 13878 6684
rect 13909 6681 13921 6684
rect 13955 6681 13967 6715
rect 14476 6712 14504 6743
rect 13909 6675 13967 6681
rect 14384 6684 14504 6712
rect 12250 6644 12256 6656
rect 11808 6616 12256 6644
rect 11517 6607 11575 6613
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12526 6604 12532 6656
rect 12584 6644 12590 6656
rect 14384 6644 14412 6684
rect 12584 6616 14412 6644
rect 12584 6604 12590 6616
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 2777 6443 2835 6449
rect 2188 6412 2452 6440
rect 2188 6400 2194 6412
rect 2424 6384 2452 6412
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 3786 6440 3792 6452
rect 2823 6412 3792 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 6917 6443 6975 6449
rect 6917 6440 6929 6443
rect 4120 6412 6929 6440
rect 4120 6400 4126 6412
rect 6917 6409 6929 6412
rect 6963 6409 6975 6443
rect 9582 6440 9588 6452
rect 6917 6403 6975 6409
rect 7484 6412 9588 6440
rect 2406 6332 2412 6384
rect 2464 6372 2470 6384
rect 6273 6375 6331 6381
rect 6273 6372 6285 6375
rect 2464 6344 2912 6372
rect 2464 6332 2470 6344
rect 1854 6264 1860 6316
rect 1912 6304 1918 6316
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 1912 6276 2145 6304
rect 1912 6264 1918 6276
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 2884 6304 2912 6344
rect 6012 6344 6285 6372
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2884 6276 3065 6304
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6236 2007 6239
rect 2406 6236 2412 6248
rect 1995 6208 2412 6236
rect 1995 6205 2007 6208
rect 1949 6199 2007 6205
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 2884 6168 2912 6276
rect 3053 6273 3065 6276
rect 3099 6273 3111 6307
rect 4890 6304 4896 6316
rect 4851 6276 4896 6304
rect 3053 6267 3111 6273
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6236 3019 6239
rect 4154 6236 4160 6248
rect 3007 6208 4160 6236
rect 3007 6205 3019 6208
rect 2961 6199 3019 6205
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 5160 6239 5218 6245
rect 5160 6205 5172 6239
rect 5206 6236 5218 6239
rect 5442 6236 5448 6248
rect 5206 6208 5448 6236
rect 5206 6205 5218 6208
rect 5160 6199 5218 6205
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 6012 6236 6040 6344
rect 6273 6341 6285 6344
rect 6319 6341 6331 6375
rect 6273 6335 6331 6341
rect 7484 6316 7512 6412
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 10226 6440 10232 6452
rect 9692 6412 10232 6440
rect 7650 6332 7656 6384
rect 7708 6332 7714 6384
rect 9122 6332 9128 6384
rect 9180 6372 9186 6384
rect 9306 6372 9312 6384
rect 9180 6344 9312 6372
rect 9180 6332 9186 6344
rect 9306 6332 9312 6344
rect 9364 6332 9370 6384
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 7466 6304 7472 6316
rect 6604 6276 7328 6304
rect 7379 6276 7472 6304
rect 6604 6264 6610 6276
rect 5684 6208 6040 6236
rect 5684 6196 5690 6208
rect 6086 6196 6092 6248
rect 6144 6236 6150 6248
rect 7190 6236 7196 6248
rect 6144 6208 7196 6236
rect 6144 6196 6150 6208
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 7300 6236 7328 6276
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 7668 6304 7696 6332
rect 8018 6304 8024 6316
rect 7668 6276 8024 6304
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 9398 6304 9404 6316
rect 9088 6276 9404 6304
rect 9088 6264 9094 6276
rect 9398 6264 9404 6276
rect 9456 6264 9462 6316
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6304 9551 6307
rect 9692 6304 9720 6412
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 10502 6440 10508 6452
rect 10463 6412 10508 6440
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 11146 6400 11152 6452
rect 11204 6440 11210 6452
rect 12250 6440 12256 6452
rect 11204 6412 12256 6440
rect 11204 6400 11210 6412
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 12492 6412 12537 6440
rect 12492 6400 12498 6412
rect 13170 6400 13176 6452
rect 13228 6440 13234 6452
rect 13633 6443 13691 6449
rect 13633 6440 13645 6443
rect 13228 6412 13645 6440
rect 13228 6400 13234 6412
rect 13633 6409 13645 6412
rect 13679 6409 13691 6443
rect 13633 6403 13691 6409
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 15010 6372 15016 6384
rect 9824 6344 14228 6372
rect 14971 6344 15016 6372
rect 9824 6332 9830 6344
rect 9539 6276 9720 6304
rect 9861 6307 9919 6313
rect 9539 6273 9551 6276
rect 9493 6267 9551 6273
rect 9861 6273 9873 6307
rect 9907 6304 9919 6307
rect 10686 6304 10692 6316
rect 9907 6276 10692 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10778 6264 10784 6316
rect 10836 6304 10842 6316
rect 11057 6307 11115 6313
rect 11057 6304 11069 6307
rect 10836 6276 11069 6304
rect 10836 6264 10842 6276
rect 11057 6273 11069 6276
rect 11103 6273 11115 6307
rect 12526 6304 12532 6316
rect 11057 6267 11115 6273
rect 11348 6276 12532 6304
rect 7377 6239 7435 6245
rect 7377 6236 7389 6239
rect 7300 6208 7389 6236
rect 7377 6205 7389 6208
rect 7423 6205 7435 6239
rect 7377 6199 7435 6205
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 7834 6236 7840 6248
rect 7708 6208 7840 6236
rect 7708 6196 7714 6208
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 11348 6236 11376 6276
rect 12526 6264 12532 6276
rect 12584 6264 12590 6316
rect 12986 6264 12992 6316
rect 13044 6304 13050 6316
rect 14200 6313 14228 6344
rect 15010 6332 15016 6344
rect 15068 6332 15074 6384
rect 14185 6307 14243 6313
rect 13044 6276 13089 6304
rect 13044 6264 13050 6276
rect 14185 6273 14197 6307
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 8128 6208 11376 6236
rect 3142 6168 3148 6180
rect 2884 6140 3148 6168
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 3320 6171 3378 6177
rect 3320 6137 3332 6171
rect 3366 6168 3378 6171
rect 3418 6168 3424 6180
rect 3366 6140 3424 6168
rect 3366 6137 3378 6140
rect 3320 6131 3378 6137
rect 3418 6128 3424 6140
rect 3476 6128 3482 6180
rect 5534 6168 5540 6180
rect 4448 6140 5540 6168
rect 1486 6060 1492 6112
rect 1544 6100 1550 6112
rect 1581 6103 1639 6109
rect 1581 6100 1593 6103
rect 1544 6072 1593 6100
rect 1544 6060 1550 6072
rect 1581 6069 1593 6072
rect 1627 6069 1639 6103
rect 1581 6063 1639 6069
rect 2041 6103 2099 6109
rect 2041 6069 2053 6103
rect 2087 6100 2099 6103
rect 4062 6100 4068 6112
rect 2087 6072 4068 6100
rect 2087 6069 2099 6072
rect 2041 6063 2099 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4448 6109 4476 6140
rect 5534 6128 5540 6140
rect 5592 6128 5598 6180
rect 5810 6128 5816 6180
rect 5868 6168 5874 6180
rect 6914 6168 6920 6180
rect 5868 6140 6920 6168
rect 5868 6128 5874 6140
rect 6914 6128 6920 6140
rect 6972 6128 6978 6180
rect 8128 6168 8156 6208
rect 8294 6177 8300 6180
rect 8288 6168 8300 6177
rect 7208 6140 8156 6168
rect 8255 6140 8300 6168
rect 4433 6103 4491 6109
rect 4433 6069 4445 6103
rect 4479 6069 4491 6103
rect 4433 6063 4491 6069
rect 4890 6060 4896 6112
rect 4948 6100 4954 6112
rect 7208 6100 7236 6140
rect 8288 6131 8300 6140
rect 8294 6128 8300 6131
rect 8352 6128 8358 6180
rect 8386 6128 8392 6180
rect 8444 6168 8450 6180
rect 9950 6168 9956 6180
rect 8444 6140 9956 6168
rect 8444 6128 8450 6140
rect 9950 6128 9956 6140
rect 10008 6128 10014 6180
rect 10594 6128 10600 6180
rect 10652 6168 10658 6180
rect 10873 6171 10931 6177
rect 10873 6168 10885 6171
rect 10652 6140 10885 6168
rect 10652 6128 10658 6140
rect 10873 6137 10885 6140
rect 10919 6137 10931 6171
rect 10980 6168 11008 6208
rect 11422 6196 11428 6248
rect 11480 6236 11486 6248
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 11480 6208 14013 6236
rect 11480 6196 11486 6208
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 11146 6168 11152 6180
rect 10980 6140 11152 6168
rect 10873 6131 10931 6137
rect 11146 6128 11152 6140
rect 11204 6128 11210 6180
rect 12250 6128 12256 6180
rect 12308 6168 12314 6180
rect 14093 6171 14151 6177
rect 14093 6168 14105 6171
rect 12308 6140 14105 6168
rect 12308 6128 12314 6140
rect 14093 6137 14105 6140
rect 14139 6137 14151 6171
rect 14844 6168 14872 6199
rect 15194 6168 15200 6180
rect 14844 6140 15200 6168
rect 14093 6131 14151 6137
rect 15194 6128 15200 6140
rect 15252 6128 15258 6180
rect 4948 6072 7236 6100
rect 7285 6103 7343 6109
rect 4948 6060 4954 6072
rect 7285 6069 7297 6103
rect 7331 6100 7343 6103
rect 8110 6100 8116 6112
rect 7331 6072 8116 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 9401 6103 9459 6109
rect 9401 6100 9413 6103
rect 8260 6072 9413 6100
rect 8260 6060 8266 6072
rect 9401 6069 9413 6072
rect 9447 6100 9459 6103
rect 10134 6100 10140 6112
rect 9447 6072 10140 6100
rect 9447 6069 9459 6072
rect 9401 6063 9459 6069
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10502 6060 10508 6112
rect 10560 6100 10566 6112
rect 10965 6103 11023 6109
rect 10965 6100 10977 6103
rect 10560 6072 10977 6100
rect 10560 6060 10566 6072
rect 10965 6069 10977 6072
rect 11011 6069 11023 6103
rect 10965 6063 11023 6069
rect 11701 6103 11759 6109
rect 11701 6069 11713 6103
rect 11747 6100 11759 6103
rect 12434 6100 12440 6112
rect 11747 6072 12440 6100
rect 11747 6069 11759 6072
rect 11701 6063 11759 6069
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 12526 6060 12532 6112
rect 12584 6100 12590 6112
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 12584 6072 12817 6100
rect 12584 6060 12590 6072
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 12805 6063 12863 6069
rect 12897 6103 12955 6109
rect 12897 6069 12909 6103
rect 12943 6100 12955 6103
rect 14182 6100 14188 6112
rect 12943 6072 14188 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 1949 5899 2007 5905
rect 1949 5865 1961 5899
rect 1995 5896 2007 5899
rect 2590 5896 2596 5908
rect 1995 5868 2596 5896
rect 1995 5865 2007 5868
rect 1949 5859 2007 5865
rect 2590 5856 2596 5868
rect 2648 5856 2654 5908
rect 2682 5856 2688 5908
rect 2740 5896 2746 5908
rect 3513 5899 3571 5905
rect 3513 5896 3525 5899
rect 2740 5868 3525 5896
rect 2740 5856 2746 5868
rect 3513 5865 3525 5868
rect 3559 5865 3571 5899
rect 4890 5896 4896 5908
rect 3513 5859 3571 5865
rect 4632 5868 4896 5896
rect 4062 5828 4068 5840
rect 1412 5800 4068 5828
rect 1412 5769 1440 5800
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5729 1455 5763
rect 1762 5760 1768 5772
rect 1723 5732 1768 5760
rect 1397 5723 1455 5729
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 2130 5760 2136 5772
rect 2091 5732 2136 5760
rect 2130 5720 2136 5732
rect 2188 5720 2194 5772
rect 2400 5763 2458 5769
rect 2400 5729 2412 5763
rect 2446 5760 2458 5763
rect 4632 5760 4660 5868
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 7653 5899 7711 5905
rect 5184 5868 7604 5896
rect 4700 5831 4758 5837
rect 4700 5797 4712 5831
rect 4746 5828 4758 5831
rect 5184 5828 5212 5868
rect 4746 5800 5212 5828
rect 4746 5797 4758 5800
rect 4700 5791 4758 5797
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 5316 5800 6684 5828
rect 5316 5788 5322 5800
rect 2446 5732 4660 5760
rect 2446 5729 2458 5732
rect 2400 5723 2458 5729
rect 5166 5720 5172 5772
rect 5224 5760 5230 5772
rect 5224 5732 5488 5760
rect 5224 5720 5230 5732
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3326 5692 3332 5704
rect 3200 5664 3332 5692
rect 3200 5652 3206 5664
rect 3326 5652 3332 5664
rect 3384 5692 3390 5704
rect 4433 5695 4491 5701
rect 4433 5692 4445 5695
rect 3384 5664 4445 5692
rect 3384 5652 3390 5664
rect 4433 5661 4445 5664
rect 4479 5661 4491 5695
rect 5460 5692 5488 5732
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 6178 5760 6184 5772
rect 5592 5732 6184 5760
rect 5592 5720 5598 5732
rect 6178 5720 6184 5732
rect 6236 5760 6242 5772
rect 6529 5763 6587 5769
rect 6529 5760 6541 5763
rect 6236 5732 6541 5760
rect 6236 5720 6242 5732
rect 6529 5729 6541 5732
rect 6575 5729 6587 5763
rect 6656 5760 6684 5800
rect 6914 5788 6920 5840
rect 6972 5828 6978 5840
rect 7282 5828 7288 5840
rect 6972 5800 7288 5828
rect 6972 5788 6978 5800
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 7576 5828 7604 5868
rect 7653 5865 7665 5899
rect 7699 5896 7711 5899
rect 8386 5896 8392 5908
rect 7699 5868 8392 5896
rect 7699 5865 7711 5868
rect 7653 5859 7711 5865
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 8757 5899 8815 5905
rect 8757 5896 8769 5899
rect 8628 5868 8769 5896
rect 8628 5856 8634 5868
rect 8757 5865 8769 5868
rect 8803 5865 8815 5899
rect 8757 5859 8815 5865
rect 8849 5899 8907 5905
rect 8849 5865 8861 5899
rect 8895 5896 8907 5899
rect 12713 5899 12771 5905
rect 8895 5868 11560 5896
rect 8895 5865 8907 5868
rect 8849 5859 8907 5865
rect 7834 5828 7840 5840
rect 7576 5800 7840 5828
rect 7834 5788 7840 5800
rect 7892 5788 7898 5840
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 8168 5800 10088 5828
rect 8168 5788 8174 5800
rect 8273 5763 8331 5769
rect 8273 5760 8285 5763
rect 6656 5732 8285 5760
rect 6529 5723 6587 5729
rect 8273 5729 8285 5732
rect 8319 5729 8331 5763
rect 8273 5723 8331 5729
rect 8386 5720 8392 5772
rect 8444 5760 8450 5772
rect 8570 5760 8576 5772
rect 8444 5732 8576 5760
rect 8444 5720 8450 5732
rect 8570 5720 8576 5732
rect 8628 5760 8634 5772
rect 8754 5760 8760 5772
rect 8628 5732 8760 5760
rect 8628 5720 8634 5732
rect 8754 5720 8760 5732
rect 8812 5720 8818 5772
rect 9030 5720 9036 5772
rect 9088 5760 9094 5772
rect 9766 5760 9772 5772
rect 9088 5732 9772 5760
rect 9088 5720 9094 5732
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 9950 5769 9956 5772
rect 9944 5760 9956 5769
rect 9911 5732 9956 5760
rect 9944 5723 9956 5732
rect 9950 5720 9956 5723
rect 10008 5720 10014 5772
rect 10060 5760 10088 5800
rect 10134 5788 10140 5840
rect 10192 5828 10198 5840
rect 11054 5828 11060 5840
rect 10192 5800 11060 5828
rect 10192 5788 10198 5800
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 11532 5760 11560 5868
rect 12713 5865 12725 5899
rect 12759 5896 12771 5899
rect 13630 5896 13636 5908
rect 12759 5868 13636 5896
rect 12759 5865 12771 5868
rect 12713 5859 12771 5865
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 13909 5899 13967 5905
rect 13909 5865 13921 5899
rect 13955 5896 13967 5899
rect 14274 5896 14280 5908
rect 13955 5868 14280 5896
rect 13955 5865 13967 5868
rect 13909 5859 13967 5865
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 15194 5896 15200 5908
rect 14415 5868 15200 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 11882 5788 11888 5840
rect 11940 5828 11946 5840
rect 12434 5828 12440 5840
rect 11940 5800 12440 5828
rect 11940 5788 11946 5800
rect 12434 5788 12440 5800
rect 12492 5788 12498 5840
rect 13814 5788 13820 5840
rect 13872 5828 13878 5840
rect 14384 5828 14412 5859
rect 15194 5856 15200 5868
rect 15252 5856 15258 5908
rect 13872 5800 14412 5828
rect 13872 5788 13878 5800
rect 11977 5763 12035 5769
rect 10060 5732 11100 5760
rect 11532 5732 11744 5760
rect 5994 5692 6000 5704
rect 5460 5664 6000 5692
rect 4433 5655 4491 5661
rect 5552 5636 5580 5664
rect 5994 5652 6000 5664
rect 6052 5692 6058 5704
rect 6273 5695 6331 5701
rect 6273 5692 6285 5695
rect 6052 5664 6285 5692
rect 6052 5652 6058 5664
rect 6273 5661 6285 5664
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 7926 5652 7932 5704
rect 7984 5692 7990 5704
rect 8938 5692 8944 5704
rect 7984 5664 8944 5692
rect 7984 5652 7990 5664
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 9490 5652 9496 5704
rect 9548 5692 9554 5704
rect 9677 5695 9735 5701
rect 9677 5692 9689 5695
rect 9548 5664 9689 5692
rect 9548 5652 9554 5664
rect 9677 5661 9689 5664
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 1581 5627 1639 5633
rect 1581 5593 1593 5627
rect 1627 5624 1639 5627
rect 1627 5596 2176 5624
rect 1627 5593 1639 5596
rect 1581 5587 1639 5593
rect 2148 5556 2176 5596
rect 3418 5584 3424 5636
rect 3476 5624 3482 5636
rect 4246 5624 4252 5636
rect 3476 5596 4252 5624
rect 3476 5584 3482 5596
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 5534 5584 5540 5636
rect 5592 5584 5598 5636
rect 8113 5627 8171 5633
rect 5644 5596 5939 5624
rect 3142 5556 3148 5568
rect 2148 5528 3148 5556
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 5074 5556 5080 5568
rect 3936 5528 5080 5556
rect 3936 5516 3942 5528
rect 5074 5516 5080 5528
rect 5132 5516 5138 5568
rect 5442 5516 5448 5568
rect 5500 5556 5506 5568
rect 5644 5556 5672 5596
rect 5810 5556 5816 5568
rect 5500 5528 5672 5556
rect 5771 5528 5816 5556
rect 5500 5516 5506 5528
rect 5810 5516 5816 5528
rect 5868 5516 5874 5568
rect 5911 5556 5939 5596
rect 7208 5596 7963 5624
rect 7208 5556 7236 5596
rect 5911 5528 7236 5556
rect 7282 5516 7288 5568
rect 7340 5556 7346 5568
rect 7834 5556 7840 5568
rect 7340 5528 7840 5556
rect 7340 5516 7346 5528
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 7935 5556 7963 5596
rect 8113 5593 8125 5627
rect 8159 5624 8171 5627
rect 8389 5627 8447 5633
rect 8159 5596 8340 5624
rect 8159 5593 8171 5596
rect 8113 5587 8171 5593
rect 8202 5556 8208 5568
rect 7935 5528 8208 5556
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 8312 5556 8340 5596
rect 8389 5593 8401 5627
rect 8435 5624 8447 5627
rect 11072 5624 11100 5732
rect 11517 5627 11575 5633
rect 11517 5624 11529 5627
rect 8435 5596 9727 5624
rect 11072 5596 11529 5624
rect 8435 5593 8447 5596
rect 8389 5587 8447 5593
rect 9030 5556 9036 5568
rect 8312 5528 9036 5556
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 9699 5556 9727 5596
rect 11517 5593 11529 5596
rect 11563 5593 11575 5627
rect 11716 5624 11744 5732
rect 11977 5729 11989 5763
rect 12023 5760 12035 5763
rect 12618 5760 12624 5772
rect 12023 5732 12624 5760
rect 12023 5729 12035 5732
rect 11977 5723 12035 5729
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 13081 5763 13139 5769
rect 13081 5729 13093 5763
rect 13127 5760 13139 5763
rect 13630 5760 13636 5772
rect 13127 5732 13636 5760
rect 13127 5729 13139 5732
rect 13081 5723 13139 5729
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 14182 5720 14188 5772
rect 14240 5760 14246 5772
rect 14277 5763 14335 5769
rect 14277 5760 14289 5763
rect 14240 5732 14289 5760
rect 14240 5720 14246 5732
rect 14277 5729 14289 5732
rect 14323 5729 14335 5763
rect 14277 5723 14335 5729
rect 11882 5652 11888 5704
rect 11940 5692 11946 5704
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 11940 5664 12081 5692
rect 11940 5652 11946 5664
rect 12069 5661 12081 5664
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 12710 5652 12716 5704
rect 12768 5692 12774 5704
rect 13173 5695 13231 5701
rect 13173 5692 13185 5695
rect 12768 5664 13185 5692
rect 12768 5652 12774 5664
rect 13173 5661 13185 5664
rect 13219 5661 13231 5695
rect 13173 5655 13231 5661
rect 13357 5695 13415 5701
rect 13357 5661 13369 5695
rect 13403 5692 13415 5695
rect 13722 5692 13728 5704
rect 13403 5664 13728 5692
rect 13403 5661 13415 5664
rect 13357 5655 13415 5661
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 14458 5652 14464 5704
rect 14516 5692 14522 5704
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 14516 5664 14565 5692
rect 14516 5652 14522 5664
rect 14553 5661 14565 5664
rect 14599 5692 14611 5695
rect 14826 5692 14832 5704
rect 14599 5664 14832 5692
rect 14599 5661 14611 5664
rect 14553 5655 14611 5661
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 12250 5624 12256 5636
rect 11716 5596 12256 5624
rect 11517 5587 11575 5593
rect 12250 5584 12256 5596
rect 12308 5624 12314 5636
rect 14918 5624 14924 5636
rect 12308 5596 14924 5624
rect 12308 5584 12314 5596
rect 14918 5584 14924 5596
rect 14976 5584 14982 5636
rect 10962 5556 10968 5568
rect 9699 5528 10968 5556
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 11057 5559 11115 5565
rect 11057 5525 11069 5559
rect 11103 5556 11115 5559
rect 11146 5556 11152 5568
rect 11103 5528 11152 5556
rect 11103 5525 11115 5528
rect 11057 5519 11115 5525
rect 11146 5516 11152 5528
rect 11204 5516 11210 5568
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 2774 5352 2780 5364
rect 2240 5324 2780 5352
rect 1946 5176 1952 5228
rect 2004 5176 2010 5228
rect 2240 5225 2268 5324
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 3326 5352 3332 5364
rect 3068 5324 3332 5352
rect 2866 5244 2872 5296
rect 2924 5244 2930 5296
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 2884 5216 2912 5244
rect 3068 5225 3096 5324
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 6730 5352 6736 5364
rect 4120 5324 6736 5352
rect 4120 5312 4126 5324
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 6825 5355 6883 5361
rect 6825 5321 6837 5355
rect 6871 5352 6883 5355
rect 6914 5352 6920 5364
rect 6871 5324 6920 5352
rect 6871 5321 6883 5324
rect 6825 5315 6883 5321
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 9217 5355 9275 5361
rect 9217 5352 9229 5355
rect 7248 5324 9229 5352
rect 7248 5312 7254 5324
rect 6270 5244 6276 5296
rect 6328 5284 6334 5296
rect 6638 5284 6644 5296
rect 6328 5256 6644 5284
rect 6328 5244 6334 5256
rect 6638 5244 6644 5256
rect 6696 5244 6702 5296
rect 2731 5188 2912 5216
rect 3053 5219 3111 5225
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 3053 5185 3065 5219
rect 3099 5185 3111 5219
rect 6457 5219 6515 5225
rect 3053 5179 3111 5185
rect 4080 5188 5028 5216
rect 1964 5148 1992 5176
rect 2409 5151 2467 5157
rect 2409 5148 2421 5151
rect 1964 5120 2421 5148
rect 2409 5117 2421 5120
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 3320 5151 3378 5157
rect 3320 5117 3332 5151
rect 3366 5148 3378 5151
rect 4080 5148 4108 5188
rect 4893 5151 4951 5157
rect 4893 5148 4905 5151
rect 3366 5120 4108 5148
rect 4172 5120 4905 5148
rect 3366 5117 3378 5120
rect 3320 5111 3378 5117
rect 1949 5083 2007 5089
rect 1949 5049 1961 5083
rect 1995 5080 2007 5083
rect 2130 5080 2136 5092
rect 1995 5052 2136 5080
rect 1995 5049 2007 5052
rect 1949 5043 2007 5049
rect 2130 5040 2136 5052
rect 2188 5040 2194 5092
rect 3970 5040 3976 5092
rect 4028 5080 4034 5092
rect 4172 5080 4200 5120
rect 4893 5117 4905 5120
rect 4939 5117 4951 5151
rect 5000 5148 5028 5188
rect 6457 5185 6469 5219
rect 6503 5216 6515 5219
rect 7006 5216 7012 5228
rect 6503 5188 7012 5216
rect 6503 5185 6515 5188
rect 6457 5179 6515 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 7190 5176 7196 5228
rect 7248 5216 7254 5228
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 7248 5188 7389 5216
rect 7248 5176 7254 5188
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 5902 5148 5908 5160
rect 5000 5120 5908 5148
rect 4893 5111 4951 5117
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 7837 5151 7895 5157
rect 7837 5148 7849 5151
rect 6052 5120 7849 5148
rect 6052 5108 6058 5120
rect 7837 5117 7849 5120
rect 7883 5117 7895 5151
rect 8864 5148 8892 5324
rect 9217 5321 9229 5324
rect 9263 5321 9275 5355
rect 9217 5315 9275 5321
rect 9582 5312 9588 5364
rect 9640 5312 9646 5364
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 10505 5355 10563 5361
rect 10505 5352 10517 5355
rect 9732 5324 10517 5352
rect 9732 5312 9738 5324
rect 10505 5321 10517 5324
rect 10551 5321 10563 5355
rect 10505 5315 10563 5321
rect 10870 5312 10876 5364
rect 10928 5352 10934 5364
rect 11882 5352 11888 5364
rect 10928 5324 11888 5352
rect 10928 5312 10934 5324
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 14458 5352 14464 5364
rect 12483 5324 14464 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 9309 5287 9367 5293
rect 9309 5253 9321 5287
rect 9355 5253 9367 5287
rect 9600 5284 9628 5312
rect 9600 5256 11100 5284
rect 9309 5247 9367 5253
rect 9324 5216 9352 5247
rect 9950 5216 9956 5228
rect 9324 5188 9727 5216
rect 9911 5188 9956 5216
rect 9214 5148 9220 5160
rect 8864 5120 9220 5148
rect 7837 5111 7895 5117
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 5138 5083 5196 5089
rect 5138 5080 5150 5083
rect 4028 5052 4200 5080
rect 4908 5052 5150 5080
rect 4028 5040 4034 5052
rect 4908 5024 4936 5052
rect 5138 5049 5150 5052
rect 5184 5049 5196 5083
rect 5138 5043 5196 5049
rect 6178 5040 6184 5092
rect 6236 5080 6242 5092
rect 6730 5080 6736 5092
rect 6236 5052 6736 5080
rect 6236 5040 6242 5052
rect 6730 5040 6736 5052
rect 6788 5040 6794 5092
rect 7006 5040 7012 5092
rect 7064 5080 7070 5092
rect 8082 5083 8140 5089
rect 8082 5080 8094 5083
rect 7064 5052 8094 5080
rect 7064 5040 7070 5052
rect 8082 5049 8094 5052
rect 8128 5080 8140 5083
rect 8202 5080 8208 5092
rect 8128 5052 8208 5080
rect 8128 5049 8140 5052
rect 8082 5043 8140 5049
rect 8202 5040 8208 5052
rect 8260 5040 8266 5092
rect 9699 5080 9727 5188
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 10318 5216 10324 5228
rect 10060 5188 10324 5216
rect 9769 5151 9827 5157
rect 9769 5117 9781 5151
rect 9815 5148 9827 5151
rect 10060 5148 10088 5188
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 10962 5216 10968 5228
rect 10923 5188 10968 5216
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 11072 5225 11100 5256
rect 11422 5244 11428 5296
rect 11480 5284 11486 5296
rect 13722 5284 13728 5296
rect 11480 5256 13728 5284
rect 11480 5244 11486 5256
rect 11057 5219 11115 5225
rect 11057 5185 11069 5219
rect 11103 5185 11115 5219
rect 11057 5179 11115 5185
rect 11698 5176 11704 5228
rect 11756 5216 11762 5228
rect 13096 5225 13124 5256
rect 13722 5244 13728 5256
rect 13780 5284 13786 5296
rect 13780 5256 14228 5284
rect 13780 5244 13786 5256
rect 13081 5219 13139 5225
rect 11756 5188 12388 5216
rect 11756 5176 11762 5188
rect 9815 5120 10088 5148
rect 10137 5151 10195 5157
rect 9815 5117 9827 5120
rect 9769 5111 9827 5117
rect 10137 5117 10149 5151
rect 10183 5148 10195 5151
rect 12360 5148 12388 5188
rect 13081 5185 13093 5219
rect 13127 5185 13139 5219
rect 14090 5216 14096 5228
rect 14051 5188 14096 5216
rect 13081 5179 13139 5185
rect 14090 5176 14096 5188
rect 14148 5176 14154 5228
rect 14200 5225 14228 5256
rect 14185 5219 14243 5225
rect 14185 5185 14197 5219
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 14001 5151 14059 5157
rect 14001 5148 14013 5151
rect 10183 5120 11928 5148
rect 12360 5120 14013 5148
rect 10183 5117 10195 5120
rect 10137 5111 10195 5117
rect 10873 5083 10931 5089
rect 10873 5080 10885 5083
rect 9699 5052 10885 5080
rect 10873 5049 10885 5052
rect 10919 5049 10931 5083
rect 11790 5080 11796 5092
rect 10873 5043 10931 5049
rect 10980 5052 11796 5080
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 2041 5015 2099 5021
rect 2041 4981 2053 5015
rect 2087 5012 2099 5015
rect 4062 5012 4068 5024
rect 2087 4984 4068 5012
rect 2087 4981 2099 4984
rect 2041 4975 2099 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 4433 5015 4491 5021
rect 4433 5012 4445 5015
rect 4304 4984 4445 5012
rect 4304 4972 4310 4984
rect 4433 4981 4445 4984
rect 4479 4981 4491 5015
rect 4433 4975 4491 4981
rect 4890 4972 4896 5024
rect 4948 4972 4954 5024
rect 6270 5012 6276 5024
rect 6231 4984 6276 5012
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 6972 4984 7205 5012
rect 6972 4972 6978 4984
rect 7193 4981 7205 4984
rect 7239 4981 7251 5015
rect 7193 4975 7251 4981
rect 7285 5015 7343 5021
rect 7285 4981 7297 5015
rect 7331 5012 7343 5015
rect 9490 5012 9496 5024
rect 7331 4984 9496 5012
rect 7331 4981 7343 4984
rect 7285 4975 7343 4981
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 9677 5015 9735 5021
rect 9677 4981 9689 5015
rect 9723 5012 9735 5015
rect 10980 5012 11008 5052
rect 11790 5040 11796 5052
rect 11848 5040 11854 5092
rect 11698 5012 11704 5024
rect 9723 4984 11008 5012
rect 11659 4984 11704 5012
rect 9723 4981 9735 4984
rect 9677 4975 9735 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 11900 5012 11928 5120
rect 14001 5117 14013 5120
rect 14047 5117 14059 5151
rect 14829 5151 14887 5157
rect 14829 5148 14841 5151
rect 14001 5111 14059 5117
rect 14108 5120 14841 5148
rect 14108 5092 14136 5120
rect 14829 5117 14841 5120
rect 14875 5117 14887 5151
rect 14829 5111 14887 5117
rect 12066 5040 12072 5092
rect 12124 5080 12130 5092
rect 12805 5083 12863 5089
rect 12805 5080 12817 5083
rect 12124 5052 12817 5080
rect 12124 5040 12130 5052
rect 12805 5049 12817 5052
rect 12851 5049 12863 5083
rect 12805 5043 12863 5049
rect 14090 5040 14096 5092
rect 14148 5040 14154 5092
rect 12526 5012 12532 5024
rect 11900 4984 12532 5012
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 12894 5012 12900 5024
rect 12855 4984 12900 5012
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 13633 5015 13691 5021
rect 13633 4981 13645 5015
rect 13679 5012 13691 5015
rect 14274 5012 14280 5024
rect 13679 4984 14280 5012
rect 13679 4981 13691 4984
rect 13633 4975 13691 4981
rect 14274 4972 14280 4984
rect 14332 4972 14338 5024
rect 15010 5012 15016 5024
rect 14971 4984 15016 5012
rect 15010 4972 15016 4984
rect 15068 4972 15074 5024
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 1578 4768 1584 4820
rect 1636 4808 1642 4820
rect 3329 4811 3387 4817
rect 3329 4808 3341 4811
rect 1636 4780 3341 4808
rect 1636 4768 1642 4780
rect 3329 4777 3341 4780
rect 3375 4777 3387 4811
rect 3329 4771 3387 4777
rect 3418 4768 3424 4820
rect 3476 4808 3482 4820
rect 4798 4808 4804 4820
rect 3476 4780 4804 4808
rect 3476 4768 3482 4780
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 5442 4808 5448 4820
rect 5403 4780 5448 4808
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 5592 4780 5939 4808
rect 5592 4768 5598 4780
rect 3237 4743 3295 4749
rect 3237 4709 3249 4743
rect 3283 4740 3295 4743
rect 5911 4740 5939 4780
rect 6270 4768 6276 4820
rect 6328 4808 6334 4820
rect 6328 4780 6875 4808
rect 6328 4768 6334 4780
rect 5994 4740 6000 4752
rect 3283 4712 5847 4740
rect 3283 4709 3295 4712
rect 3237 4703 3295 4709
rect 1664 4675 1722 4681
rect 1664 4641 1676 4675
rect 1710 4672 1722 4675
rect 3418 4672 3424 4684
rect 1710 4644 3424 4672
rect 1710 4641 1722 4644
rect 1664 4635 1722 4641
rect 3418 4632 3424 4644
rect 3476 4632 3482 4684
rect 4332 4675 4390 4681
rect 4332 4672 4344 4675
rect 3528 4644 4344 4672
rect 3528 4613 3556 4644
rect 4332 4641 4344 4644
rect 4378 4672 4390 4675
rect 5534 4672 5540 4684
rect 4378 4644 5540 4672
rect 4378 4641 4390 4644
rect 4332 4635 4390 4641
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 3970 4564 3976 4616
rect 4028 4604 4034 4616
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 4028 4576 4077 4604
rect 4028 4564 4034 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 5819 4604 5847 4712
rect 5911 4712 6000 4740
rect 5911 4681 5939 4712
rect 5994 4700 6000 4712
rect 6052 4700 6058 4752
rect 6730 4740 6736 4752
rect 6104 4712 6736 4740
rect 5905 4675 5963 4681
rect 5905 4641 5917 4675
rect 5951 4641 5963 4675
rect 6104 4672 6132 4712
rect 6730 4700 6736 4712
rect 6788 4700 6794 4752
rect 6847 4740 6875 4780
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 10873 4811 10931 4817
rect 10873 4808 10885 4811
rect 6972 4780 10885 4808
rect 6972 4768 6978 4780
rect 10873 4777 10885 4780
rect 10919 4777 10931 4811
rect 11238 4808 11244 4820
rect 11199 4780 11244 4808
rect 10873 4771 10931 4777
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 12250 4768 12256 4820
rect 12308 4808 12314 4820
rect 12434 4808 12440 4820
rect 12308 4780 12440 4808
rect 12308 4768 12314 4780
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 13078 4768 13084 4820
rect 13136 4808 13142 4820
rect 13722 4808 13728 4820
rect 13136 4780 13728 4808
rect 13136 4768 13142 4780
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 10137 4743 10195 4749
rect 6847 4712 9904 4740
rect 5905 4635 5963 4641
rect 6012 4644 6132 4672
rect 6172 4675 6230 4681
rect 6012 4604 6040 4644
rect 6172 4641 6184 4675
rect 6218 4672 6230 4675
rect 6546 4672 6552 4684
rect 6218 4644 6552 4672
rect 6218 4641 6230 4644
rect 6172 4635 6230 4641
rect 6546 4632 6552 4644
rect 6604 4672 6610 4684
rect 7190 4672 7196 4684
rect 6604 4644 7196 4672
rect 6604 4632 6610 4644
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 7282 4632 7288 4684
rect 7340 4672 7346 4684
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 7340 4644 7389 4672
rect 7340 4632 7346 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 8012 4675 8070 4681
rect 8012 4672 8024 4675
rect 7377 4635 7435 4641
rect 7668 4644 8024 4672
rect 5819 4576 6040 4604
rect 4065 4567 4123 4573
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7466 4604 7472 4616
rect 6972 4576 7472 4604
rect 6972 4564 6978 4576
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 2777 4539 2835 4545
rect 2777 4505 2789 4539
rect 2823 4536 2835 4539
rect 3786 4536 3792 4548
rect 2823 4508 3792 4536
rect 2823 4505 2835 4508
rect 2777 4499 2835 4505
rect 3786 4496 3792 4508
rect 3844 4496 3850 4548
rect 5166 4496 5172 4548
rect 5224 4536 5230 4548
rect 7561 4539 7619 4545
rect 7561 4536 7573 4539
rect 5224 4508 5580 4536
rect 5224 4496 5230 4508
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 3878 4468 3884 4480
rect 2915 4440 3884 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 5552 4468 5580 4508
rect 6840 4508 7573 4536
rect 6840 4468 6868 4508
rect 7561 4505 7573 4508
rect 7607 4505 7619 4539
rect 7561 4499 7619 4505
rect 5552 4440 6868 4468
rect 7285 4471 7343 4477
rect 7285 4437 7297 4471
rect 7331 4468 7343 4471
rect 7668 4468 7696 4644
rect 8012 4641 8024 4644
rect 8058 4672 8070 4675
rect 9674 4672 9680 4684
rect 8058 4644 9680 4672
rect 8058 4641 8070 4644
rect 8012 4635 8070 4641
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 7331 4440 7696 4468
rect 7760 4468 7788 4567
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 9766 4604 9772 4616
rect 8812 4576 9772 4604
rect 8812 4564 8818 4576
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 9876 4604 9904 4712
rect 10137 4709 10149 4743
rect 10183 4740 10195 4743
rect 10410 4740 10416 4752
rect 10183 4712 10416 4740
rect 10183 4709 10195 4712
rect 10137 4703 10195 4709
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 10962 4700 10968 4752
rect 11020 4740 11026 4752
rect 11790 4740 11796 4752
rect 11020 4712 11796 4740
rect 11020 4700 11026 4712
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 11882 4700 11888 4752
rect 11940 4740 11946 4752
rect 13633 4743 13691 4749
rect 13633 4740 13645 4743
rect 11940 4712 13645 4740
rect 11940 4700 11946 4712
rect 13633 4709 13645 4712
rect 13679 4709 13691 4743
rect 13633 4703 13691 4709
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10318 4672 10324 4684
rect 10091 4644 10324 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10318 4632 10324 4644
rect 10376 4672 10382 4684
rect 11146 4672 11152 4684
rect 10376 4644 11152 4672
rect 10376 4632 10382 4644
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4672 11391 4675
rect 13998 4672 14004 4684
rect 11379 4644 14004 4672
rect 11379 4641 11391 4644
rect 11333 4635 11391 4641
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 14461 4675 14519 4681
rect 14461 4641 14473 4675
rect 14507 4672 14519 4675
rect 14550 4672 14556 4684
rect 14507 4644 14556 4672
rect 14507 4641 14519 4644
rect 14461 4635 14519 4641
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 9876 4576 10241 4604
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 11238 4564 11244 4616
rect 11296 4604 11302 4616
rect 11425 4607 11483 4613
rect 11425 4604 11437 4607
rect 11296 4576 11437 4604
rect 11296 4564 11302 4576
rect 11425 4573 11437 4576
rect 11471 4573 11483 4607
rect 12526 4604 12532 4616
rect 12487 4576 12532 4604
rect 11425 4567 11483 4573
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 12621 4607 12679 4613
rect 12621 4573 12633 4607
rect 12667 4604 12679 4607
rect 13817 4607 13875 4613
rect 13817 4604 13829 4607
rect 12667 4576 13829 4604
rect 12667 4573 12679 4576
rect 12621 4567 12679 4573
rect 13817 4573 13829 4576
rect 13863 4573 13875 4607
rect 13817 4567 13875 4573
rect 8938 4496 8944 4548
rect 8996 4536 9002 4548
rect 9125 4539 9183 4545
rect 9125 4536 9137 4539
rect 8996 4508 9137 4536
rect 8996 4496 9002 4508
rect 9125 4505 9137 4508
rect 9171 4536 9183 4539
rect 9950 4536 9956 4548
rect 9171 4508 9956 4536
rect 9171 4505 9183 4508
rect 9125 4499 9183 4505
rect 9950 4496 9956 4508
rect 10008 4496 10014 4548
rect 10870 4496 10876 4548
rect 10928 4536 10934 4548
rect 10928 4508 12204 4536
rect 10928 4496 10934 4508
rect 7926 4468 7932 4480
rect 7760 4440 7932 4468
rect 7331 4437 7343 4440
rect 7285 4431 7343 4437
rect 7926 4428 7932 4440
rect 7984 4428 7990 4480
rect 8110 4428 8116 4480
rect 8168 4468 8174 4480
rect 8754 4468 8760 4480
rect 8168 4440 8760 4468
rect 8168 4428 8174 4440
rect 8754 4428 8760 4440
rect 8812 4428 8818 4480
rect 9674 4468 9680 4480
rect 9635 4440 9680 4468
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 9766 4428 9772 4480
rect 9824 4468 9830 4480
rect 10686 4468 10692 4480
rect 9824 4440 10692 4468
rect 9824 4428 9830 4440
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 11882 4428 11888 4480
rect 11940 4468 11946 4480
rect 12069 4471 12127 4477
rect 12069 4468 12081 4471
rect 11940 4440 12081 4468
rect 11940 4428 11946 4440
rect 12069 4437 12081 4440
rect 12115 4437 12127 4471
rect 12176 4468 12204 4508
rect 12342 4496 12348 4548
rect 12400 4536 12406 4548
rect 12636 4536 12664 4567
rect 12710 4536 12716 4548
rect 12400 4508 12716 4536
rect 12400 4496 12406 4508
rect 12710 4496 12716 4508
rect 12768 4496 12774 4548
rect 15010 4536 15016 4548
rect 13188 4508 15016 4536
rect 13188 4468 13216 4508
rect 15010 4496 15016 4508
rect 15068 4496 15074 4548
rect 12176 4440 13216 4468
rect 13265 4471 13323 4477
rect 12069 4431 12127 4437
rect 13265 4437 13277 4471
rect 13311 4468 13323 4471
rect 13998 4468 14004 4480
rect 13311 4440 14004 4468
rect 13311 4437 13323 4440
rect 13265 4431 13323 4437
rect 13998 4428 14004 4440
rect 14056 4428 14062 4480
rect 14642 4468 14648 4480
rect 14603 4440 14648 4468
rect 14642 4428 14648 4440
rect 14700 4428 14706 4480
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 2590 4224 2596 4276
rect 2648 4264 2654 4276
rect 2774 4264 2780 4276
rect 2648 4236 2780 4264
rect 2648 4224 2654 4236
rect 2774 4224 2780 4236
rect 2832 4224 2838 4276
rect 2866 4224 2872 4276
rect 2924 4264 2930 4276
rect 4798 4264 4804 4276
rect 2924 4236 4804 4264
rect 2924 4224 2930 4236
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 6273 4267 6331 4273
rect 6273 4264 6285 4267
rect 5592 4236 6285 4264
rect 5592 4224 5598 4236
rect 6273 4233 6285 4236
rect 6319 4233 6331 4267
rect 7466 4264 7472 4276
rect 6273 4227 6331 4233
rect 6847 4236 7472 4264
rect 5902 4156 5908 4208
rect 5960 4196 5966 4208
rect 6847 4196 6875 4236
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 8297 4267 8355 4273
rect 8297 4233 8309 4267
rect 8343 4264 8355 4267
rect 8662 4264 8668 4276
rect 8343 4236 8668 4264
rect 8343 4233 8355 4236
rect 8297 4227 8355 4233
rect 8662 4224 8668 4236
rect 8720 4224 8726 4276
rect 9490 4224 9496 4276
rect 9548 4264 9554 4276
rect 9861 4267 9919 4273
rect 9861 4264 9873 4267
rect 9548 4236 9873 4264
rect 9548 4224 9554 4236
rect 9861 4233 9873 4236
rect 9907 4233 9919 4267
rect 9861 4227 9919 4233
rect 10410 4224 10416 4276
rect 10468 4264 10474 4276
rect 11606 4264 11612 4276
rect 10468 4236 11612 4264
rect 10468 4224 10474 4236
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 13630 4264 13636 4276
rect 11716 4236 13636 4264
rect 7926 4196 7932 4208
rect 5960 4168 6875 4196
rect 7852 4168 7932 4196
rect 5960 4156 5966 4168
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4893 4131 4951 4137
rect 4893 4128 4905 4131
rect 4028 4100 4905 4128
rect 4028 4088 4034 4100
rect 4893 4097 4905 4100
rect 4939 4097 4951 4131
rect 4893 4091 4951 4097
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 6638 4128 6644 4140
rect 6052 4100 6644 4128
rect 6052 4088 6058 4100
rect 6638 4088 6644 4100
rect 6696 4128 6702 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6696 4100 6837 4128
rect 6696 4088 6702 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 1394 4060 1400 4072
rect 1307 4032 1400 4060
rect 1394 4020 1400 4032
rect 1452 4060 1458 4072
rect 1664 4063 1722 4069
rect 1452 4032 1624 4060
rect 1452 4020 1458 4032
rect 1596 3992 1624 4032
rect 1664 4029 1676 4063
rect 1710 4060 1722 4063
rect 1710 4032 4752 4060
rect 1710 4029 1722 4032
rect 1664 4023 1722 4029
rect 3136 3995 3194 4001
rect 1596 3964 2820 3992
rect 1670 3884 1676 3936
rect 1728 3924 1734 3936
rect 2682 3924 2688 3936
rect 1728 3896 2688 3924
rect 1728 3884 1734 3896
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 2792 3924 2820 3964
rect 3136 3961 3148 3995
rect 3182 3992 3194 3995
rect 3786 3992 3792 4004
rect 3182 3964 3792 3992
rect 3182 3961 3194 3964
rect 3136 3955 3194 3961
rect 3786 3952 3792 3964
rect 3844 3952 3850 4004
rect 4724 3992 4752 4032
rect 4798 4020 4804 4072
rect 4856 4060 4862 4072
rect 4856 4032 5203 4060
rect 4856 4020 4862 4032
rect 4982 3992 4988 4004
rect 4724 3964 4988 3992
rect 4982 3952 4988 3964
rect 5040 3952 5046 4004
rect 5175 4001 5203 4032
rect 5160 3995 5218 4001
rect 5160 3961 5172 3995
rect 5206 3992 5218 3995
rect 5442 3992 5448 4004
rect 5206 3964 5448 3992
rect 5206 3961 5218 3964
rect 5160 3955 5218 3961
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 6840 3992 6868 4091
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 7081 4063 7139 4069
rect 7081 4060 7093 4063
rect 6972 4032 7093 4060
rect 6972 4020 6978 4032
rect 7081 4029 7093 4032
rect 7127 4029 7139 4063
rect 7081 4023 7139 4029
rect 7852 3992 7880 4168
rect 7926 4156 7932 4168
rect 7984 4156 7990 4208
rect 8754 4156 8760 4208
rect 8812 4196 8818 4208
rect 9769 4199 9827 4205
rect 8812 4168 8892 4196
rect 8812 4156 8818 4168
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 8864 4137 8892 4168
rect 9769 4165 9781 4199
rect 9815 4196 9827 4199
rect 10318 4196 10324 4208
rect 9815 4168 10324 4196
rect 9815 4165 9827 4168
rect 9769 4159 9827 4165
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 11238 4196 11244 4208
rect 10428 4168 11244 4196
rect 10428 4137 10456 4168
rect 11238 4156 11244 4168
rect 11296 4156 11302 4208
rect 11716 4196 11744 4236
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 14182 4224 14188 4276
rect 14240 4264 14246 4276
rect 14458 4264 14464 4276
rect 14240 4236 14464 4264
rect 14240 4224 14246 4236
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 11348 4168 11744 4196
rect 8849 4131 8907 4137
rect 8260 4100 8800 4128
rect 8260 4088 8266 4100
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 7984 4032 8677 4060
rect 7984 4020 7990 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 8772 4060 8800 4100
rect 8849 4097 8861 4131
rect 8895 4097 8907 4131
rect 10413 4131 10471 4137
rect 10413 4128 10425 4131
rect 8849 4091 8907 4097
rect 9048 4100 10425 4128
rect 9048 4060 9076 4100
rect 10413 4097 10425 4100
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 10502 4088 10508 4140
rect 10560 4088 10566 4140
rect 8772 4032 9076 4060
rect 8665 4023 8723 4029
rect 9490 4020 9496 4072
rect 9548 4060 9554 4072
rect 9677 4063 9735 4069
rect 9548 4032 9628 4060
rect 9548 4020 9554 4032
rect 9600 3992 9628 4032
rect 9677 4029 9689 4063
rect 9723 4060 9735 4063
rect 9858 4060 9864 4072
rect 9723 4032 9864 4060
rect 9723 4029 9735 4032
rect 9677 4023 9735 4029
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 10520 4060 10548 4088
rect 11348 4060 11376 4168
rect 12434 4156 12440 4208
rect 12492 4196 12498 4208
rect 12492 4168 12537 4196
rect 12492 4156 12498 4168
rect 13814 4156 13820 4208
rect 13872 4196 13878 4208
rect 13872 4168 14228 4196
rect 13872 4156 13878 4168
rect 11514 4088 11520 4140
rect 11572 4128 11578 4140
rect 11609 4131 11667 4137
rect 11609 4128 11621 4131
rect 11572 4100 11621 4128
rect 11572 4088 11578 4100
rect 11609 4097 11621 4100
rect 11655 4097 11667 4131
rect 11609 4091 11667 4097
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 11848 4100 13001 4128
rect 11848 4088 11854 4100
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13630 4088 13636 4140
rect 13688 4128 13694 4140
rect 14200 4137 14228 4168
rect 14185 4131 14243 4137
rect 13688 4100 14136 4128
rect 13688 4088 13694 4100
rect 10275 4032 11376 4060
rect 11425 4063 11483 4069
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 11425 4029 11437 4063
rect 11471 4060 11483 4063
rect 11698 4060 11704 4072
rect 11471 4032 11704 4060
rect 11471 4029 11483 4032
rect 11425 4023 11483 4029
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12544 4032 12817 4060
rect 9769 3995 9827 4001
rect 9769 3992 9781 3995
rect 6840 3964 9536 3992
rect 9600 3964 9781 3992
rect 3970 3924 3976 3936
rect 2792 3896 3976 3924
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 4249 3927 4307 3933
rect 4249 3893 4261 3927
rect 4295 3924 4307 3927
rect 5534 3924 5540 3936
rect 4295 3896 5540 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 7340 3896 8217 3924
rect 7340 3884 7346 3896
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 8205 3887 8263 3893
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 9508 3933 9536 3964
rect 9769 3961 9781 3964
rect 9815 3961 9827 3995
rect 9769 3955 9827 3961
rect 9950 3952 9956 4004
rect 10008 3992 10014 4004
rect 10870 3992 10876 4004
rect 10008 3964 10876 3992
rect 10008 3952 10014 3964
rect 10870 3952 10876 3964
rect 10928 3952 10934 4004
rect 10962 3952 10968 4004
rect 11020 3952 11026 4004
rect 12544 3992 12572 4032
rect 12805 4029 12817 4032
rect 12851 4029 12863 4063
rect 13998 4060 14004 4072
rect 13959 4032 14004 4060
rect 12805 4023 12863 4029
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14108 4060 14136 4100
rect 14185 4097 14197 4131
rect 14231 4097 14243 4131
rect 14185 4091 14243 4097
rect 14642 4060 14648 4072
rect 14108 4032 14648 4060
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 14829 4063 14887 4069
rect 14829 4029 14841 4063
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 11072 3964 12572 3992
rect 9493 3927 9551 3933
rect 8812 3896 8857 3924
rect 8812 3884 8818 3896
rect 9493 3893 9505 3927
rect 9539 3893 9551 3927
rect 9493 3887 9551 3893
rect 10226 3884 10232 3936
rect 10284 3924 10290 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 10284 3896 10333 3924
rect 10284 3884 10290 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 10321 3887 10379 3893
rect 10502 3884 10508 3936
rect 10560 3924 10566 3936
rect 10980 3924 11008 3952
rect 11072 3933 11100 3964
rect 13262 3952 13268 4004
rect 13320 3992 13326 4004
rect 14844 3992 14872 4023
rect 13320 3964 14872 3992
rect 13320 3952 13326 3964
rect 10560 3896 11008 3924
rect 11057 3927 11115 3933
rect 10560 3884 10566 3896
rect 11057 3893 11069 3927
rect 11103 3893 11115 3927
rect 11057 3887 11115 3893
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11388 3896 11529 3924
rect 11388 3884 11394 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 11664 3896 12909 3924
rect 11664 3884 11670 3896
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 13630 3924 13636 3936
rect 13591 3896 13636 3924
rect 12897 3887 12955 3893
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 14093 3927 14151 3933
rect 14093 3924 14105 3927
rect 13872 3896 14105 3924
rect 13872 3884 13878 3896
rect 14093 3893 14105 3896
rect 14139 3893 14151 3927
rect 15010 3924 15016 3936
rect 14971 3896 15016 3924
rect 14093 3887 14151 3893
rect 15010 3884 15016 3896
rect 15068 3884 15074 3936
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 2869 3723 2927 3729
rect 2869 3689 2881 3723
rect 2915 3720 2927 3723
rect 4433 3723 4491 3729
rect 4433 3720 4445 3723
rect 2915 3692 4445 3720
rect 2915 3689 2927 3692
rect 2869 3683 2927 3689
rect 4433 3689 4445 3692
rect 4479 3689 4491 3723
rect 4433 3683 4491 3689
rect 4614 3680 4620 3732
rect 4672 3720 4678 3732
rect 4672 3692 4936 3720
rect 4672 3680 4678 3692
rect 1664 3655 1722 3661
rect 1664 3621 1676 3655
rect 1710 3652 1722 3655
rect 2038 3652 2044 3664
rect 1710 3624 2044 3652
rect 1710 3621 1722 3624
rect 1664 3615 1722 3621
rect 2038 3612 2044 3624
rect 2096 3612 2102 3664
rect 2958 3612 2964 3664
rect 3016 3652 3022 3664
rect 3329 3655 3387 3661
rect 3329 3652 3341 3655
rect 3016 3624 3341 3652
rect 3016 3612 3022 3624
rect 3329 3621 3341 3624
rect 3375 3652 3387 3655
rect 3878 3652 3884 3664
rect 3375 3624 3884 3652
rect 3375 3621 3387 3624
rect 3329 3615 3387 3621
rect 3878 3612 3884 3624
rect 3936 3612 3942 3664
rect 4525 3655 4583 3661
rect 4525 3621 4537 3655
rect 4571 3652 4583 3655
rect 4798 3652 4804 3664
rect 4571 3624 4804 3652
rect 4571 3621 4583 3624
rect 4525 3615 4583 3621
rect 4798 3612 4804 3624
rect 4856 3612 4862 3664
rect 4908 3652 4936 3692
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 5500 3692 6837 3720
rect 5500 3680 5506 3692
rect 6825 3689 6837 3692
rect 6871 3720 6883 3723
rect 6914 3720 6920 3732
rect 6871 3692 6920 3720
rect 6871 3689 6883 3692
rect 6825 3683 6883 3689
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 7190 3680 7196 3732
rect 7248 3720 7254 3732
rect 7377 3723 7435 3729
rect 7377 3720 7389 3723
rect 7248 3692 7389 3720
rect 7248 3680 7254 3692
rect 7377 3689 7389 3692
rect 7423 3689 7435 3723
rect 7377 3683 7435 3689
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 7524 3692 8953 3720
rect 7524 3680 7530 3692
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 8941 3683 8999 3689
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 10318 3720 10324 3732
rect 9088 3692 10324 3720
rect 9088 3680 9094 3692
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 10873 3723 10931 3729
rect 10873 3689 10885 3723
rect 10919 3720 10931 3723
rect 11606 3720 11612 3732
rect 10919 3692 11612 3720
rect 10919 3689 10931 3692
rect 10873 3683 10931 3689
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 12069 3723 12127 3729
rect 12069 3720 12081 3723
rect 11940 3692 12081 3720
rect 11940 3680 11946 3692
rect 12069 3689 12081 3692
rect 12115 3689 12127 3723
rect 12894 3720 12900 3732
rect 12855 3692 12900 3720
rect 12069 3683 12127 3689
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 13262 3720 13268 3732
rect 13223 3692 13268 3720
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 14737 3723 14795 3729
rect 14737 3720 14749 3723
rect 13780 3692 14749 3720
rect 13780 3680 13786 3692
rect 14737 3689 14749 3692
rect 14783 3689 14795 3723
rect 14737 3683 14795 3689
rect 5718 3661 5724 3664
rect 5701 3655 5724 3661
rect 5701 3652 5713 3655
rect 4908 3624 5713 3652
rect 5701 3621 5713 3624
rect 5776 3652 5782 3664
rect 6546 3652 6552 3664
rect 5776 3624 6552 3652
rect 5701 3615 5724 3621
rect 5718 3612 5724 3615
rect 5776 3612 5782 3624
rect 6546 3612 6552 3624
rect 6604 3612 6610 3664
rect 7285 3655 7343 3661
rect 7285 3621 7297 3655
rect 7331 3652 7343 3655
rect 7650 3652 7656 3664
rect 7331 3624 7656 3652
rect 7331 3621 7343 3624
rect 7285 3615 7343 3621
rect 7650 3612 7656 3624
rect 7708 3612 7714 3664
rect 8205 3655 8263 3661
rect 8205 3621 8217 3655
rect 8251 3652 8263 3655
rect 9674 3652 9680 3664
rect 8251 3624 9680 3652
rect 8251 3621 8263 3624
rect 8205 3615 8263 3621
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 10410 3612 10416 3664
rect 10468 3652 10474 3664
rect 11238 3652 11244 3664
rect 10468 3624 11008 3652
rect 11199 3624 11244 3652
rect 10468 3612 10474 3624
rect 3237 3587 3295 3593
rect 3237 3553 3249 3587
rect 3283 3553 3295 3587
rect 3237 3547 3295 3553
rect 3252 3448 3280 3547
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4893 3587 4951 3593
rect 4028 3556 4743 3584
rect 4028 3544 4034 3556
rect 3513 3519 3571 3525
rect 3513 3485 3525 3519
rect 3559 3516 3571 3519
rect 3786 3516 3792 3528
rect 3559 3488 3792 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 3786 3476 3792 3488
rect 3844 3516 3850 3528
rect 4154 3516 4160 3528
rect 3844 3488 4160 3516
rect 3844 3476 3850 3488
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4614 3516 4620 3528
rect 4575 3488 4620 3516
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 4430 3448 4436 3460
rect 3252 3420 4436 3448
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 4715 3448 4743 3556
rect 4893 3553 4905 3587
rect 4939 3584 4951 3587
rect 7834 3584 7840 3596
rect 4939 3556 7840 3584
rect 4939 3553 4951 3556
rect 4893 3547 4951 3553
rect 7834 3544 7840 3556
rect 7892 3544 7898 3596
rect 8110 3584 8116 3596
rect 8071 3556 8116 3584
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 8220 3556 9352 3584
rect 5074 3516 5080 3528
rect 5035 3488 5080 3516
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 5445 3519 5503 3525
rect 5445 3485 5457 3519
rect 5491 3485 5503 3519
rect 5445 3479 5503 3485
rect 5460 3448 5488 3479
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 7469 3519 7527 3525
rect 7469 3516 7481 3519
rect 6972 3488 7481 3516
rect 6972 3476 6978 3488
rect 7469 3485 7481 3488
rect 7515 3485 7527 3519
rect 8220 3516 8248 3556
rect 8386 3516 8392 3528
rect 7469 3479 7527 3485
rect 7576 3488 8248 3516
rect 8347 3488 8392 3516
rect 7576 3448 7604 3488
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 9033 3519 9091 3525
rect 9033 3516 9045 3519
rect 8496 3488 9045 3516
rect 4715 3420 5488 3448
rect 6847 3420 7604 3448
rect 7745 3451 7803 3457
rect 2777 3383 2835 3389
rect 2777 3349 2789 3383
rect 2823 3380 2835 3383
rect 2866 3380 2872 3392
rect 2823 3352 2872 3380
rect 2823 3349 2835 3352
rect 2777 3343 2835 3349
rect 2866 3340 2872 3352
rect 2924 3340 2930 3392
rect 3878 3340 3884 3392
rect 3936 3380 3942 3392
rect 4065 3383 4123 3389
rect 4065 3380 4077 3383
rect 3936 3352 4077 3380
rect 3936 3340 3942 3352
rect 4065 3349 4077 3352
rect 4111 3349 4123 3383
rect 4065 3343 4123 3349
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 5166 3380 5172 3392
rect 4212 3352 5172 3380
rect 4212 3340 4218 3352
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 5258 3340 5264 3392
rect 5316 3380 5322 3392
rect 6847 3380 6875 3420
rect 7745 3417 7757 3451
rect 7791 3448 7803 3451
rect 8496 3448 8524 3488
rect 9033 3485 9045 3488
rect 9079 3485 9091 3519
rect 9214 3516 9220 3528
rect 9175 3488 9220 3516
rect 9033 3479 9091 3485
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 7791 3420 8524 3448
rect 7791 3417 7803 3420
rect 7745 3411 7803 3417
rect 8570 3408 8576 3460
rect 8628 3448 8634 3460
rect 8628 3420 8673 3448
rect 8628 3408 8634 3420
rect 5316 3352 6875 3380
rect 6917 3383 6975 3389
rect 5316 3340 5322 3352
rect 6917 3349 6929 3383
rect 6963 3380 6975 3383
rect 8846 3380 8852 3392
rect 6963 3352 8852 3380
rect 6963 3349 6975 3352
rect 6917 3343 6975 3349
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 9324 3380 9352 3556
rect 9490 3544 9496 3596
rect 9548 3544 9554 3596
rect 9766 3544 9772 3596
rect 9824 3584 9830 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 9824 3556 10057 3584
rect 9824 3544 9830 3556
rect 10045 3553 10057 3556
rect 10091 3584 10103 3587
rect 10091 3556 10916 3584
rect 10091 3553 10103 3556
rect 10045 3547 10103 3553
rect 9508 3516 9536 3544
rect 9674 3516 9680 3528
rect 9508 3488 9680 3516
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 10137 3519 10195 3525
rect 10137 3485 10149 3519
rect 10183 3516 10195 3519
rect 10226 3516 10232 3528
rect 10183 3488 10232 3516
rect 10183 3485 10195 3488
rect 10137 3479 10195 3485
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3516 10379 3519
rect 10367 3488 10456 3516
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 9490 3408 9496 3460
rect 9548 3448 9554 3460
rect 9766 3448 9772 3460
rect 9548 3420 9772 3448
rect 9548 3408 9554 3420
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 9677 3383 9735 3389
rect 9677 3380 9689 3383
rect 9324 3352 9689 3380
rect 9677 3349 9689 3352
rect 9723 3349 9735 3383
rect 10428 3380 10456 3488
rect 10888 3448 10916 3556
rect 10980 3516 11008 3624
rect 11238 3612 11244 3624
rect 11296 3612 11302 3664
rect 11333 3655 11391 3661
rect 11333 3621 11345 3655
rect 11379 3652 11391 3655
rect 12158 3652 12164 3664
rect 11379 3624 12164 3652
rect 11379 3621 11391 3624
rect 11333 3615 11391 3621
rect 12158 3612 12164 3624
rect 12216 3612 12222 3664
rect 12526 3652 12532 3664
rect 12487 3624 12532 3652
rect 12526 3612 12532 3624
rect 12584 3612 12590 3664
rect 13354 3652 13360 3664
rect 13315 3624 13360 3652
rect 13354 3612 13360 3624
rect 13412 3612 13418 3664
rect 13446 3612 13452 3664
rect 13504 3652 13510 3664
rect 13504 3624 14320 3652
rect 13504 3612 13510 3624
rect 11054 3544 11060 3596
rect 11112 3584 11118 3596
rect 12437 3587 12495 3593
rect 12437 3584 12449 3587
rect 11112 3556 12449 3584
rect 11112 3544 11118 3556
rect 12437 3553 12449 3556
rect 12483 3584 12495 3587
rect 14090 3584 14096 3596
rect 12483 3556 13952 3584
rect 14051 3556 14096 3584
rect 12483 3553 12495 3556
rect 12437 3547 12495 3553
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 10980 3488 11437 3516
rect 11425 3485 11437 3488
rect 11471 3516 11483 3519
rect 11514 3516 11520 3528
rect 11471 3488 11520 3516
rect 11471 3485 11483 3488
rect 11425 3479 11483 3485
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 12710 3516 12716 3528
rect 12671 3488 12716 3516
rect 12710 3476 12716 3488
rect 12768 3516 12774 3528
rect 12986 3516 12992 3528
rect 12768 3488 12992 3516
rect 12768 3476 12774 3488
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 13170 3476 13176 3528
rect 13228 3516 13234 3528
rect 13449 3519 13507 3525
rect 13449 3516 13461 3519
rect 13228 3488 13461 3516
rect 13228 3476 13234 3488
rect 13449 3485 13461 3488
rect 13495 3485 13507 3519
rect 13449 3479 13507 3485
rect 13078 3448 13084 3460
rect 10888 3420 13084 3448
rect 13078 3408 13084 3420
rect 13136 3408 13142 3460
rect 13262 3408 13268 3460
rect 13320 3408 13326 3460
rect 13924 3448 13952 3556
rect 14090 3544 14096 3556
rect 14148 3544 14154 3596
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14292 3525 14320 3624
rect 14458 3544 14464 3596
rect 14516 3584 14522 3596
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 14516 3556 14565 3584
rect 14516 3544 14522 3556
rect 14553 3553 14565 3556
rect 14599 3553 14611 3587
rect 14553 3547 14611 3553
rect 14185 3519 14243 3525
rect 14185 3516 14197 3519
rect 14056 3488 14197 3516
rect 14056 3476 14062 3488
rect 14185 3485 14197 3488
rect 14231 3485 14243 3519
rect 14185 3479 14243 3485
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 14458 3448 14464 3460
rect 13924 3420 14464 3448
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 10594 3380 10600 3392
rect 10428 3352 10600 3380
rect 9677 3343 9735 3349
rect 10594 3340 10600 3352
rect 10652 3380 10658 3392
rect 11974 3380 11980 3392
rect 10652 3352 11980 3380
rect 10652 3340 10658 3352
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 12434 3340 12440 3392
rect 12492 3380 12498 3392
rect 13280 3380 13308 3408
rect 12492 3352 13308 3380
rect 13725 3383 13783 3389
rect 12492 3340 12498 3352
rect 13725 3349 13737 3383
rect 13771 3380 13783 3383
rect 15286 3380 15292 3392
rect 13771 3352 15292 3380
rect 13771 3349 13783 3352
rect 13725 3343 13783 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 2038 3136 2044 3188
rect 2096 3176 2102 3188
rect 6730 3176 6736 3188
rect 2096 3148 4200 3176
rect 2096 3136 2102 3148
rect 4172 3108 4200 3148
rect 4356 3148 6736 3176
rect 4356 3108 4384 3148
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 7524 3148 8217 3176
rect 7524 3136 7530 3148
rect 8205 3145 8217 3148
rect 8251 3145 8263 3179
rect 8205 3139 8263 3145
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3176 8355 3179
rect 9122 3176 9128 3188
rect 8343 3148 9128 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 9493 3179 9551 3185
rect 9493 3145 9505 3179
rect 9539 3176 9551 3179
rect 9582 3176 9588 3188
rect 9539 3148 9588 3176
rect 9539 3145 9551 3148
rect 9493 3139 9551 3145
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 10962 3176 10968 3188
rect 10284 3148 10968 3176
rect 10284 3136 10290 3148
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 11057 3179 11115 3185
rect 11057 3145 11069 3179
rect 11103 3176 11115 3179
rect 12526 3176 12532 3188
rect 11103 3148 12532 3176
rect 11103 3145 11115 3148
rect 11057 3139 11115 3145
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 14090 3176 14096 3188
rect 13136 3148 14096 3176
rect 13136 3136 13142 3148
rect 14090 3136 14096 3148
rect 14148 3136 14154 3188
rect 14366 3136 14372 3188
rect 14424 3176 14430 3188
rect 14461 3179 14519 3185
rect 14461 3176 14473 3179
rect 14424 3148 14473 3176
rect 14424 3136 14430 3148
rect 14461 3145 14473 3148
rect 14507 3145 14519 3179
rect 14461 3139 14519 3145
rect 4172 3080 4384 3108
rect 5350 3068 5356 3120
rect 5408 3108 5414 3120
rect 5721 3111 5779 3117
rect 5721 3108 5733 3111
rect 5408 3080 5733 3108
rect 5408 3068 5414 3080
rect 5721 3077 5733 3080
rect 5767 3077 5779 3111
rect 5721 3071 5779 3077
rect 7834 3068 7840 3120
rect 7892 3108 7898 3120
rect 12253 3111 12311 3117
rect 7892 3080 12020 3108
rect 7892 3068 7898 3080
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 5626 3000 5632 3052
rect 5684 3040 5690 3052
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 5684 3012 6377 3040
rect 5684 3000 5690 3012
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6696 3012 6837 3040
rect 6696 3000 6702 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 7926 3000 7932 3052
rect 7984 3040 7990 3052
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 7984 3012 8861 3040
rect 7984 3000 7990 3012
rect 8849 3009 8861 3012
rect 8895 3009 8907 3043
rect 8849 3003 8907 3009
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 9088 3012 10425 3040
rect 9088 3000 9094 3012
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 10686 3000 10692 3052
rect 10744 3040 10750 3052
rect 11609 3043 11667 3049
rect 11609 3040 11621 3043
rect 10744 3012 11621 3040
rect 10744 3000 10750 3012
rect 11609 3009 11621 3012
rect 11655 3009 11667 3043
rect 11609 3003 11667 3009
rect 11882 3000 11888 3052
rect 11940 3000 11946 3052
rect 11992 3040 12020 3080
rect 12253 3077 12265 3111
rect 12299 3108 12311 3111
rect 12437 3111 12495 3117
rect 12437 3108 12449 3111
rect 12299 3080 12449 3108
rect 12299 3077 12311 3080
rect 12253 3071 12311 3077
rect 12437 3077 12449 3080
rect 12483 3077 12495 3111
rect 13633 3111 13691 3117
rect 13633 3108 13645 3111
rect 12437 3071 12495 3077
rect 12544 3080 13645 3108
rect 12544 3040 12572 3080
rect 13633 3077 13645 3080
rect 13679 3077 13691 3111
rect 13998 3108 14004 3120
rect 13633 3071 13691 3077
rect 13740 3080 14004 3108
rect 13078 3040 13084 3052
rect 11992 3012 12572 3040
rect 13039 3012 13084 3040
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 13740 3040 13768 3080
rect 13998 3068 14004 3080
rect 14056 3068 14062 3120
rect 14090 3040 14096 3052
rect 13464 3012 13768 3040
rect 14051 3012 14096 3040
rect 5166 2972 5172 2984
rect 2332 2944 5172 2972
rect 2332 2916 2360 2944
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 6273 2975 6331 2981
rect 6273 2941 6285 2975
rect 6319 2972 6331 2975
rect 6454 2972 6460 2984
rect 6319 2944 6460 2972
rect 6319 2941 6331 2944
rect 6273 2935 6331 2941
rect 6454 2932 6460 2944
rect 6512 2932 6518 2984
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 8386 2972 8392 2984
rect 6604 2944 8392 2972
rect 6604 2932 6610 2944
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 8478 2932 8484 2984
rect 8536 2972 8542 2984
rect 9214 2972 9220 2984
rect 8536 2944 9220 2972
rect 8536 2932 8542 2944
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 9677 2975 9735 2981
rect 9677 2941 9689 2975
rect 9723 2972 9735 2975
rect 9858 2972 9864 2984
rect 9723 2944 9864 2972
rect 9723 2941 9735 2944
rect 9677 2935 9735 2941
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 11900 2972 11928 3000
rect 10060 2944 11928 2972
rect 12253 2975 12311 2981
rect 1664 2907 1722 2913
rect 1664 2873 1676 2907
rect 1710 2904 1722 2907
rect 1854 2904 1860 2916
rect 1710 2876 1860 2904
rect 1710 2873 1722 2876
rect 1664 2867 1722 2873
rect 1854 2864 1860 2876
rect 1912 2864 1918 2916
rect 2314 2864 2320 2916
rect 2372 2864 2378 2916
rect 3136 2907 3194 2913
rect 3136 2873 3148 2907
rect 3182 2904 3194 2907
rect 4430 2904 4436 2916
rect 3182 2876 4436 2904
rect 3182 2873 3194 2876
rect 3136 2867 3194 2873
rect 4430 2864 4436 2876
rect 4488 2864 4494 2916
rect 4608 2907 4666 2913
rect 4608 2873 4620 2907
rect 4654 2904 4666 2907
rect 6181 2907 6239 2913
rect 4654 2876 6132 2904
rect 4654 2873 4666 2876
rect 4608 2867 4666 2873
rect 2777 2839 2835 2845
rect 2777 2805 2789 2839
rect 2823 2836 2835 2839
rect 4154 2836 4160 2848
rect 2823 2808 4160 2836
rect 2823 2805 2835 2808
rect 2777 2799 2835 2805
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 4249 2839 4307 2845
rect 4249 2805 4261 2839
rect 4295 2836 4307 2839
rect 4338 2836 4344 2848
rect 4295 2808 4344 2836
rect 4295 2805 4307 2808
rect 4249 2799 4307 2805
rect 4338 2796 4344 2808
rect 4396 2796 4402 2848
rect 5810 2796 5816 2848
rect 5868 2836 5874 2848
rect 6104 2836 6132 2876
rect 6181 2873 6193 2907
rect 6227 2904 6239 2907
rect 6362 2904 6368 2916
rect 6227 2876 6368 2904
rect 6227 2873 6239 2876
rect 6181 2867 6239 2873
rect 6362 2864 6368 2876
rect 6420 2864 6426 2916
rect 7092 2907 7150 2913
rect 7092 2873 7104 2907
rect 7138 2904 7150 2907
rect 9306 2904 9312 2916
rect 7138 2876 9312 2904
rect 7138 2873 7150 2876
rect 7092 2867 7150 2873
rect 9306 2864 9312 2876
rect 9364 2864 9370 2916
rect 10060 2904 10088 2944
rect 12253 2941 12265 2975
rect 12299 2972 12311 2975
rect 12618 2972 12624 2984
rect 12299 2944 12624 2972
rect 12299 2941 12311 2944
rect 12253 2935 12311 2941
rect 12618 2932 12624 2944
rect 12676 2932 12682 2984
rect 12710 2932 12716 2984
rect 12768 2972 12774 2984
rect 12805 2975 12863 2981
rect 12805 2972 12817 2975
rect 12768 2944 12817 2972
rect 12768 2932 12774 2944
rect 12805 2941 12817 2944
rect 12851 2972 12863 2975
rect 13354 2972 13360 2984
rect 12851 2944 13360 2972
rect 12851 2941 12863 2944
rect 12805 2935 12863 2941
rect 13354 2932 13360 2944
rect 13412 2932 13418 2984
rect 9699 2876 10088 2904
rect 6270 2836 6276 2848
rect 5868 2808 5913 2836
rect 6104 2808 6276 2836
rect 5868 2796 5874 2808
rect 6270 2796 6276 2808
rect 6328 2796 6334 2848
rect 6638 2796 6644 2848
rect 6696 2836 6702 2848
rect 7006 2836 7012 2848
rect 6696 2808 7012 2836
rect 6696 2796 6702 2808
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 8570 2796 8576 2848
rect 8628 2836 8634 2848
rect 8665 2839 8723 2845
rect 8665 2836 8677 2839
rect 8628 2808 8677 2836
rect 8628 2796 8634 2808
rect 8665 2805 8677 2808
rect 8711 2805 8723 2839
rect 8665 2799 8723 2805
rect 8757 2839 8815 2845
rect 8757 2805 8769 2839
rect 8803 2836 8815 2839
rect 9699 2836 9727 2876
rect 10134 2864 10140 2916
rect 10192 2904 10198 2916
rect 10229 2907 10287 2913
rect 10229 2904 10241 2907
rect 10192 2876 10241 2904
rect 10192 2864 10198 2876
rect 10229 2873 10241 2876
rect 10275 2873 10287 2907
rect 10229 2867 10287 2873
rect 10318 2864 10324 2916
rect 10376 2904 10382 2916
rect 10376 2876 10421 2904
rect 10376 2864 10382 2876
rect 10594 2864 10600 2916
rect 10652 2904 10658 2916
rect 11517 2907 11575 2913
rect 11517 2904 11529 2907
rect 10652 2876 11529 2904
rect 10652 2864 10658 2876
rect 11517 2873 11529 2876
rect 11563 2904 11575 2907
rect 13464 2904 13492 3012
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14185 3043 14243 3049
rect 14185 3009 14197 3043
rect 14231 3009 14243 3043
rect 14185 3003 14243 3009
rect 13538 2932 13544 2984
rect 13596 2972 13602 2984
rect 14200 2972 14228 3003
rect 14826 3000 14832 3052
rect 14884 3040 14890 3052
rect 15013 3043 15071 3049
rect 15013 3040 15025 3043
rect 14884 3012 15025 3040
rect 14884 3000 14890 3012
rect 15013 3009 15025 3012
rect 15059 3009 15071 3043
rect 15013 3003 15071 3009
rect 13596 2944 14228 2972
rect 14921 2975 14979 2981
rect 13596 2932 13602 2944
rect 14921 2941 14933 2975
rect 14967 2972 14979 2975
rect 15286 2972 15292 2984
rect 14967 2944 15292 2972
rect 14967 2941 14979 2944
rect 14921 2935 14979 2941
rect 15286 2932 15292 2944
rect 15344 2932 15350 2984
rect 11563 2876 13492 2904
rect 11563 2873 11575 2876
rect 11517 2867 11575 2873
rect 13906 2864 13912 2916
rect 13964 2904 13970 2916
rect 14001 2907 14059 2913
rect 14001 2904 14013 2907
rect 13964 2876 14013 2904
rect 13964 2864 13970 2876
rect 14001 2873 14013 2876
rect 14047 2873 14059 2907
rect 14001 2867 14059 2873
rect 9858 2836 9864 2848
rect 8803 2808 9727 2836
rect 9819 2808 9864 2836
rect 8803 2805 8815 2808
rect 8757 2799 8815 2805
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 11422 2836 11428 2848
rect 11383 2808 11428 2836
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 12897 2839 12955 2845
rect 12897 2836 12909 2839
rect 11664 2808 12909 2836
rect 11664 2796 11670 2808
rect 12897 2805 12909 2808
rect 12943 2805 12955 2839
rect 12897 2799 12955 2805
rect 14458 2796 14464 2848
rect 14516 2836 14522 2848
rect 14829 2839 14887 2845
rect 14829 2836 14841 2839
rect 14516 2808 14841 2836
rect 14516 2796 14522 2808
rect 14829 2805 14841 2808
rect 14875 2805 14887 2839
rect 14829 2799 14887 2805
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 1762 2592 1768 2644
rect 1820 2632 1826 2644
rect 2774 2632 2780 2644
rect 1820 2604 2780 2632
rect 1820 2592 1826 2604
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 2866 2592 2872 2644
rect 2924 2632 2930 2644
rect 2924 2604 5396 2632
rect 2924 2592 2930 2604
rect 1673 2567 1731 2573
rect 1673 2533 1685 2567
rect 1719 2564 1731 2567
rect 1946 2564 1952 2576
rect 1719 2536 1952 2564
rect 1719 2533 1731 2536
rect 1673 2527 1731 2533
rect 1946 2524 1952 2536
rect 2004 2524 2010 2576
rect 3050 2524 3056 2576
rect 3108 2524 3114 2576
rect 3326 2524 3332 2576
rect 3384 2564 3390 2576
rect 4332 2567 4390 2573
rect 3384 2536 4292 2564
rect 3384 2524 3390 2536
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 2222 2496 2228 2508
rect 1443 2468 2228 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 2400 2499 2458 2505
rect 2400 2465 2412 2499
rect 2446 2496 2458 2499
rect 2774 2496 2780 2508
rect 2446 2468 2780 2496
rect 2446 2465 2458 2468
rect 2400 2459 2458 2465
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 3068 2496 3096 2524
rect 3605 2499 3663 2505
rect 3605 2496 3617 2499
rect 3068 2468 3617 2496
rect 3605 2465 3617 2468
rect 3651 2496 3663 2499
rect 3786 2496 3792 2508
rect 3651 2468 3792 2496
rect 3651 2465 3663 2468
rect 3605 2459 3663 2465
rect 3786 2456 3792 2468
rect 3844 2456 3850 2508
rect 4264 2496 4292 2536
rect 4332 2533 4344 2567
rect 4378 2564 4390 2567
rect 4430 2564 4436 2576
rect 4378 2536 4436 2564
rect 4378 2533 4390 2536
rect 4332 2527 4390 2533
rect 4430 2524 4436 2536
rect 4488 2524 4494 2576
rect 5368 2564 5396 2604
rect 5442 2592 5448 2644
rect 5500 2632 5506 2644
rect 5537 2635 5595 2641
rect 5537 2632 5549 2635
rect 5500 2604 5549 2632
rect 5500 2592 5506 2604
rect 5537 2601 5549 2604
rect 5583 2601 5595 2635
rect 5537 2595 5595 2601
rect 5626 2592 5632 2644
rect 5684 2632 5690 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5684 2604 6009 2632
rect 5684 2592 5690 2604
rect 5997 2601 6009 2604
rect 6043 2632 6055 2635
rect 7190 2632 7196 2644
rect 6043 2604 7196 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 7285 2635 7343 2641
rect 7285 2601 7297 2635
rect 7331 2632 7343 2635
rect 7742 2632 7748 2644
rect 7331 2604 7748 2632
rect 7331 2601 7343 2604
rect 7285 2595 7343 2601
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 8754 2632 8760 2644
rect 8619 2604 8760 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 8754 2592 8760 2604
rect 8812 2592 8818 2644
rect 8846 2592 8852 2644
rect 8904 2632 8910 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8904 2604 8953 2632
rect 8904 2592 8910 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 9858 2592 9864 2644
rect 9916 2632 9922 2644
rect 10229 2635 10287 2641
rect 10229 2632 10241 2635
rect 9916 2604 10241 2632
rect 9916 2592 9922 2604
rect 10229 2601 10241 2604
rect 10275 2601 10287 2635
rect 10229 2595 10287 2601
rect 10965 2635 11023 2641
rect 10965 2601 10977 2635
rect 11011 2601 11023 2635
rect 10965 2595 11023 2601
rect 11425 2635 11483 2641
rect 11425 2601 11437 2635
rect 11471 2632 11483 2635
rect 13630 2632 13636 2644
rect 11471 2604 13636 2632
rect 11471 2601 11483 2604
rect 11425 2595 11483 2601
rect 8113 2567 8171 2573
rect 5368 2536 6592 2564
rect 5902 2496 5908 2508
rect 4264 2468 5120 2496
rect 5863 2468 5908 2496
rect 1486 2388 1492 2440
rect 1544 2428 1550 2440
rect 2133 2431 2191 2437
rect 2133 2428 2145 2431
rect 1544 2400 2145 2428
rect 1544 2388 1550 2400
rect 2133 2397 2145 2400
rect 2179 2397 2191 2431
rect 2133 2391 2191 2397
rect 3789 2363 3847 2369
rect 3789 2360 3801 2363
rect 3068 2332 3801 2360
rect 198 2252 204 2304
rect 256 2292 262 2304
rect 3068 2292 3096 2332
rect 3789 2329 3801 2332
rect 3835 2329 3847 2363
rect 5092 2360 5120 2468
rect 5902 2456 5908 2468
rect 5960 2456 5966 2508
rect 6365 2499 6423 2505
rect 6365 2465 6377 2499
rect 6411 2496 6423 2499
rect 6454 2496 6460 2508
rect 6411 2468 6460 2496
rect 6411 2465 6423 2468
rect 6365 2459 6423 2465
rect 6454 2456 6460 2468
rect 6512 2456 6518 2508
rect 6089 2431 6147 2437
rect 6089 2428 6101 2431
rect 6012 2400 6101 2428
rect 6012 2372 6040 2400
rect 6089 2397 6101 2400
rect 6135 2397 6147 2431
rect 6564 2428 6592 2536
rect 8113 2533 8125 2567
rect 8159 2564 8171 2567
rect 8159 2536 8616 2564
rect 8159 2533 8171 2536
rect 8113 2527 8171 2533
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 7377 2499 7435 2505
rect 7377 2496 7389 2499
rect 6788 2468 7389 2496
rect 6788 2456 6794 2468
rect 7377 2465 7389 2468
rect 7423 2465 7435 2499
rect 7377 2459 7435 2465
rect 7558 2456 7564 2508
rect 7616 2496 7622 2508
rect 8588 2496 8616 2536
rect 8662 2524 8668 2576
rect 8720 2564 8726 2576
rect 9033 2567 9091 2573
rect 9033 2564 9045 2567
rect 8720 2536 9045 2564
rect 8720 2524 8726 2536
rect 9033 2533 9045 2536
rect 9079 2533 9091 2567
rect 10980 2564 11008 2595
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 13817 2635 13875 2641
rect 13817 2601 13829 2635
rect 13863 2632 13875 2635
rect 14090 2632 14096 2644
rect 13863 2604 14096 2632
rect 13863 2601 13875 2604
rect 13817 2595 13875 2601
rect 14090 2592 14096 2604
rect 14148 2592 14154 2644
rect 14274 2632 14280 2644
rect 14235 2604 14280 2632
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 11698 2564 11704 2576
rect 10980 2536 11704 2564
rect 9033 2527 9091 2533
rect 11698 2524 11704 2536
rect 11756 2524 11762 2576
rect 12802 2524 12808 2576
rect 12860 2564 12866 2576
rect 12989 2567 13047 2573
rect 12989 2564 13001 2567
rect 12860 2536 13001 2564
rect 12860 2524 12866 2536
rect 12989 2533 13001 2536
rect 13035 2533 13047 2567
rect 14182 2564 14188 2576
rect 14143 2536 14188 2564
rect 12989 2527 13047 2533
rect 14182 2524 14188 2536
rect 14240 2524 14246 2576
rect 8938 2496 8944 2508
rect 7616 2468 8340 2496
rect 8588 2468 8944 2496
rect 7616 2456 7622 2468
rect 8312 2437 8340 2468
rect 8938 2456 8944 2468
rect 8996 2456 9002 2508
rect 10137 2499 10195 2505
rect 10137 2465 10149 2499
rect 10183 2496 10195 2499
rect 11330 2496 11336 2508
rect 10183 2468 10824 2496
rect 11291 2468 11336 2496
rect 10183 2465 10195 2468
rect 10137 2459 10195 2465
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 6564 2400 7481 2428
rect 6089 2391 6147 2397
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 5092 2332 5571 2360
rect 3789 2323 3847 2329
rect 256 2264 3096 2292
rect 3513 2295 3571 2301
rect 256 2252 262 2264
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 3878 2292 3884 2304
rect 3559 2264 3884 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 3878 2252 3884 2264
rect 3936 2252 3942 2304
rect 4706 2252 4712 2304
rect 4764 2292 4770 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 4764 2264 5457 2292
rect 4764 2252 4770 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5543 2292 5571 2332
rect 5994 2320 6000 2372
rect 6052 2320 6058 2372
rect 6546 2360 6552 2372
rect 6507 2332 6552 2360
rect 6546 2320 6552 2332
rect 6604 2320 6610 2372
rect 6822 2320 6828 2372
rect 6880 2360 6886 2372
rect 6880 2332 7236 2360
rect 6880 2320 6886 2332
rect 6917 2295 6975 2301
rect 6917 2292 6929 2295
rect 5543 2264 6929 2292
rect 5445 2255 5503 2261
rect 6917 2261 6929 2264
rect 6963 2261 6975 2295
rect 7208 2292 7236 2332
rect 7558 2320 7564 2372
rect 7616 2360 7622 2372
rect 8220 2360 8248 2391
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8812 2400 9137 2428
rect 8812 2388 8818 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2428 10379 2431
rect 10410 2428 10416 2440
rect 10367 2400 10416 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 7616 2332 8248 2360
rect 7616 2320 7622 2332
rect 7745 2295 7803 2301
rect 7745 2292 7757 2295
rect 7208 2264 7757 2292
rect 6917 2255 6975 2261
rect 7745 2261 7757 2264
rect 7791 2261 7803 2295
rect 8220 2292 8248 2332
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 10336 2360 10364 2391
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 8444 2332 10364 2360
rect 10796 2360 10824 2468
rect 11330 2456 11336 2468
rect 11388 2456 11394 2508
rect 11882 2456 11888 2508
rect 11940 2496 11946 2508
rect 12710 2496 12716 2508
rect 11940 2468 12716 2496
rect 11940 2456 11946 2468
rect 12710 2456 12716 2468
rect 12768 2456 12774 2508
rect 13078 2496 13084 2508
rect 13039 2468 13084 2496
rect 13078 2456 13084 2468
rect 13136 2456 13142 2508
rect 13354 2456 13360 2508
rect 13412 2496 13418 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 13412 2468 14841 2496
rect 13412 2456 13418 2468
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 14829 2459 14887 2465
rect 11609 2431 11667 2437
rect 11609 2397 11621 2431
rect 11655 2428 11667 2431
rect 11698 2428 11704 2440
rect 11655 2400 11704 2428
rect 11655 2397 11667 2400
rect 11609 2391 11667 2397
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 12986 2388 12992 2440
rect 13044 2428 13050 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 13044 2400 13185 2428
rect 13044 2388 13050 2400
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 14918 2428 14924 2440
rect 14507 2400 14924 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 12894 2360 12900 2372
rect 10796 2332 12900 2360
rect 8444 2320 8450 2332
rect 12894 2320 12900 2332
rect 12952 2320 12958 2372
rect 13538 2320 13544 2372
rect 13596 2320 13602 2372
rect 9490 2292 9496 2304
rect 8220 2264 9496 2292
rect 7745 2255 7803 2261
rect 9490 2252 9496 2264
rect 9548 2252 9554 2304
rect 9766 2292 9772 2304
rect 9727 2264 9772 2292
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 10134 2252 10140 2304
rect 10192 2292 10198 2304
rect 12434 2292 12440 2304
rect 10192 2264 12440 2292
rect 10192 2252 10198 2264
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 12618 2292 12624 2304
rect 12579 2264 12624 2292
rect 12618 2252 12624 2264
rect 12676 2252 12682 2304
rect 12710 2252 12716 2304
rect 12768 2292 12774 2304
rect 13556 2292 13584 2320
rect 15010 2292 15016 2304
rect 12768 2264 13584 2292
rect 14971 2264 15016 2292
rect 12768 2252 12774 2264
rect 15010 2252 15016 2264
rect 15068 2252 15074 2304
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 3142 2048 3148 2100
rect 3200 2088 3206 2100
rect 15010 2088 15016 2100
rect 3200 2060 15016 2088
rect 3200 2048 3206 2060
rect 15010 2048 15016 2060
rect 15068 2048 15074 2100
rect 2406 1980 2412 2032
rect 2464 2020 2470 2032
rect 12618 2020 12624 2032
rect 2464 1992 12624 2020
rect 2464 1980 2470 1992
rect 12618 1980 12624 1992
rect 12676 1980 12682 2032
rect 1578 1912 1584 1964
rect 1636 1952 1642 1964
rect 11330 1952 11336 1964
rect 1636 1924 11336 1952
rect 1636 1912 1642 1924
rect 11330 1912 11336 1924
rect 11388 1912 11394 1964
rect 12250 1912 12256 1964
rect 12308 1952 12314 1964
rect 14182 1952 14188 1964
rect 12308 1924 14188 1952
rect 12308 1912 12314 1924
rect 14182 1912 14188 1924
rect 14240 1912 14246 1964
rect 3878 1844 3884 1896
rect 3936 1884 3942 1896
rect 5994 1884 6000 1896
rect 3936 1856 6000 1884
rect 3936 1844 3942 1856
rect 5994 1844 6000 1856
rect 6052 1844 6058 1896
rect 6089 1887 6147 1893
rect 6089 1853 6101 1887
rect 6135 1884 6147 1887
rect 9766 1884 9772 1896
rect 6135 1856 9772 1884
rect 6135 1853 6147 1856
rect 6089 1847 6147 1853
rect 9766 1844 9772 1856
rect 9824 1844 9830 1896
rect 10318 1844 10324 1896
rect 10376 1884 10382 1896
rect 12342 1884 12348 1896
rect 10376 1856 12348 1884
rect 10376 1844 10382 1856
rect 12342 1844 12348 1856
rect 12400 1844 12406 1896
rect 5810 1776 5816 1828
rect 5868 1816 5874 1828
rect 6730 1816 6736 1828
rect 5868 1788 6736 1816
rect 5868 1776 5874 1788
rect 6730 1776 6736 1788
rect 6788 1776 6794 1828
rect 7190 1776 7196 1828
rect 7248 1816 7254 1828
rect 8662 1816 8668 1828
rect 7248 1788 8668 1816
rect 7248 1776 7254 1788
rect 8662 1776 8668 1788
rect 8720 1776 8726 1828
rect 11146 1776 11152 1828
rect 11204 1816 11210 1828
rect 15470 1816 15476 1828
rect 11204 1788 15476 1816
rect 11204 1776 11210 1788
rect 15470 1776 15476 1788
rect 15528 1776 15534 1828
rect 4062 1708 4068 1760
rect 4120 1748 4126 1760
rect 15102 1748 15108 1760
rect 4120 1720 15108 1748
rect 4120 1708 4126 1720
rect 15102 1708 15108 1720
rect 15160 1708 15166 1760
rect 4338 1640 4344 1692
rect 4396 1680 4402 1692
rect 8754 1680 8760 1692
rect 4396 1652 8760 1680
rect 4396 1640 4402 1652
rect 8754 1640 8760 1652
rect 8812 1640 8818 1692
rect 3786 1572 3792 1624
rect 3844 1612 3850 1624
rect 5902 1612 5908 1624
rect 3844 1584 5908 1612
rect 3844 1572 3850 1584
rect 5902 1572 5908 1584
rect 5960 1612 5966 1624
rect 9674 1612 9680 1624
rect 5960 1584 9680 1612
rect 5960 1572 5966 1584
rect 9674 1572 9680 1584
rect 9732 1572 9738 1624
rect 4154 1504 4160 1556
rect 4212 1544 4218 1556
rect 4890 1544 4896 1556
rect 4212 1516 4896 1544
rect 4212 1504 4218 1516
rect 4890 1504 4896 1516
rect 4948 1544 4954 1556
rect 11698 1544 11704 1556
rect 4948 1516 11704 1544
rect 4948 1504 4954 1516
rect 11698 1504 11704 1516
rect 11756 1504 11762 1556
rect 2130 1436 2136 1488
rect 2188 1476 2194 1488
rect 6089 1479 6147 1485
rect 6089 1476 6101 1479
rect 2188 1448 6101 1476
rect 2188 1436 2194 1448
rect 6089 1445 6101 1448
rect 6135 1445 6147 1479
rect 6089 1439 6147 1445
rect 6454 1436 6460 1488
rect 6512 1476 6518 1488
rect 11146 1476 11152 1488
rect 6512 1448 11152 1476
rect 6512 1436 6518 1448
rect 11146 1436 11152 1448
rect 11204 1436 11210 1488
rect 8110 1368 8116 1420
rect 8168 1408 8174 1420
rect 9490 1408 9496 1420
rect 8168 1380 9496 1408
rect 8168 1368 8174 1380
rect 9490 1368 9496 1380
rect 9548 1368 9554 1420
rect 6086 1300 6092 1352
rect 6144 1340 6150 1352
rect 8018 1340 8024 1352
rect 6144 1312 8024 1340
rect 6144 1300 6150 1312
rect 8018 1300 8024 1312
rect 8076 1300 8082 1352
rect 9122 824 9128 876
rect 9180 864 9186 876
rect 10594 864 10600 876
rect 9180 836 10600 864
rect 9180 824 9186 836
rect 10594 824 10600 836
rect 10652 824 10658 876
<< via1 >>
rect 1400 16464 1452 16516
rect 6644 16464 6696 16516
rect 2412 16396 2464 16448
rect 8208 16396 8260 16448
rect 1768 16328 1820 16380
rect 10324 16328 10376 16380
rect 4988 16260 5040 16312
rect 10140 16260 10192 16312
rect 11244 16260 11296 16312
rect 4068 16192 4120 16244
rect 8852 16192 8904 16244
rect 204 16124 256 16176
rect 13728 16124 13780 16176
rect 6368 16056 6420 16108
rect 12624 16056 12676 16108
rect 2780 15988 2832 16040
rect 6092 15988 6144 16040
rect 6920 15988 6972 16040
rect 9404 15988 9456 16040
rect 11336 15988 11388 16040
rect 3056 15920 3108 15972
rect 12900 15920 12952 15972
rect 572 15852 624 15904
rect 14464 15852 14516 15904
rect 5912 15750 5964 15802
rect 5976 15750 6028 15802
rect 6040 15750 6092 15802
rect 6104 15750 6156 15802
rect 10843 15750 10895 15802
rect 10907 15750 10959 15802
rect 10971 15750 11023 15802
rect 11035 15750 11087 15802
rect 2688 15648 2740 15700
rect 4160 15648 4212 15700
rect 6552 15648 6604 15700
rect 10324 15648 10376 15700
rect 13728 15691 13780 15700
rect 13728 15657 13737 15691
rect 13737 15657 13771 15691
rect 13771 15657 13780 15691
rect 13728 15648 13780 15657
rect 14464 15691 14516 15700
rect 14464 15657 14473 15691
rect 14473 15657 14507 15691
rect 14507 15657 14516 15691
rect 14464 15648 14516 15657
rect 4988 15580 5040 15632
rect 8300 15580 8352 15632
rect 2228 15512 2280 15564
rect 2872 15512 2924 15564
rect 4068 15512 4120 15564
rect 4712 15555 4764 15564
rect 4712 15521 4721 15555
rect 4721 15521 4755 15555
rect 4755 15521 4764 15555
rect 4712 15512 4764 15521
rect 7196 15512 7248 15564
rect 2136 15487 2188 15496
rect 2136 15453 2145 15487
rect 2145 15453 2179 15487
rect 2179 15453 2188 15487
rect 2136 15444 2188 15453
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 2780 15308 2832 15360
rect 6736 15444 6788 15496
rect 7656 15512 7708 15564
rect 8668 15580 8720 15632
rect 9588 15580 9640 15632
rect 12164 15580 12216 15632
rect 12900 15623 12952 15632
rect 8392 15444 8444 15496
rect 5540 15376 5592 15428
rect 9680 15512 9732 15564
rect 11980 15512 12032 15564
rect 12624 15555 12676 15564
rect 12624 15521 12633 15555
rect 12633 15521 12667 15555
rect 12667 15521 12676 15555
rect 12624 15512 12676 15521
rect 12900 15589 12909 15623
rect 12909 15589 12943 15623
rect 12943 15589 12952 15623
rect 12900 15580 12952 15589
rect 9312 15376 9364 15428
rect 13728 15444 13780 15496
rect 12256 15376 12308 15428
rect 4528 15308 4580 15360
rect 11244 15308 11296 15360
rect 13636 15308 13688 15360
rect 3447 15206 3499 15258
rect 3511 15206 3563 15258
rect 3575 15206 3627 15258
rect 3639 15206 3691 15258
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 13308 15206 13360 15258
rect 13372 15206 13424 15258
rect 13436 15206 13488 15258
rect 13500 15206 13552 15258
rect 2320 15104 2372 15156
rect 5172 15104 5224 15156
rect 5264 15104 5316 15156
rect 7380 15104 7432 15156
rect 8668 15104 8720 15156
rect 1860 15036 1912 15088
rect 5724 15036 5776 15088
rect 11152 15104 11204 15156
rect 15476 15104 15528 15156
rect 8944 15036 8996 15088
rect 13544 15036 13596 15088
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4068 14968 4120 14977
rect 4252 15011 4304 15020
rect 4252 14977 4261 15011
rect 4261 14977 4295 15011
rect 4295 14977 4304 15011
rect 4252 14968 4304 14977
rect 1492 14943 1544 14952
rect 1492 14909 1501 14943
rect 1501 14909 1535 14943
rect 1535 14909 1544 14943
rect 1492 14900 1544 14909
rect 4896 14968 4948 15020
rect 5448 15011 5500 15020
rect 5448 14977 5457 15011
rect 5457 14977 5491 15011
rect 5491 14977 5500 15011
rect 5448 14968 5500 14977
rect 7748 14968 7800 15020
rect 9220 15011 9272 15020
rect 9220 14977 9229 15011
rect 9229 14977 9263 15011
rect 9263 14977 9272 15011
rect 9220 14968 9272 14977
rect 11704 15011 11756 15020
rect 4804 14900 4856 14952
rect 5632 14832 5684 14884
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 3976 14807 4028 14816
rect 3976 14773 3985 14807
rect 3985 14773 4019 14807
rect 4019 14773 4028 14807
rect 3976 14764 4028 14773
rect 5724 14764 5776 14816
rect 7288 14900 7340 14952
rect 10324 14900 10376 14952
rect 10508 14900 10560 14952
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 12900 14968 12952 15020
rect 13084 15011 13136 15020
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13084 14968 13136 14977
rect 12348 14900 12400 14952
rect 12992 14900 13044 14952
rect 8760 14832 8812 14884
rect 11152 14832 11204 14884
rect 12072 14832 12124 14884
rect 14004 14900 14056 14952
rect 7380 14764 7432 14816
rect 9220 14764 9272 14816
rect 10692 14764 10744 14816
rect 11428 14764 11480 14816
rect 11796 14764 11848 14816
rect 12440 14807 12492 14816
rect 12440 14773 12449 14807
rect 12449 14773 12483 14807
rect 12483 14773 12492 14807
rect 12440 14764 12492 14773
rect 12624 14764 12676 14816
rect 15108 14832 15160 14884
rect 16304 14832 16356 14884
rect 14556 14807 14608 14816
rect 14556 14773 14565 14807
rect 14565 14773 14599 14807
rect 14599 14773 14608 14807
rect 14556 14764 14608 14773
rect 5912 14662 5964 14714
rect 5976 14662 6028 14714
rect 6040 14662 6092 14714
rect 6104 14662 6156 14714
rect 10843 14662 10895 14714
rect 10907 14662 10959 14714
rect 10971 14662 11023 14714
rect 11035 14662 11087 14714
rect 3332 14560 3384 14612
rect 3608 14560 3660 14612
rect 2136 14492 2188 14544
rect 2504 14467 2556 14476
rect 2504 14433 2513 14467
rect 2513 14433 2547 14467
rect 2547 14433 2556 14467
rect 2504 14424 2556 14433
rect 3884 14492 3936 14544
rect 5172 14560 5224 14612
rect 6368 14560 6420 14612
rect 7472 14560 7524 14612
rect 7656 14560 7708 14612
rect 7932 14560 7984 14612
rect 6460 14492 6512 14544
rect 7104 14492 7156 14544
rect 2964 14356 3016 14408
rect 3792 14424 3844 14476
rect 4252 14424 4304 14476
rect 8116 14492 8168 14544
rect 8852 14535 8904 14544
rect 8208 14424 8260 14476
rect 8852 14501 8861 14535
rect 8861 14501 8895 14535
rect 8895 14501 8904 14535
rect 8852 14492 8904 14501
rect 10048 14492 10100 14544
rect 9956 14467 10008 14476
rect 9956 14433 9990 14467
rect 9990 14433 10008 14467
rect 9956 14424 10008 14433
rect 10232 14424 10284 14476
rect 10508 14424 10560 14476
rect 11428 14560 11480 14612
rect 13084 14560 13136 14612
rect 11796 14492 11848 14544
rect 13544 14535 13596 14544
rect 12072 14424 12124 14476
rect 13268 14467 13320 14476
rect 13268 14433 13277 14467
rect 13277 14433 13311 14467
rect 13311 14433 13320 14467
rect 13268 14424 13320 14433
rect 13544 14501 13553 14535
rect 13553 14501 13587 14535
rect 13587 14501 13596 14535
rect 13544 14492 13596 14501
rect 16764 14424 16816 14476
rect 4344 14399 4396 14408
rect 4344 14365 4353 14399
rect 4353 14365 4387 14399
rect 4387 14365 4396 14399
rect 4344 14356 4396 14365
rect 5356 14356 5408 14408
rect 6736 14399 6788 14408
rect 6736 14365 6745 14399
rect 6745 14365 6779 14399
rect 6779 14365 6788 14399
rect 6736 14356 6788 14365
rect 8300 14356 8352 14408
rect 8484 14356 8536 14408
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 12716 14399 12768 14408
rect 12716 14365 12725 14399
rect 12725 14365 12759 14399
rect 12759 14365 12768 14399
rect 12716 14356 12768 14365
rect 12808 14356 12860 14408
rect 14096 14356 14148 14408
rect 6092 14288 6144 14340
rect 6184 14331 6236 14340
rect 6184 14297 6193 14331
rect 6193 14297 6227 14331
rect 6227 14297 6236 14331
rect 6184 14288 6236 14297
rect 3332 14220 3384 14272
rect 6552 14220 6604 14272
rect 9220 14288 9272 14340
rect 11980 14288 12032 14340
rect 10692 14220 10744 14272
rect 11336 14220 11388 14272
rect 11428 14220 11480 14272
rect 12808 14220 12860 14272
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 3447 14118 3499 14170
rect 3511 14118 3563 14170
rect 3575 14118 3627 14170
rect 3639 14118 3691 14170
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 13308 14118 13360 14170
rect 13372 14118 13424 14170
rect 13436 14118 13488 14170
rect 13500 14118 13552 14170
rect 2412 14016 2464 14068
rect 3792 14016 3844 14068
rect 5632 14016 5684 14068
rect 6368 14016 6420 14068
rect 6920 14016 6972 14068
rect 7564 14016 7616 14068
rect 7656 14016 7708 14068
rect 10508 14016 10560 14068
rect 3056 13948 3108 14000
rect 5172 13948 5224 14000
rect 6828 13948 6880 14000
rect 7472 13948 7524 14000
rect 8024 13948 8076 14000
rect 9864 13991 9916 14000
rect 1676 13812 1728 13864
rect 4620 13880 4672 13932
rect 4804 13923 4856 13932
rect 4804 13889 4813 13923
rect 4813 13889 4847 13923
rect 4847 13889 4856 13923
rect 4804 13880 4856 13889
rect 5540 13880 5592 13932
rect 5908 13923 5960 13932
rect 5908 13889 5917 13923
rect 5917 13889 5951 13923
rect 5951 13889 5960 13923
rect 5908 13880 5960 13889
rect 7196 13880 7248 13932
rect 3332 13812 3384 13864
rect 4528 13787 4580 13796
rect 4528 13753 4537 13787
rect 4537 13753 4571 13787
rect 4571 13753 4580 13787
rect 4528 13744 4580 13753
rect 6184 13812 6236 13864
rect 6644 13812 6696 13864
rect 7564 13812 7616 13864
rect 7748 13880 7800 13932
rect 7840 13812 7892 13864
rect 9864 13957 9873 13991
rect 9873 13957 9907 13991
rect 9907 13957 9916 13991
rect 9864 13948 9916 13957
rect 12716 13948 12768 14000
rect 9772 13880 9824 13932
rect 11244 13880 11296 13932
rect 13176 13880 13228 13932
rect 15016 13991 15068 14000
rect 15016 13957 15025 13991
rect 15025 13957 15059 13991
rect 15059 13957 15068 13991
rect 15016 13948 15068 13957
rect 8208 13744 8260 13796
rect 2872 13676 2924 13728
rect 3424 13676 3476 13728
rect 7564 13676 7616 13728
rect 7748 13719 7800 13728
rect 7748 13685 7757 13719
rect 7757 13685 7791 13719
rect 7791 13685 7800 13719
rect 7748 13676 7800 13685
rect 8300 13676 8352 13728
rect 8852 13744 8904 13796
rect 9128 13744 9180 13796
rect 14004 13787 14056 13796
rect 14004 13753 14013 13787
rect 14013 13753 14047 13787
rect 14047 13753 14056 13787
rect 14004 13744 14056 13753
rect 9036 13676 9088 13728
rect 11244 13676 11296 13728
rect 11888 13676 11940 13728
rect 12256 13676 12308 13728
rect 12716 13676 12768 13728
rect 5912 13574 5964 13626
rect 5976 13574 6028 13626
rect 6040 13574 6092 13626
rect 6104 13574 6156 13626
rect 10843 13574 10895 13626
rect 10907 13574 10959 13626
rect 10971 13574 11023 13626
rect 11035 13574 11087 13626
rect 1584 13472 1636 13524
rect 5540 13472 5592 13524
rect 5724 13472 5776 13524
rect 2136 13379 2188 13388
rect 2136 13345 2145 13379
rect 2145 13345 2179 13379
rect 2179 13345 2188 13379
rect 2136 13336 2188 13345
rect 2872 13336 2924 13388
rect 3148 13404 3200 13456
rect 4620 13404 4672 13456
rect 5264 13447 5316 13456
rect 5264 13413 5298 13447
rect 5298 13413 5316 13447
rect 5264 13404 5316 13413
rect 5632 13404 5684 13456
rect 9128 13472 9180 13524
rect 9496 13472 9548 13524
rect 12532 13472 12584 13524
rect 13084 13472 13136 13524
rect 14096 13472 14148 13524
rect 14740 13472 14792 13524
rect 7012 13336 7064 13388
rect 7196 13379 7248 13388
rect 7196 13345 7205 13379
rect 7205 13345 7239 13379
rect 7239 13345 7248 13379
rect 7196 13336 7248 13345
rect 7748 13336 7800 13388
rect 8668 13404 8720 13456
rect 9036 13404 9088 13456
rect 9680 13404 9732 13456
rect 9864 13404 9916 13456
rect 11612 13404 11664 13456
rect 13268 13404 13320 13456
rect 13728 13404 13780 13456
rect 10508 13336 10560 13388
rect 11704 13336 11756 13388
rect 12808 13336 12860 13388
rect 14832 13336 14884 13388
rect 4160 13200 4212 13252
rect 3332 13132 3384 13184
rect 4436 13268 4488 13320
rect 7380 13268 7432 13320
rect 6092 13132 6144 13184
rect 6460 13132 6512 13184
rect 7196 13132 7248 13184
rect 7932 13268 7984 13320
rect 8392 13268 8444 13320
rect 8852 13268 8904 13320
rect 7748 13200 7800 13252
rect 8024 13175 8076 13184
rect 8024 13141 8033 13175
rect 8033 13141 8067 13175
rect 8067 13141 8076 13175
rect 8024 13132 8076 13141
rect 8208 13200 8260 13252
rect 9128 13200 9180 13252
rect 9864 13268 9916 13320
rect 10232 13200 10284 13252
rect 9864 13132 9916 13184
rect 11428 13268 11480 13320
rect 12256 13268 12308 13320
rect 11980 13200 12032 13252
rect 12900 13200 12952 13252
rect 14004 13132 14056 13184
rect 3447 13030 3499 13082
rect 3511 13030 3563 13082
rect 3575 13030 3627 13082
rect 3639 13030 3691 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 13308 13030 13360 13082
rect 13372 13030 13424 13082
rect 13436 13030 13488 13082
rect 13500 13030 13552 13082
rect 5356 12928 5408 12980
rect 5448 12928 5500 12980
rect 2136 12860 2188 12912
rect 2320 12860 2372 12912
rect 4804 12860 4856 12912
rect 5264 12860 5316 12912
rect 6736 12860 6788 12912
rect 7012 12928 7064 12980
rect 7840 12928 7892 12980
rect 7932 12928 7984 12980
rect 8760 12928 8812 12980
rect 9036 12928 9088 12980
rect 9956 12928 10008 12980
rect 3608 12792 3660 12844
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 4436 12792 4488 12844
rect 4620 12792 4672 12844
rect 5080 12792 5132 12844
rect 5908 12792 5960 12844
rect 6092 12835 6144 12844
rect 6092 12801 6101 12835
rect 6101 12801 6135 12835
rect 6135 12801 6144 12835
rect 6092 12792 6144 12801
rect 2412 12724 2464 12776
rect 2688 12724 2740 12776
rect 7932 12792 7984 12844
rect 8392 12792 8444 12844
rect 8852 12792 8904 12844
rect 9312 12792 9364 12844
rect 10048 12792 10100 12844
rect 11336 12835 11388 12844
rect 11336 12801 11345 12835
rect 11345 12801 11379 12835
rect 11379 12801 11388 12835
rect 11336 12792 11388 12801
rect 11612 12928 11664 12980
rect 11520 12860 11572 12912
rect 12532 12860 12584 12912
rect 14188 12835 14240 12844
rect 14188 12801 14197 12835
rect 14197 12801 14231 12835
rect 14231 12801 14240 12835
rect 14188 12792 14240 12801
rect 3792 12656 3844 12708
rect 3976 12656 4028 12708
rect 4160 12656 4212 12708
rect 5448 12656 5500 12708
rect 7288 12724 7340 12776
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 8760 12724 8812 12776
rect 7012 12656 7064 12708
rect 7564 12656 7616 12708
rect 9036 12656 9088 12708
rect 9496 12656 9548 12708
rect 10508 12724 10560 12776
rect 11244 12724 11296 12776
rect 12532 12724 12584 12776
rect 13912 12724 13964 12776
rect 14832 12767 14884 12776
rect 14832 12733 14841 12767
rect 14841 12733 14875 12767
rect 14875 12733 14884 12767
rect 14832 12724 14884 12733
rect 15108 12724 15160 12776
rect 11520 12656 11572 12708
rect 13636 12656 13688 12708
rect 2412 12631 2464 12640
rect 2412 12597 2421 12631
rect 2421 12597 2455 12631
rect 2455 12597 2464 12631
rect 2412 12588 2464 12597
rect 3056 12588 3108 12640
rect 4344 12631 4396 12640
rect 4344 12597 4353 12631
rect 4353 12597 4387 12631
rect 4387 12597 4396 12631
rect 4344 12588 4396 12597
rect 4436 12588 4488 12640
rect 5816 12588 5868 12640
rect 7748 12631 7800 12640
rect 7748 12597 7757 12631
rect 7757 12597 7791 12631
rect 7791 12597 7800 12631
rect 7748 12588 7800 12597
rect 7932 12588 7984 12640
rect 8944 12588 8996 12640
rect 10048 12588 10100 12640
rect 10416 12588 10468 12640
rect 12164 12588 12216 12640
rect 13912 12588 13964 12640
rect 5912 12486 5964 12538
rect 5976 12486 6028 12538
rect 6040 12486 6092 12538
rect 6104 12486 6156 12538
rect 10843 12486 10895 12538
rect 10907 12486 10959 12538
rect 10971 12486 11023 12538
rect 11035 12486 11087 12538
rect 2044 12384 2096 12436
rect 3148 12427 3200 12436
rect 3148 12393 3157 12427
rect 3157 12393 3191 12427
rect 3191 12393 3200 12427
rect 3148 12384 3200 12393
rect 3240 12427 3292 12436
rect 3240 12393 3249 12427
rect 3249 12393 3283 12427
rect 3283 12393 3292 12427
rect 3240 12384 3292 12393
rect 2780 12248 2832 12300
rect 3056 12248 3108 12300
rect 4436 12248 4488 12300
rect 4712 12291 4764 12300
rect 4712 12257 4721 12291
rect 4721 12257 4755 12291
rect 4755 12257 4764 12291
rect 4712 12248 4764 12257
rect 5264 12248 5316 12300
rect 6644 12316 6696 12368
rect 7472 12384 7524 12436
rect 7564 12384 7616 12436
rect 8024 12384 8076 12436
rect 6920 12316 6972 12368
rect 6000 12180 6052 12232
rect 8392 12248 8444 12300
rect 3056 12112 3108 12164
rect 3240 12112 3292 12164
rect 4344 12112 4396 12164
rect 4712 12112 4764 12164
rect 5724 12112 5776 12164
rect 6184 12112 6236 12164
rect 4160 12044 4212 12096
rect 4620 12044 4672 12096
rect 5448 12044 5500 12096
rect 6092 12087 6144 12096
rect 6092 12053 6101 12087
rect 6101 12053 6135 12087
rect 6135 12053 6144 12087
rect 6092 12044 6144 12053
rect 7564 12180 7616 12232
rect 8760 12180 8812 12232
rect 11336 12384 11388 12436
rect 11428 12384 11480 12436
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 8392 12155 8444 12164
rect 8392 12121 8401 12155
rect 8401 12121 8435 12155
rect 8435 12121 8444 12155
rect 8392 12112 8444 12121
rect 8668 12112 8720 12164
rect 14648 12316 14700 12368
rect 7288 12044 7340 12096
rect 8852 12044 8904 12096
rect 9772 12248 9824 12300
rect 9680 12223 9732 12232
rect 9680 12189 9689 12223
rect 9689 12189 9723 12223
rect 9723 12189 9732 12223
rect 9680 12180 9732 12189
rect 10968 12180 11020 12232
rect 9312 12044 9364 12096
rect 9680 12044 9732 12096
rect 10692 12044 10744 12096
rect 11244 12112 11296 12164
rect 11612 12180 11664 12232
rect 12256 12248 12308 12300
rect 13268 12291 13320 12300
rect 12532 12223 12584 12232
rect 12532 12189 12541 12223
rect 12541 12189 12575 12223
rect 12575 12189 12584 12223
rect 12532 12180 12584 12189
rect 13268 12257 13277 12291
rect 13277 12257 13311 12291
rect 13311 12257 13320 12291
rect 13268 12248 13320 12257
rect 14188 12291 14240 12300
rect 14188 12257 14197 12291
rect 14197 12257 14231 12291
rect 14231 12257 14240 12291
rect 14188 12248 14240 12257
rect 13452 12223 13504 12232
rect 13452 12189 13461 12223
rect 13461 12189 13495 12223
rect 13495 12189 13504 12223
rect 13452 12180 13504 12189
rect 13544 12180 13596 12232
rect 10876 12044 10928 12096
rect 12072 12044 12124 12096
rect 13084 12044 13136 12096
rect 3447 11942 3499 11994
rect 3511 11942 3563 11994
rect 3575 11942 3627 11994
rect 3639 11942 3691 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 13308 11942 13360 11994
rect 13372 11942 13424 11994
rect 13436 11942 13488 11994
rect 13500 11942 13552 11994
rect 1860 11883 1912 11892
rect 1860 11849 1869 11883
rect 1869 11849 1903 11883
rect 1903 11849 1912 11883
rect 1860 11840 1912 11849
rect 2044 11840 2096 11892
rect 6000 11840 6052 11892
rect 6092 11840 6144 11892
rect 8944 11840 8996 11892
rect 9220 11840 9272 11892
rect 10324 11840 10376 11892
rect 11612 11840 11664 11892
rect 2320 11772 2372 11824
rect 6184 11772 6236 11824
rect 6828 11772 6880 11824
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 2228 11636 2280 11645
rect 2688 11636 2740 11688
rect 4896 11679 4948 11688
rect 4896 11645 4905 11679
rect 4905 11645 4939 11679
rect 4939 11645 4948 11679
rect 4896 11636 4948 11645
rect 5908 11704 5960 11756
rect 6644 11704 6696 11756
rect 6276 11636 6328 11688
rect 2412 11568 2464 11620
rect 3148 11568 3200 11620
rect 3424 11568 3476 11620
rect 5264 11568 5316 11620
rect 6736 11568 6788 11620
rect 7472 11636 7524 11688
rect 10876 11772 10928 11824
rect 11152 11772 11204 11824
rect 11520 11772 11572 11824
rect 13820 11772 13872 11824
rect 8484 11704 8536 11756
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 8852 11636 8904 11688
rect 6920 11568 6972 11620
rect 9312 11704 9364 11756
rect 11060 11704 11112 11756
rect 11612 11704 11664 11756
rect 9680 11636 9732 11688
rect 10968 11636 11020 11688
rect 11152 11636 11204 11688
rect 3792 11500 3844 11552
rect 10324 11568 10376 11620
rect 11336 11568 11388 11620
rect 13176 11636 13228 11688
rect 14464 11636 14516 11688
rect 15936 11636 15988 11688
rect 8208 11500 8260 11552
rect 8944 11500 8996 11552
rect 9680 11500 9732 11552
rect 9956 11500 10008 11552
rect 12532 11568 12584 11620
rect 12716 11568 12768 11620
rect 13268 11568 13320 11620
rect 12440 11543 12492 11552
rect 12440 11509 12449 11543
rect 12449 11509 12483 11543
rect 12483 11509 12492 11543
rect 12900 11543 12952 11552
rect 12440 11500 12492 11509
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 13544 11500 13596 11552
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 6104 11398 6156 11450
rect 10843 11398 10895 11450
rect 10907 11398 10959 11450
rect 10971 11398 11023 11450
rect 11035 11398 11087 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 2688 11296 2740 11348
rect 2044 11271 2096 11280
rect 2044 11237 2053 11271
rect 2053 11237 2087 11271
rect 2087 11237 2096 11271
rect 2044 11228 2096 11237
rect 3056 11296 3108 11348
rect 4068 11296 4120 11348
rect 4344 11339 4396 11348
rect 4344 11305 4353 11339
rect 4353 11305 4387 11339
rect 4387 11305 4396 11339
rect 4344 11296 4396 11305
rect 6552 11296 6604 11348
rect 6736 11296 6788 11348
rect 7656 11271 7708 11280
rect 7656 11237 7668 11271
rect 7668 11237 7708 11271
rect 7656 11228 7708 11237
rect 8116 11296 8168 11348
rect 9220 11339 9272 11348
rect 8576 11228 8628 11280
rect 9220 11305 9229 11339
rect 9229 11305 9263 11339
rect 9263 11305 9272 11339
rect 9220 11296 9272 11305
rect 9680 11339 9732 11348
rect 9680 11305 9689 11339
rect 9689 11305 9723 11339
rect 9723 11305 9732 11339
rect 9680 11296 9732 11305
rect 11612 11296 11664 11348
rect 12716 11296 12768 11348
rect 13636 11296 13688 11348
rect 9312 11228 9364 11280
rect 10048 11271 10100 11280
rect 10048 11237 10057 11271
rect 10057 11237 10091 11271
rect 10091 11237 10100 11271
rect 10048 11228 10100 11237
rect 11520 11228 11572 11280
rect 14280 11228 14332 11280
rect 3056 11092 3108 11144
rect 3240 11135 3292 11144
rect 3240 11101 3249 11135
rect 3249 11101 3283 11135
rect 3283 11101 3292 11135
rect 3240 11092 3292 11101
rect 3332 11135 3384 11144
rect 3332 11101 3341 11135
rect 3341 11101 3375 11135
rect 3375 11101 3384 11135
rect 4160 11160 4212 11212
rect 5448 11160 5500 11212
rect 6552 11160 6604 11212
rect 6920 11160 6972 11212
rect 8484 11160 8536 11212
rect 9864 11160 9916 11212
rect 4988 11135 5040 11144
rect 3332 11092 3384 11101
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 5356 11092 5408 11144
rect 8668 11092 8720 11144
rect 1676 11024 1728 11076
rect 5080 11024 5132 11076
rect 6552 11024 6604 11076
rect 7104 11024 7156 11076
rect 8392 11024 8444 11076
rect 11336 11160 11388 11212
rect 12256 11160 12308 11212
rect 12808 11160 12860 11212
rect 13268 11160 13320 11212
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 13912 11160 13964 11212
rect 11980 11092 12032 11144
rect 12348 11092 12400 11144
rect 12624 11135 12676 11144
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 12624 11092 12676 11101
rect 3056 10956 3108 11008
rect 4896 10956 4948 11008
rect 5724 10956 5776 11008
rect 6736 10956 6788 11008
rect 6828 10956 6880 11008
rect 9772 11024 9824 11076
rect 11244 11024 11296 11076
rect 9220 10956 9272 11008
rect 13268 11067 13320 11076
rect 13268 11033 13277 11067
rect 13277 11033 13311 11067
rect 13311 11033 13320 11067
rect 13268 11024 13320 11033
rect 13912 11024 13964 11076
rect 15476 11160 15528 11212
rect 13084 10956 13136 11008
rect 3447 10854 3499 10906
rect 3511 10854 3563 10906
rect 3575 10854 3627 10906
rect 3639 10854 3691 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 13308 10854 13360 10906
rect 13372 10854 13424 10906
rect 13436 10854 13488 10906
rect 13500 10854 13552 10906
rect 2688 10752 2740 10804
rect 2688 10659 2740 10668
rect 2688 10625 2697 10659
rect 2697 10625 2731 10659
rect 2731 10625 2740 10659
rect 2688 10616 2740 10625
rect 2872 10659 2924 10668
rect 2872 10625 2881 10659
rect 2881 10625 2915 10659
rect 2915 10625 2924 10659
rect 2872 10616 2924 10625
rect 3792 10752 3844 10804
rect 3056 10659 3108 10668
rect 3056 10625 3065 10659
rect 3065 10625 3099 10659
rect 3099 10625 3108 10659
rect 3056 10616 3108 10625
rect 2412 10480 2464 10532
rect 3608 10548 3660 10600
rect 5908 10752 5960 10804
rect 6460 10752 6512 10804
rect 7564 10752 7616 10804
rect 8024 10752 8076 10804
rect 9956 10752 10008 10804
rect 10232 10752 10284 10804
rect 10692 10752 10744 10804
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 5724 10548 5776 10600
rect 6460 10548 6512 10600
rect 4712 10480 4764 10532
rect 8116 10616 8168 10668
rect 6920 10548 6972 10600
rect 7104 10591 7156 10600
rect 7104 10557 7138 10591
rect 7138 10557 7156 10591
rect 7104 10548 7156 10557
rect 7656 10548 7708 10600
rect 9680 10684 9732 10736
rect 12992 10752 13044 10804
rect 11152 10684 11204 10736
rect 9864 10616 9916 10668
rect 10784 10616 10836 10668
rect 11520 10616 11572 10668
rect 12072 10684 12124 10736
rect 12624 10616 12676 10668
rect 3056 10412 3108 10464
rect 6276 10412 6328 10464
rect 7840 10480 7892 10532
rect 8024 10480 8076 10532
rect 8668 10480 8720 10532
rect 9680 10480 9732 10532
rect 10140 10548 10192 10600
rect 10416 10548 10468 10600
rect 10784 10480 10836 10532
rect 14740 10659 14792 10668
rect 14740 10625 14749 10659
rect 14749 10625 14783 10659
rect 14783 10625 14792 10659
rect 14740 10616 14792 10625
rect 13268 10548 13320 10600
rect 12072 10480 12124 10532
rect 12992 10480 13044 10532
rect 13728 10548 13780 10600
rect 13912 10523 13964 10532
rect 13912 10489 13921 10523
rect 13921 10489 13955 10523
rect 13955 10489 13964 10523
rect 13912 10480 13964 10489
rect 8300 10412 8352 10464
rect 11428 10412 11480 10464
rect 11980 10412 12032 10464
rect 12256 10412 12308 10464
rect 12348 10412 12400 10464
rect 15200 10412 15252 10464
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 6104 10310 6156 10362
rect 10843 10310 10895 10362
rect 10907 10310 10959 10362
rect 10971 10310 11023 10362
rect 11035 10310 11087 10362
rect 2688 10208 2740 10260
rect 4528 10140 4580 10192
rect 5724 10140 5776 10192
rect 5816 10140 5868 10192
rect 2780 10072 2832 10124
rect 1860 10004 1912 10056
rect 3056 10072 3108 10124
rect 3424 10072 3476 10124
rect 3148 10004 3200 10056
rect 5540 10072 5592 10124
rect 7196 10208 7248 10260
rect 7656 10208 7708 10260
rect 7932 10208 7984 10260
rect 8392 10208 8444 10260
rect 8668 10208 8720 10260
rect 9220 10208 9272 10260
rect 6276 10140 6328 10192
rect 9772 10140 9824 10192
rect 10324 10140 10376 10192
rect 10508 10208 10560 10260
rect 11980 10208 12032 10260
rect 12624 10140 12676 10192
rect 12808 10140 12860 10192
rect 8116 10072 8168 10124
rect 8300 10072 8352 10124
rect 8392 10072 8444 10124
rect 10048 10115 10100 10124
rect 10048 10081 10057 10115
rect 10057 10081 10091 10115
rect 10091 10081 10100 10115
rect 10048 10072 10100 10081
rect 2320 9911 2372 9920
rect 2320 9877 2329 9911
rect 2329 9877 2363 9911
rect 2363 9877 2372 9911
rect 2320 9868 2372 9877
rect 2412 9868 2464 9920
rect 2964 9868 3016 9920
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 4436 10004 4488 10056
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 5448 10004 5500 10056
rect 6920 10004 6972 10056
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 9680 10004 9732 10056
rect 10508 10072 10560 10124
rect 10692 10072 10744 10124
rect 11152 10004 11204 10056
rect 11428 10004 11480 10056
rect 12900 10072 12952 10124
rect 13176 10140 13228 10192
rect 13544 10072 13596 10124
rect 14280 10072 14332 10124
rect 14740 10072 14792 10124
rect 12532 10047 12584 10056
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 5632 9936 5684 9988
rect 8944 9936 8996 9988
rect 10600 9936 10652 9988
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 13728 10004 13780 10013
rect 13084 9936 13136 9988
rect 14648 9979 14700 9988
rect 14648 9945 14657 9979
rect 14657 9945 14691 9979
rect 14691 9945 14700 9979
rect 14648 9936 14700 9945
rect 6092 9868 6144 9920
rect 6736 9868 6788 9920
rect 10048 9868 10100 9920
rect 12900 9868 12952 9920
rect 3447 9766 3499 9818
rect 3511 9766 3563 9818
rect 3575 9766 3627 9818
rect 3639 9766 3691 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 13308 9766 13360 9818
rect 13372 9766 13424 9818
rect 13436 9766 13488 9818
rect 13500 9766 13552 9818
rect 1492 9664 1544 9716
rect 3056 9664 3108 9716
rect 3608 9596 3660 9648
rect 3148 9460 3200 9512
rect 1952 9435 2004 9444
rect 1952 9401 1961 9435
rect 1961 9401 1995 9435
rect 1995 9401 2004 9435
rect 1952 9392 2004 9401
rect 2688 9392 2740 9444
rect 3700 9528 3752 9580
rect 5448 9664 5500 9716
rect 5540 9664 5592 9716
rect 11428 9664 11480 9716
rect 14648 9664 14700 9716
rect 6552 9596 6604 9648
rect 7932 9596 7984 9648
rect 8300 9596 8352 9648
rect 8576 9596 8628 9648
rect 9680 9596 9732 9648
rect 11152 9596 11204 9648
rect 7840 9528 7892 9580
rect 10232 9528 10284 9580
rect 10600 9528 10652 9580
rect 12808 9596 12860 9648
rect 4059 9503 4111 9512
rect 4059 9469 4091 9503
rect 4091 9469 4111 9503
rect 4059 9460 4111 9469
rect 5080 9460 5132 9512
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 3148 9367 3200 9376
rect 3148 9333 3157 9367
rect 3157 9333 3191 9367
rect 3191 9333 3200 9367
rect 3148 9324 3200 9333
rect 3792 9324 3844 9376
rect 5540 9435 5592 9444
rect 5540 9401 5574 9435
rect 5574 9401 5592 9435
rect 6920 9460 6972 9512
rect 8576 9460 8628 9512
rect 8668 9460 8720 9512
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 10048 9460 10100 9512
rect 12624 9528 12676 9580
rect 13636 9596 13688 9648
rect 14280 9596 14332 9648
rect 14832 9596 14884 9648
rect 15016 9639 15068 9648
rect 15016 9605 15025 9639
rect 15025 9605 15059 9639
rect 15059 9605 15068 9639
rect 15016 9596 15068 9605
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 13360 9528 13412 9580
rect 5540 9392 5592 9401
rect 9772 9392 9824 9444
rect 12164 9460 12216 9512
rect 13912 9460 13964 9512
rect 14648 9460 14700 9512
rect 11888 9392 11940 9444
rect 6736 9324 6788 9376
rect 7840 9324 7892 9376
rect 9680 9324 9732 9376
rect 10416 9324 10468 9376
rect 10600 9324 10652 9376
rect 11428 9367 11480 9376
rect 11428 9333 11437 9367
rect 11437 9333 11471 9367
rect 11471 9333 11480 9367
rect 11428 9324 11480 9333
rect 13268 9324 13320 9376
rect 13636 9367 13688 9376
rect 13636 9333 13645 9367
rect 13645 9333 13679 9367
rect 13679 9333 13688 9367
rect 13636 9324 13688 9333
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 6104 9222 6156 9274
rect 10843 9222 10895 9274
rect 10907 9222 10959 9274
rect 10971 9222 11023 9274
rect 11035 9222 11087 9274
rect 4896 9120 4948 9172
rect 5080 9120 5132 9172
rect 11612 9120 11664 9172
rect 13728 9120 13780 9172
rect 1676 9095 1728 9104
rect 1676 9061 1685 9095
rect 1685 9061 1719 9095
rect 1719 9061 1728 9095
rect 1676 9052 1728 9061
rect 3056 9052 3108 9104
rect 6920 9052 6972 9104
rect 7012 9052 7064 9104
rect 8024 9052 8076 9104
rect 8300 9052 8352 9104
rect 9772 9052 9824 9104
rect 2320 8984 2372 9036
rect 2412 8959 2464 8968
rect 2412 8925 2421 8959
rect 2421 8925 2455 8959
rect 2455 8925 2464 8959
rect 2412 8916 2464 8925
rect 5632 8984 5684 9036
rect 5816 9027 5868 9036
rect 5816 8993 5825 9027
rect 5825 8993 5859 9027
rect 5859 8993 5868 9027
rect 5816 8984 5868 8993
rect 6276 8984 6328 9036
rect 4436 8916 4488 8968
rect 7104 8984 7156 9036
rect 7564 8984 7616 9036
rect 3056 8848 3108 8900
rect 4160 8848 4212 8900
rect 1952 8823 2004 8832
rect 1952 8789 1961 8823
rect 1961 8789 1995 8823
rect 1995 8789 2004 8823
rect 1952 8780 2004 8789
rect 2780 8823 2832 8832
rect 2780 8789 2789 8823
rect 2789 8789 2823 8823
rect 2823 8789 2832 8823
rect 2780 8780 2832 8789
rect 3792 8780 3844 8832
rect 4068 8780 4120 8832
rect 4896 8848 4948 8900
rect 6184 8848 6236 8900
rect 8760 8916 8812 8968
rect 7564 8848 7616 8900
rect 10508 8984 10560 9036
rect 11060 8984 11112 9036
rect 11152 8984 11204 9036
rect 11336 9027 11388 9036
rect 11336 8993 11345 9027
rect 11345 8993 11379 9027
rect 11379 8993 11388 9027
rect 11336 8984 11388 8993
rect 11704 9052 11756 9104
rect 12440 9095 12492 9104
rect 12440 9061 12449 9095
rect 12449 9061 12483 9095
rect 12483 9061 12492 9095
rect 12440 9052 12492 9061
rect 12072 8984 12124 9036
rect 12256 8984 12308 9036
rect 12348 8984 12400 9036
rect 13360 9052 13412 9104
rect 12808 8984 12860 9036
rect 14188 9027 14240 9036
rect 14188 8993 14197 9027
rect 14197 8993 14231 9027
rect 14231 8993 14240 9027
rect 14188 8984 14240 8993
rect 10416 8848 10468 8900
rect 11336 8848 11388 8900
rect 12992 8916 13044 8968
rect 15108 8916 15160 8968
rect 6828 8780 6880 8832
rect 6920 8780 6972 8832
rect 8024 8780 8076 8832
rect 8760 8780 8812 8832
rect 13084 8848 13136 8900
rect 13268 8848 13320 8900
rect 15292 8848 15344 8900
rect 12440 8780 12492 8832
rect 13176 8780 13228 8832
rect 3447 8678 3499 8730
rect 3511 8678 3563 8730
rect 3575 8678 3627 8730
rect 3639 8678 3691 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 13308 8678 13360 8730
rect 13372 8678 13424 8730
rect 13436 8678 13488 8730
rect 13500 8678 13552 8730
rect 2504 8576 2556 8628
rect 2688 8619 2740 8628
rect 2688 8585 2697 8619
rect 2697 8585 2731 8619
rect 2731 8585 2740 8619
rect 2688 8576 2740 8585
rect 3148 8576 3200 8628
rect 4436 8576 4488 8628
rect 6276 8619 6328 8628
rect 6276 8585 6285 8619
rect 6285 8585 6319 8619
rect 6319 8585 6328 8619
rect 6276 8576 6328 8585
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 3332 8440 3384 8492
rect 4528 8483 4580 8492
rect 4528 8449 4537 8483
rect 4537 8449 4571 8483
rect 4571 8449 4580 8483
rect 4528 8440 4580 8449
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 2320 8372 2372 8424
rect 2964 8372 3016 8424
rect 4896 8415 4948 8424
rect 4896 8381 4905 8415
rect 4905 8381 4939 8415
rect 4939 8381 4948 8415
rect 4896 8372 4948 8381
rect 4344 8304 4396 8356
rect 5540 8372 5592 8424
rect 7104 8576 7156 8628
rect 7564 8576 7616 8628
rect 10416 8576 10468 8628
rect 10600 8576 10652 8628
rect 11428 8576 11480 8628
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 8300 8508 8352 8560
rect 7932 8440 7984 8492
rect 5632 8304 5684 8356
rect 6736 8304 6788 8356
rect 6920 8372 6972 8424
rect 8484 8372 8536 8424
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 10968 8508 11020 8560
rect 11980 8508 12032 8560
rect 10784 8440 10836 8492
rect 11612 8440 11664 8492
rect 14464 8576 14516 8628
rect 14280 8508 14332 8560
rect 10048 8372 10100 8424
rect 13452 8440 13504 8492
rect 13728 8440 13780 8492
rect 14372 8372 14424 8424
rect 14740 8372 14792 8424
rect 2320 8279 2372 8288
rect 2320 8245 2329 8279
rect 2329 8245 2363 8279
rect 2363 8245 2372 8279
rect 2320 8236 2372 8245
rect 2964 8236 3016 8288
rect 3424 8236 3476 8288
rect 4620 8236 4672 8288
rect 4896 8236 4948 8288
rect 7840 8236 7892 8288
rect 8208 8304 8260 8356
rect 9588 8236 9640 8288
rect 10416 8304 10468 8356
rect 11060 8304 11112 8356
rect 10692 8236 10744 8288
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 13452 8236 13504 8288
rect 14464 8236 14516 8288
rect 14648 8236 14700 8288
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 6104 8134 6156 8186
rect 10843 8134 10895 8186
rect 10907 8134 10959 8186
rect 10971 8134 11023 8186
rect 11035 8134 11087 8186
rect 2320 8032 2372 8084
rect 2780 8032 2832 8084
rect 6552 8032 6604 8084
rect 6736 8032 6788 8084
rect 9772 8032 9824 8084
rect 10232 8032 10284 8084
rect 10600 8032 10652 8084
rect 2504 7964 2556 8016
rect 2044 7939 2096 7948
rect 2044 7905 2053 7939
rect 2053 7905 2087 7939
rect 2087 7905 2096 7939
rect 2044 7896 2096 7905
rect 2780 7939 2832 7948
rect 2780 7905 2789 7939
rect 2789 7905 2823 7939
rect 2823 7905 2832 7939
rect 2780 7896 2832 7905
rect 2964 7896 3016 7948
rect 3424 7896 3476 7948
rect 2688 7828 2740 7880
rect 3148 7828 3200 7880
rect 3792 7939 3844 7948
rect 3792 7905 3801 7939
rect 3801 7905 3835 7939
rect 3835 7905 3844 7939
rect 3792 7896 3844 7905
rect 5080 7896 5132 7948
rect 4344 7828 4396 7880
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 5264 7828 5316 7880
rect 7012 7964 7064 8016
rect 7288 7964 7340 8016
rect 7564 7964 7616 8016
rect 7840 7964 7892 8016
rect 8576 7964 8628 8016
rect 5632 7939 5684 7948
rect 5632 7905 5641 7939
rect 5641 7905 5675 7939
rect 5675 7905 5684 7939
rect 5632 7896 5684 7905
rect 5448 7760 5500 7812
rect 3332 7692 3384 7744
rect 3976 7692 4028 7744
rect 5264 7735 5316 7744
rect 5264 7701 5273 7735
rect 5273 7701 5307 7735
rect 5307 7701 5316 7735
rect 5264 7692 5316 7701
rect 6736 7828 6788 7880
rect 9588 7896 9640 7948
rect 10508 7896 10560 7948
rect 11152 8032 11204 8084
rect 11612 8032 11664 8084
rect 12348 8032 12400 8084
rect 13176 8032 13228 8084
rect 14280 8075 14332 8084
rect 14280 8041 14289 8075
rect 14289 8041 14323 8075
rect 14323 8041 14332 8075
rect 14280 8032 14332 8041
rect 11980 8007 12032 8016
rect 11980 7973 11989 8007
rect 11989 7973 12023 8007
rect 12023 7973 12032 8007
rect 11980 7964 12032 7973
rect 11888 7896 11940 7948
rect 12532 7896 12584 7948
rect 8576 7828 8628 7880
rect 6920 7692 6972 7744
rect 8760 7692 8812 7744
rect 8944 7692 8996 7744
rect 9496 7760 9548 7812
rect 10692 7828 10744 7880
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 13636 7828 13688 7880
rect 15384 7828 15436 7880
rect 11152 7692 11204 7744
rect 11612 7692 11664 7744
rect 13912 7735 13964 7744
rect 13912 7701 13921 7735
rect 13921 7701 13955 7735
rect 13955 7701 13964 7735
rect 13912 7692 13964 7701
rect 14004 7692 14056 7744
rect 14372 7692 14424 7744
rect 3447 7590 3499 7642
rect 3511 7590 3563 7642
rect 3575 7590 3627 7642
rect 3639 7590 3691 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 13308 7590 13360 7642
rect 13372 7590 13424 7642
rect 13436 7590 13488 7642
rect 13500 7590 13552 7642
rect 2964 7420 3016 7472
rect 1492 7352 1544 7404
rect 1676 7352 1728 7404
rect 2504 7352 2556 7404
rect 6000 7488 6052 7540
rect 6276 7531 6328 7540
rect 6276 7497 6285 7531
rect 6285 7497 6319 7531
rect 6319 7497 6328 7531
rect 6276 7488 6328 7497
rect 6828 7488 6880 7540
rect 4344 7420 4396 7472
rect 5908 7420 5960 7472
rect 6184 7420 6236 7472
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 6828 7395 6880 7404
rect 1768 7284 1820 7336
rect 2228 7284 2280 7336
rect 2412 7284 2464 7336
rect 2780 7216 2832 7268
rect 3148 7216 3200 7268
rect 6000 7284 6052 7336
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 11060 7488 11112 7540
rect 12992 7488 13044 7540
rect 13176 7488 13228 7540
rect 14740 7488 14792 7540
rect 14924 7488 14976 7540
rect 9680 7420 9732 7472
rect 13268 7420 13320 7472
rect 10232 7352 10284 7404
rect 10508 7352 10560 7404
rect 10692 7352 10744 7404
rect 12072 7352 12124 7404
rect 12440 7352 12492 7404
rect 12624 7352 12676 7404
rect 13360 7352 13412 7404
rect 14464 7352 14516 7404
rect 14556 7352 14608 7404
rect 5172 7259 5224 7268
rect 5172 7225 5206 7259
rect 5206 7225 5224 7259
rect 5172 7216 5224 7225
rect 5448 7216 5500 7268
rect 7472 7284 7524 7336
rect 7932 7284 7984 7336
rect 8024 7284 8076 7336
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 9496 7284 9548 7336
rect 10048 7284 10100 7336
rect 10416 7284 10468 7336
rect 11612 7284 11664 7336
rect 7104 7259 7156 7268
rect 1584 7148 1636 7200
rect 1768 7191 1820 7200
rect 1768 7157 1777 7191
rect 1777 7157 1811 7191
rect 1811 7157 1820 7191
rect 1768 7148 1820 7157
rect 4068 7148 4120 7200
rect 4712 7148 4764 7200
rect 5356 7148 5408 7200
rect 6276 7148 6328 7200
rect 7104 7225 7138 7259
rect 7138 7225 7156 7259
rect 7104 7216 7156 7225
rect 7288 7148 7340 7200
rect 7472 7148 7524 7200
rect 8116 7148 8168 7200
rect 11152 7216 11204 7268
rect 12716 7284 12768 7336
rect 12900 7284 12952 7336
rect 13176 7284 13228 7336
rect 9772 7148 9824 7200
rect 10140 7148 10192 7200
rect 10416 7148 10468 7200
rect 12256 7148 12308 7200
rect 14096 7216 14148 7268
rect 14556 7216 14608 7268
rect 13268 7148 13320 7200
rect 15936 7148 15988 7200
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 6104 7046 6156 7098
rect 10843 7046 10895 7098
rect 10907 7046 10959 7098
rect 10971 7046 11023 7098
rect 11035 7046 11087 7098
rect 1768 6944 1820 6996
rect 2320 6944 2372 6996
rect 3056 6944 3108 6996
rect 4436 6987 4488 6996
rect 4436 6953 4445 6987
rect 4445 6953 4479 6987
rect 4479 6953 4488 6987
rect 4436 6944 4488 6953
rect 5172 6944 5224 6996
rect 9772 6944 9824 6996
rect 10600 6944 10652 6996
rect 12624 6944 12676 6996
rect 1584 6876 1636 6928
rect 4620 6876 4672 6928
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 2688 6808 2740 6860
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 4436 6740 4488 6792
rect 5356 6876 5408 6928
rect 6828 6876 6880 6928
rect 6092 6808 6144 6860
rect 7656 6876 7708 6928
rect 8300 6876 8352 6928
rect 8944 6919 8996 6928
rect 8944 6885 8953 6919
rect 8953 6885 8987 6919
rect 8987 6885 8996 6919
rect 8944 6876 8996 6885
rect 9036 6919 9088 6928
rect 9036 6885 9045 6919
rect 9045 6885 9079 6919
rect 9079 6885 9088 6919
rect 9036 6876 9088 6885
rect 12440 6876 12492 6928
rect 4896 6740 4948 6792
rect 5172 6740 5224 6792
rect 6276 6740 6328 6792
rect 7932 6808 7984 6860
rect 9772 6808 9824 6860
rect 10416 6808 10468 6860
rect 11060 6808 11112 6860
rect 11152 6808 11204 6860
rect 8392 6740 8444 6792
rect 9220 6740 9272 6792
rect 9496 6740 9548 6792
rect 10692 6740 10744 6792
rect 12256 6808 12308 6860
rect 12808 6876 12860 6928
rect 15292 6876 15344 6928
rect 16304 6876 16356 6928
rect 12624 6808 12676 6860
rect 14280 6851 14332 6860
rect 2504 6604 2556 6656
rect 4528 6604 4580 6656
rect 6736 6604 6788 6656
rect 9588 6604 9640 6656
rect 11704 6672 11756 6724
rect 11428 6604 11480 6656
rect 12164 6740 12216 6792
rect 12992 6740 13044 6792
rect 13176 6783 13228 6792
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 14280 6817 14289 6851
rect 14289 6817 14323 6851
rect 14323 6817 14332 6851
rect 14280 6808 14332 6817
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 13820 6672 13872 6724
rect 12256 6604 12308 6656
rect 12532 6604 12584 6656
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 2136 6400 2188 6452
rect 3792 6400 3844 6452
rect 4068 6400 4120 6452
rect 2412 6332 2464 6384
rect 1860 6264 1912 6316
rect 2412 6196 2464 6248
rect 4896 6307 4948 6316
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 4160 6196 4212 6248
rect 5448 6196 5500 6248
rect 5632 6196 5684 6248
rect 9588 6400 9640 6452
rect 7656 6332 7708 6384
rect 9128 6332 9180 6384
rect 9312 6332 9364 6384
rect 6552 6264 6604 6316
rect 7472 6307 7524 6316
rect 6092 6196 6144 6248
rect 7196 6196 7248 6248
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 9036 6264 9088 6316
rect 9404 6264 9456 6316
rect 10232 6400 10284 6452
rect 10508 6443 10560 6452
rect 10508 6409 10517 6443
rect 10517 6409 10551 6443
rect 10551 6409 10560 6443
rect 10508 6400 10560 6409
rect 11152 6400 11204 6452
rect 12256 6400 12308 6452
rect 12440 6443 12492 6452
rect 12440 6409 12449 6443
rect 12449 6409 12483 6443
rect 12483 6409 12492 6443
rect 12440 6400 12492 6409
rect 13176 6400 13228 6452
rect 9772 6332 9824 6384
rect 15016 6375 15068 6384
rect 10692 6264 10744 6316
rect 10784 6264 10836 6316
rect 7656 6196 7708 6248
rect 7840 6196 7892 6248
rect 12532 6264 12584 6316
rect 12992 6307 13044 6316
rect 12992 6273 13001 6307
rect 13001 6273 13035 6307
rect 13035 6273 13044 6307
rect 15016 6341 15025 6375
rect 15025 6341 15059 6375
rect 15059 6341 15068 6375
rect 15016 6332 15068 6341
rect 12992 6264 13044 6273
rect 3148 6128 3200 6180
rect 3424 6128 3476 6180
rect 1492 6060 1544 6112
rect 4068 6060 4120 6112
rect 5540 6128 5592 6180
rect 5816 6128 5868 6180
rect 6920 6128 6972 6180
rect 8300 6171 8352 6180
rect 4896 6060 4948 6112
rect 8300 6137 8334 6171
rect 8334 6137 8352 6171
rect 8300 6128 8352 6137
rect 8392 6128 8444 6180
rect 9956 6128 10008 6180
rect 10600 6128 10652 6180
rect 11428 6196 11480 6248
rect 11152 6128 11204 6180
rect 12256 6128 12308 6180
rect 15200 6128 15252 6180
rect 8116 6060 8168 6112
rect 8208 6060 8260 6112
rect 10140 6060 10192 6112
rect 10508 6060 10560 6112
rect 12440 6060 12492 6112
rect 12532 6060 12584 6112
rect 14188 6060 14240 6112
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 2596 5856 2648 5908
rect 2688 5856 2740 5908
rect 4068 5788 4120 5840
rect 1768 5763 1820 5772
rect 1768 5729 1777 5763
rect 1777 5729 1811 5763
rect 1811 5729 1820 5763
rect 1768 5720 1820 5729
rect 2136 5763 2188 5772
rect 2136 5729 2145 5763
rect 2145 5729 2179 5763
rect 2179 5729 2188 5763
rect 2136 5720 2188 5729
rect 4896 5856 4948 5908
rect 5264 5788 5316 5840
rect 5172 5720 5224 5772
rect 3148 5652 3200 5704
rect 3332 5652 3384 5704
rect 5540 5720 5592 5772
rect 6184 5720 6236 5772
rect 6920 5788 6972 5840
rect 7288 5788 7340 5840
rect 8392 5856 8444 5908
rect 8576 5856 8628 5908
rect 7840 5788 7892 5840
rect 8116 5788 8168 5840
rect 8392 5720 8444 5772
rect 8576 5720 8628 5772
rect 8760 5720 8812 5772
rect 9036 5720 9088 5772
rect 9772 5720 9824 5772
rect 9956 5763 10008 5772
rect 9956 5729 9990 5763
rect 9990 5729 10008 5763
rect 9956 5720 10008 5729
rect 10140 5788 10192 5840
rect 11060 5788 11112 5840
rect 13636 5856 13688 5908
rect 14280 5856 14332 5908
rect 11888 5831 11940 5840
rect 11888 5797 11897 5831
rect 11897 5797 11931 5831
rect 11931 5797 11940 5831
rect 11888 5788 11940 5797
rect 12440 5788 12492 5840
rect 13820 5788 13872 5840
rect 15200 5856 15252 5908
rect 6000 5652 6052 5704
rect 7932 5652 7984 5704
rect 8944 5695 8996 5704
rect 8944 5661 8953 5695
rect 8953 5661 8987 5695
rect 8987 5661 8996 5695
rect 8944 5652 8996 5661
rect 9496 5652 9548 5704
rect 3424 5584 3476 5636
rect 4252 5584 4304 5636
rect 5540 5584 5592 5636
rect 3148 5516 3200 5568
rect 3884 5516 3936 5568
rect 5080 5516 5132 5568
rect 5448 5516 5500 5568
rect 5816 5559 5868 5568
rect 5816 5525 5825 5559
rect 5825 5525 5859 5559
rect 5859 5525 5868 5559
rect 5816 5516 5868 5525
rect 7288 5516 7340 5568
rect 7840 5516 7892 5568
rect 8208 5516 8260 5568
rect 9036 5516 9088 5568
rect 12624 5720 12676 5772
rect 13636 5720 13688 5772
rect 14188 5720 14240 5772
rect 11888 5652 11940 5704
rect 12716 5652 12768 5704
rect 13728 5652 13780 5704
rect 14464 5652 14516 5704
rect 14832 5652 14884 5704
rect 12256 5584 12308 5636
rect 14924 5584 14976 5636
rect 10968 5516 11020 5568
rect 11152 5516 11204 5568
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 1952 5176 2004 5228
rect 2780 5312 2832 5364
rect 2872 5244 2924 5296
rect 3332 5312 3384 5364
rect 4068 5312 4120 5364
rect 6736 5312 6788 5364
rect 6920 5312 6972 5364
rect 7196 5312 7248 5364
rect 6276 5244 6328 5296
rect 6644 5244 6696 5296
rect 2136 5040 2188 5092
rect 3976 5040 4028 5092
rect 7012 5176 7064 5228
rect 7196 5176 7248 5228
rect 5908 5108 5960 5160
rect 6000 5108 6052 5160
rect 9588 5312 9640 5364
rect 9680 5312 9732 5364
rect 10876 5312 10928 5364
rect 11888 5312 11940 5364
rect 14464 5312 14516 5364
rect 9956 5219 10008 5228
rect 9220 5108 9272 5160
rect 6184 5040 6236 5092
rect 6736 5040 6788 5092
rect 7012 5040 7064 5092
rect 8208 5040 8260 5092
rect 9956 5185 9965 5219
rect 9965 5185 9999 5219
rect 9999 5185 10008 5219
rect 9956 5176 10008 5185
rect 10324 5176 10376 5228
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 11428 5244 11480 5296
rect 11704 5176 11756 5228
rect 13728 5244 13780 5296
rect 14096 5219 14148 5228
rect 14096 5185 14105 5219
rect 14105 5185 14139 5219
rect 14139 5185 14148 5219
rect 14096 5176 14148 5185
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 4068 4972 4120 5024
rect 4252 4972 4304 5024
rect 4896 4972 4948 5024
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 6920 4972 6972 5024
rect 9496 4972 9548 5024
rect 11796 5040 11848 5092
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 12072 5040 12124 5092
rect 14096 5040 14148 5092
rect 12532 4972 12584 5024
rect 12900 5015 12952 5024
rect 12900 4981 12909 5015
rect 12909 4981 12943 5015
rect 12943 4981 12952 5015
rect 12900 4972 12952 4981
rect 14280 4972 14332 5024
rect 15016 5015 15068 5024
rect 15016 4981 15025 5015
rect 15025 4981 15059 5015
rect 15059 4981 15068 5015
rect 15016 4972 15068 4981
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 1584 4768 1636 4820
rect 3424 4768 3476 4820
rect 4804 4768 4856 4820
rect 5448 4811 5500 4820
rect 5448 4777 5457 4811
rect 5457 4777 5491 4811
rect 5491 4777 5500 4811
rect 5448 4768 5500 4777
rect 5540 4768 5592 4820
rect 6276 4768 6328 4820
rect 3424 4632 3476 4684
rect 5540 4632 5592 4684
rect 3976 4564 4028 4616
rect 6000 4700 6052 4752
rect 6736 4700 6788 4752
rect 6920 4768 6972 4820
rect 11244 4811 11296 4820
rect 11244 4777 11253 4811
rect 11253 4777 11287 4811
rect 11287 4777 11296 4811
rect 11244 4768 11296 4777
rect 12256 4768 12308 4820
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 13084 4768 13136 4820
rect 13728 4811 13780 4820
rect 13728 4777 13737 4811
rect 13737 4777 13771 4811
rect 13771 4777 13780 4811
rect 13728 4768 13780 4777
rect 6552 4632 6604 4684
rect 7196 4632 7248 4684
rect 7288 4632 7340 4684
rect 6920 4564 6972 4616
rect 7472 4564 7524 4616
rect 3792 4496 3844 4548
rect 5172 4496 5224 4548
rect 3884 4428 3936 4480
rect 9680 4632 9732 4684
rect 8760 4564 8812 4616
rect 9772 4564 9824 4616
rect 10416 4700 10468 4752
rect 10968 4700 11020 4752
rect 11796 4700 11848 4752
rect 11888 4700 11940 4752
rect 10324 4632 10376 4684
rect 11152 4632 11204 4684
rect 14004 4632 14056 4684
rect 14556 4632 14608 4684
rect 11244 4564 11296 4616
rect 12532 4607 12584 4616
rect 12532 4573 12541 4607
rect 12541 4573 12575 4607
rect 12575 4573 12584 4607
rect 12532 4564 12584 4573
rect 8944 4496 8996 4548
rect 9956 4496 10008 4548
rect 10876 4496 10928 4548
rect 7932 4428 7984 4480
rect 8116 4428 8168 4480
rect 8760 4428 8812 4480
rect 9680 4471 9732 4480
rect 9680 4437 9689 4471
rect 9689 4437 9723 4471
rect 9723 4437 9732 4471
rect 9680 4428 9732 4437
rect 9772 4428 9824 4480
rect 10692 4428 10744 4480
rect 11888 4428 11940 4480
rect 12348 4496 12400 4548
rect 12716 4496 12768 4548
rect 15016 4496 15068 4548
rect 14004 4428 14056 4480
rect 14648 4471 14700 4480
rect 14648 4437 14657 4471
rect 14657 4437 14691 4471
rect 14691 4437 14700 4471
rect 14648 4428 14700 4437
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 2596 4224 2648 4276
rect 2780 4267 2832 4276
rect 2780 4233 2789 4267
rect 2789 4233 2823 4267
rect 2823 4233 2832 4267
rect 2780 4224 2832 4233
rect 2872 4224 2924 4276
rect 4804 4224 4856 4276
rect 5540 4224 5592 4276
rect 5908 4156 5960 4208
rect 7472 4224 7524 4276
rect 8668 4224 8720 4276
rect 9496 4224 9548 4276
rect 10416 4224 10468 4276
rect 11612 4224 11664 4276
rect 3976 4088 4028 4140
rect 6000 4088 6052 4140
rect 6644 4088 6696 4140
rect 1400 4063 1452 4072
rect 1400 4029 1409 4063
rect 1409 4029 1443 4063
rect 1443 4029 1452 4063
rect 1400 4020 1452 4029
rect 1676 3884 1728 3936
rect 2688 3884 2740 3936
rect 3792 3952 3844 4004
rect 4804 4020 4856 4072
rect 4988 3952 5040 4004
rect 5448 3952 5500 4004
rect 6920 4020 6972 4072
rect 7932 4156 7984 4208
rect 8760 4156 8812 4208
rect 8208 4088 8260 4140
rect 10324 4156 10376 4208
rect 11244 4156 11296 4208
rect 13636 4224 13688 4276
rect 14188 4224 14240 4276
rect 14464 4224 14516 4276
rect 7932 4020 7984 4072
rect 10508 4088 10560 4140
rect 9496 4020 9548 4072
rect 9864 4020 9916 4072
rect 12440 4199 12492 4208
rect 12440 4165 12449 4199
rect 12449 4165 12483 4199
rect 12483 4165 12492 4199
rect 12440 4156 12492 4165
rect 13820 4156 13872 4208
rect 11520 4088 11572 4140
rect 11796 4088 11848 4140
rect 13636 4088 13688 4140
rect 11704 4020 11756 4072
rect 3976 3884 4028 3936
rect 5540 3884 5592 3936
rect 7288 3884 7340 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 9956 3952 10008 4004
rect 10876 3952 10928 4004
rect 10968 3952 11020 4004
rect 14004 4063 14056 4072
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 14648 4020 14700 4072
rect 8760 3884 8812 3893
rect 10232 3884 10284 3936
rect 10508 3884 10560 3936
rect 13268 3952 13320 4004
rect 11336 3884 11388 3936
rect 11612 3884 11664 3936
rect 13636 3927 13688 3936
rect 13636 3893 13645 3927
rect 13645 3893 13679 3927
rect 13679 3893 13688 3927
rect 13636 3884 13688 3893
rect 13820 3884 13872 3936
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 4620 3680 4672 3732
rect 2044 3612 2096 3664
rect 2964 3612 3016 3664
rect 3884 3612 3936 3664
rect 4804 3612 4856 3664
rect 5448 3680 5500 3732
rect 6920 3680 6972 3732
rect 7196 3680 7248 3732
rect 7472 3680 7524 3732
rect 9036 3680 9088 3732
rect 10324 3680 10376 3732
rect 11612 3680 11664 3732
rect 11888 3680 11940 3732
rect 12900 3723 12952 3732
rect 12900 3689 12909 3723
rect 12909 3689 12943 3723
rect 12943 3689 12952 3723
rect 12900 3680 12952 3689
rect 13268 3723 13320 3732
rect 13268 3689 13277 3723
rect 13277 3689 13311 3723
rect 13311 3689 13320 3723
rect 13268 3680 13320 3689
rect 13728 3680 13780 3732
rect 5724 3655 5776 3664
rect 5724 3621 5747 3655
rect 5747 3621 5776 3655
rect 5724 3612 5776 3621
rect 6552 3612 6604 3664
rect 7656 3612 7708 3664
rect 9680 3612 9732 3664
rect 10416 3612 10468 3664
rect 11244 3655 11296 3664
rect 3976 3544 4028 3596
rect 3792 3476 3844 3528
rect 4160 3476 4212 3528
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 4436 3408 4488 3460
rect 7840 3544 7892 3596
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 6920 3476 6972 3528
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 2872 3340 2924 3392
rect 3884 3340 3936 3392
rect 4160 3340 4212 3392
rect 5172 3340 5224 3392
rect 5264 3340 5316 3392
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 8576 3451 8628 3460
rect 8576 3417 8585 3451
rect 8585 3417 8619 3451
rect 8619 3417 8628 3451
rect 8576 3408 8628 3417
rect 8852 3340 8904 3392
rect 9496 3544 9548 3596
rect 9772 3544 9824 3596
rect 9680 3476 9732 3528
rect 10232 3476 10284 3528
rect 9496 3408 9548 3460
rect 9772 3408 9824 3460
rect 11244 3621 11253 3655
rect 11253 3621 11287 3655
rect 11287 3621 11296 3655
rect 11244 3612 11296 3621
rect 12164 3612 12216 3664
rect 12532 3655 12584 3664
rect 12532 3621 12541 3655
rect 12541 3621 12575 3655
rect 12575 3621 12584 3655
rect 12532 3612 12584 3621
rect 13360 3655 13412 3664
rect 13360 3621 13369 3655
rect 13369 3621 13403 3655
rect 13403 3621 13412 3655
rect 13360 3612 13412 3621
rect 13452 3612 13504 3664
rect 11060 3544 11112 3596
rect 14096 3587 14148 3596
rect 11520 3476 11572 3528
rect 12716 3519 12768 3528
rect 12716 3485 12725 3519
rect 12725 3485 12759 3519
rect 12759 3485 12768 3519
rect 12716 3476 12768 3485
rect 12992 3476 13044 3528
rect 13176 3476 13228 3528
rect 13084 3408 13136 3460
rect 13268 3408 13320 3460
rect 14096 3553 14105 3587
rect 14105 3553 14139 3587
rect 14139 3553 14148 3587
rect 14096 3544 14148 3553
rect 14004 3476 14056 3528
rect 14464 3544 14516 3596
rect 14464 3408 14516 3460
rect 10600 3340 10652 3392
rect 11980 3340 12032 3392
rect 12440 3340 12492 3392
rect 15292 3340 15344 3392
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 2044 3136 2096 3188
rect 6736 3136 6788 3188
rect 7472 3136 7524 3188
rect 9128 3136 9180 3188
rect 9588 3136 9640 3188
rect 10232 3136 10284 3188
rect 10968 3136 11020 3188
rect 12532 3136 12584 3188
rect 13084 3136 13136 3188
rect 14096 3136 14148 3188
rect 14372 3136 14424 3188
rect 5356 3068 5408 3120
rect 7840 3068 7892 3120
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 5632 3000 5684 3052
rect 6644 3000 6696 3052
rect 7932 3000 7984 3052
rect 9036 3000 9088 3052
rect 10692 3000 10744 3052
rect 11888 3000 11940 3052
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 14004 3068 14056 3120
rect 14096 3043 14148 3052
rect 5172 2932 5224 2984
rect 6460 2932 6512 2984
rect 6552 2932 6604 2984
rect 8392 2932 8444 2984
rect 8484 2932 8536 2984
rect 9220 2932 9272 2984
rect 9864 2932 9916 2984
rect 1860 2864 1912 2916
rect 2320 2864 2372 2916
rect 4436 2864 4488 2916
rect 4160 2796 4212 2848
rect 4344 2796 4396 2848
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 6368 2864 6420 2916
rect 9312 2864 9364 2916
rect 12624 2932 12676 2984
rect 12716 2932 12768 2984
rect 13360 2932 13412 2984
rect 5816 2796 5868 2805
rect 6276 2796 6328 2848
rect 6644 2796 6696 2848
rect 7012 2796 7064 2848
rect 8576 2796 8628 2848
rect 10140 2864 10192 2916
rect 10324 2907 10376 2916
rect 10324 2873 10333 2907
rect 10333 2873 10367 2907
rect 10367 2873 10376 2907
rect 10324 2864 10376 2873
rect 10600 2864 10652 2916
rect 14096 3009 14105 3043
rect 14105 3009 14139 3043
rect 14139 3009 14148 3043
rect 14096 3000 14148 3009
rect 13544 2932 13596 2984
rect 14832 3000 14884 3052
rect 15292 2932 15344 2984
rect 13912 2864 13964 2916
rect 9864 2839 9916 2848
rect 9864 2805 9873 2839
rect 9873 2805 9907 2839
rect 9907 2805 9916 2839
rect 9864 2796 9916 2805
rect 11428 2839 11480 2848
rect 11428 2805 11437 2839
rect 11437 2805 11471 2839
rect 11471 2805 11480 2839
rect 11428 2796 11480 2805
rect 11612 2796 11664 2848
rect 14464 2796 14516 2848
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 1768 2592 1820 2644
rect 2780 2592 2832 2644
rect 2872 2592 2924 2644
rect 1952 2524 2004 2576
rect 3056 2524 3108 2576
rect 3332 2524 3384 2576
rect 2228 2456 2280 2508
rect 2780 2456 2832 2508
rect 3792 2456 3844 2508
rect 4436 2524 4488 2576
rect 5448 2592 5500 2644
rect 5632 2592 5684 2644
rect 7196 2592 7248 2644
rect 7748 2592 7800 2644
rect 8760 2592 8812 2644
rect 8852 2592 8904 2644
rect 9864 2592 9916 2644
rect 5908 2499 5960 2508
rect 1492 2388 1544 2440
rect 204 2252 256 2304
rect 5908 2465 5917 2499
rect 5917 2465 5951 2499
rect 5951 2465 5960 2499
rect 5908 2456 5960 2465
rect 6460 2456 6512 2508
rect 6736 2456 6788 2508
rect 7564 2456 7616 2508
rect 8668 2524 8720 2576
rect 13636 2592 13688 2644
rect 14096 2592 14148 2644
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 11704 2524 11756 2576
rect 12808 2524 12860 2576
rect 14188 2567 14240 2576
rect 14188 2533 14197 2567
rect 14197 2533 14231 2567
rect 14231 2533 14240 2567
rect 14188 2524 14240 2533
rect 8944 2456 8996 2508
rect 11336 2499 11388 2508
rect 3884 2252 3936 2304
rect 4712 2252 4764 2304
rect 6000 2320 6052 2372
rect 6552 2363 6604 2372
rect 6552 2329 6561 2363
rect 6561 2329 6595 2363
rect 6595 2329 6604 2363
rect 6552 2320 6604 2329
rect 6828 2320 6880 2372
rect 7564 2320 7616 2372
rect 8760 2388 8812 2440
rect 8392 2320 8444 2372
rect 10416 2388 10468 2440
rect 11336 2465 11345 2499
rect 11345 2465 11379 2499
rect 11379 2465 11388 2499
rect 11336 2456 11388 2465
rect 11888 2456 11940 2508
rect 12716 2456 12768 2508
rect 13084 2499 13136 2508
rect 13084 2465 13093 2499
rect 13093 2465 13127 2499
rect 13127 2465 13136 2499
rect 13084 2456 13136 2465
rect 13360 2456 13412 2508
rect 11704 2388 11756 2440
rect 12992 2388 13044 2440
rect 14924 2388 14976 2440
rect 12900 2320 12952 2372
rect 13544 2320 13596 2372
rect 9496 2252 9548 2304
rect 9772 2295 9824 2304
rect 9772 2261 9781 2295
rect 9781 2261 9815 2295
rect 9815 2261 9824 2295
rect 9772 2252 9824 2261
rect 10140 2252 10192 2304
rect 12440 2252 12492 2304
rect 12624 2295 12676 2304
rect 12624 2261 12633 2295
rect 12633 2261 12667 2295
rect 12667 2261 12676 2295
rect 12624 2252 12676 2261
rect 12716 2252 12768 2304
rect 15016 2295 15068 2304
rect 15016 2261 15025 2295
rect 15025 2261 15059 2295
rect 15059 2261 15068 2295
rect 15016 2252 15068 2261
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 3148 2048 3200 2100
rect 15016 2048 15068 2100
rect 2412 1980 2464 2032
rect 12624 1980 12676 2032
rect 1584 1912 1636 1964
rect 11336 1912 11388 1964
rect 12256 1912 12308 1964
rect 14188 1912 14240 1964
rect 3884 1844 3936 1896
rect 6000 1844 6052 1896
rect 9772 1844 9824 1896
rect 10324 1844 10376 1896
rect 12348 1844 12400 1896
rect 5816 1776 5868 1828
rect 6736 1776 6788 1828
rect 7196 1776 7248 1828
rect 8668 1776 8720 1828
rect 11152 1776 11204 1828
rect 15476 1776 15528 1828
rect 4068 1708 4120 1760
rect 15108 1708 15160 1760
rect 4344 1640 4396 1692
rect 8760 1640 8812 1692
rect 3792 1572 3844 1624
rect 5908 1572 5960 1624
rect 9680 1572 9732 1624
rect 4160 1504 4212 1556
rect 4896 1504 4948 1556
rect 11704 1504 11756 1556
rect 2136 1436 2188 1488
rect 6460 1436 6512 1488
rect 11152 1436 11204 1488
rect 8116 1368 8168 1420
rect 9496 1368 9548 1420
rect 6092 1300 6144 1352
rect 8024 1300 8076 1352
rect 9128 824 9180 876
rect 10600 824 10652 876
<< metal2 >>
rect 202 17520 258 18000
rect 570 17520 626 18000
rect 1030 17520 1086 18000
rect 1398 17520 1454 18000
rect 1858 17520 1914 18000
rect 2318 17520 2374 18000
rect 2686 17520 2742 18000
rect 3146 17520 3202 18000
rect 3606 17520 3662 18000
rect 3974 17520 4030 18000
rect 4434 17520 4490 18000
rect 4802 17520 4858 18000
rect 5262 17520 5318 18000
rect 5722 17520 5778 18000
rect 6090 17520 6146 18000
rect 6550 17520 6606 18000
rect 7010 17520 7066 18000
rect 7378 17520 7434 18000
rect 7838 17520 7894 18000
rect 8206 17520 8262 18000
rect 8666 17520 8722 18000
rect 9126 17520 9182 18000
rect 9494 17520 9550 18000
rect 9954 17520 10010 18000
rect 10414 17520 10470 18000
rect 10782 17520 10838 18000
rect 11242 17520 11298 18000
rect 11610 17520 11666 18000
rect 12070 17520 12126 18000
rect 12530 17520 12586 18000
rect 12898 17520 12954 18000
rect 13358 17520 13414 18000
rect 13818 17520 13874 18000
rect 14186 17520 14242 18000
rect 14646 17520 14702 18000
rect 15014 17520 15070 18000
rect 15474 17520 15530 18000
rect 15934 17520 15990 18000
rect 16302 17520 16358 18000
rect 16762 17520 16818 18000
rect 216 16182 244 17520
rect 204 16176 256 16182
rect 204 16118 256 16124
rect 584 15910 612 17520
rect 572 15904 624 15910
rect 572 15846 624 15852
rect 1044 14929 1072 17520
rect 1412 16522 1440 17520
rect 1400 16516 1452 16522
rect 1400 16458 1452 16464
rect 1768 16380 1820 16386
rect 1768 16322 1820 16328
rect 1492 14952 1544 14958
rect 1030 14920 1086 14929
rect 1492 14894 1544 14900
rect 1030 14855 1086 14864
rect 1504 14385 1532 14894
rect 1490 14376 1546 14385
rect 1490 14311 1546 14320
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1596 11354 1624 13466
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1688 11082 1716 13806
rect 1676 11076 1728 11082
rect 1676 11018 1728 11024
rect 1674 9888 1730 9897
rect 1674 9823 1730 9832
rect 1492 9716 1544 9722
rect 1492 9658 1544 9664
rect 1504 7410 1532 9658
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9081 1624 9318
rect 1688 9110 1716 9823
rect 1676 9104 1728 9110
rect 1582 9072 1638 9081
rect 1676 9046 1728 9052
rect 1582 9007 1638 9016
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6934 1624 7142
rect 1584 6928 1636 6934
rect 1398 6896 1454 6905
rect 1584 6870 1636 6876
rect 1398 6831 1400 6840
rect 1452 6831 1454 6840
rect 1400 6802 1452 6808
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 570 3496 626 3505
rect 570 3431 626 3440
rect 204 2304 256 2310
rect 204 2246 256 2252
rect 216 480 244 2246
rect 584 480 612 3431
rect 1412 3058 1440 4014
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1030 2952 1086 2961
rect 1030 2887 1086 2896
rect 1044 480 1072 2887
rect 1412 2428 1440 2994
rect 1504 2666 1532 6054
rect 1688 5522 1716 7346
rect 1780 7342 1808 16322
rect 1872 15094 1900 17520
rect 1950 17368 2006 17377
rect 1950 17303 2006 17312
rect 1860 15088 1912 15094
rect 1860 15030 1912 15036
rect 1858 13424 1914 13433
rect 1858 13359 1914 13368
rect 1872 11898 1900 13359
rect 1964 12594 1992 17303
rect 2228 15564 2280 15570
rect 2228 15506 2280 15512
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 2148 14550 2176 15438
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 2148 13394 2176 14486
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2148 12918 2176 13330
rect 2136 12912 2188 12918
rect 2136 12854 2188 12860
rect 1964 12566 2176 12594
rect 1950 12472 2006 12481
rect 1950 12407 2006 12416
rect 2044 12436 2096 12442
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1872 9897 1900 9998
rect 1858 9888 1914 9897
rect 1858 9823 1914 9832
rect 1964 9738 1992 12407
rect 2044 12378 2096 12384
rect 2056 11898 2084 12378
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 2044 11280 2096 11286
rect 2042 11248 2044 11257
rect 2096 11248 2098 11257
rect 2042 11183 2098 11192
rect 1872 9710 1992 9738
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1780 7002 1808 7142
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1872 6497 1900 9710
rect 1950 9480 2006 9489
rect 1950 9415 1952 9424
rect 2004 9415 2006 9424
rect 1952 9386 2004 9392
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1858 6488 1914 6497
rect 1780 6446 1858 6474
rect 1780 5778 1808 6446
rect 1858 6423 1914 6432
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1688 5494 1808 5522
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1596 4826 1624 4966
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1504 2638 1624 2666
rect 1492 2440 1544 2446
rect 1412 2400 1492 2428
rect 1492 2382 1544 2388
rect 1596 1970 1624 2638
rect 1584 1964 1636 1970
rect 1584 1906 1636 1912
rect 1688 1850 1716 3878
rect 1780 2650 1808 5494
rect 1872 5273 1900 6258
rect 1858 5264 1914 5273
rect 1964 5234 1992 8774
rect 2042 7984 2098 7993
rect 2042 7919 2044 7928
rect 2096 7919 2098 7928
rect 2044 7890 2096 7896
rect 2148 7324 2176 12566
rect 2240 12345 2268 15506
rect 2332 15162 2360 17520
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 2424 14074 2452 16390
rect 2700 15706 2728 17520
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 2792 15450 2820 15982
rect 3056 15972 3108 15978
rect 3056 15914 3108 15920
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 2700 15422 2820 15450
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2410 13832 2466 13841
rect 2410 13767 2466 13776
rect 2320 12912 2372 12918
rect 2320 12854 2372 12860
rect 2226 12336 2282 12345
rect 2226 12271 2282 12280
rect 2332 11830 2360 12854
rect 2424 12782 2452 13767
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2320 11824 2372 11830
rect 2320 11766 2372 11772
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2240 7426 2268 11630
rect 2424 11626 2452 12582
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2412 10532 2464 10538
rect 2412 10474 2464 10480
rect 2424 9926 2452 10474
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2332 9042 2360 9862
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2412 8968 2464 8974
rect 2410 8936 2412 8945
rect 2464 8936 2466 8945
rect 2410 8871 2466 8880
rect 2516 8634 2544 14418
rect 2700 13682 2728 15422
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2608 13654 2728 13682
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2318 8528 2374 8537
rect 2318 8463 2374 8472
rect 2504 8492 2556 8498
rect 2332 8430 2360 8463
rect 2504 8434 2556 8440
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2332 8090 2360 8230
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2516 8022 2544 8434
rect 2504 8016 2556 8022
rect 2504 7958 2556 7964
rect 2502 7848 2558 7857
rect 2502 7783 2558 7792
rect 2240 7398 2360 7426
rect 2516 7410 2544 7783
rect 2056 7296 2176 7324
rect 2228 7336 2280 7342
rect 1858 5199 1914 5208
rect 1952 5228 2004 5234
rect 1872 2922 1900 5199
rect 1952 5170 2004 5176
rect 2056 5114 2084 7296
rect 2228 7278 2280 7284
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2148 6458 2176 6734
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2148 5778 2176 6394
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 1964 5086 2084 5114
rect 2136 5092 2188 5098
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 1964 2582 1992 5086
rect 2136 5034 2188 5040
rect 2148 4808 2176 5034
rect 2056 4780 2176 4808
rect 2056 3890 2084 4780
rect 2056 3862 2176 3890
rect 2042 3768 2098 3777
rect 2042 3703 2098 3712
rect 2056 3670 2084 3703
rect 2044 3664 2096 3670
rect 2044 3606 2096 3612
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 1952 2576 2004 2582
rect 1952 2518 2004 2524
rect 1412 1822 1716 1850
rect 1412 480 1440 1822
rect 2056 1442 2084 3130
rect 2148 1494 2176 3862
rect 2240 2514 2268 7278
rect 2332 7002 2360 7398
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2424 6390 2452 7278
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2320 2916 2372 2922
rect 2320 2858 2372 2864
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 1872 1414 2084 1442
rect 2136 1488 2188 1494
rect 2136 1430 2188 1436
rect 1872 480 1900 1414
rect 2332 480 2360 2858
rect 2424 2038 2452 6190
rect 2516 3754 2544 6598
rect 2608 5914 2636 13654
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2700 11694 2728 12718
rect 2792 12306 2820 15302
rect 2884 13734 2912 15506
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2884 12209 2912 13330
rect 2870 12200 2926 12209
rect 2870 12135 2926 12144
rect 2976 11880 3004 14350
rect 3068 14113 3096 15914
rect 3054 14104 3110 14113
rect 3054 14039 3110 14048
rect 3056 14000 3108 14006
rect 3160 13988 3188 17520
rect 3620 15348 3648 17520
rect 3988 15688 4016 17520
rect 4066 16280 4122 16289
rect 4066 16215 4068 16224
rect 4120 16215 4122 16224
rect 4068 16186 4120 16192
rect 4160 15700 4212 15706
rect 3988 15660 4160 15688
rect 4160 15642 4212 15648
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 4080 15473 4108 15506
rect 4066 15464 4122 15473
rect 4066 15399 4122 15408
rect 3344 15320 3648 15348
rect 3344 14618 3372 15320
rect 3421 15260 3717 15280
rect 3477 15258 3501 15260
rect 3557 15258 3581 15260
rect 3637 15258 3661 15260
rect 3499 15206 3501 15258
rect 3563 15206 3575 15258
rect 3637 15206 3639 15258
rect 3477 15204 3501 15206
rect 3557 15204 3581 15206
rect 3637 15204 3661 15206
rect 3421 15184 3717 15204
rect 4066 15056 4122 15065
rect 4066 14991 4068 15000
rect 4120 14991 4122 15000
rect 4252 15020 4304 15026
rect 4068 14962 4120 14968
rect 4252 14962 4304 14968
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3620 14618 3648 14758
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3884 14544 3936 14550
rect 3988 14521 4016 14758
rect 4264 14657 4292 14962
rect 4250 14648 4306 14657
rect 4250 14583 4306 14592
rect 3884 14486 3936 14492
rect 3974 14512 4030 14521
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3108 13960 3188 13988
rect 3056 13942 3108 13948
rect 3344 13870 3372 14214
rect 3421 14172 3717 14192
rect 3477 14170 3501 14172
rect 3557 14170 3581 14172
rect 3637 14170 3661 14172
rect 3499 14118 3501 14170
rect 3563 14118 3575 14170
rect 3637 14118 3639 14170
rect 3477 14116 3501 14118
rect 3557 14116 3581 14118
rect 3637 14116 3661 14118
rect 3421 14096 3717 14116
rect 3804 14074 3832 14418
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3424 13728 3476 13734
rect 3476 13688 3832 13716
rect 3424 13670 3476 13676
rect 3148 13456 3200 13462
rect 3148 13398 3200 13404
rect 3054 13288 3110 13297
rect 3054 13223 3110 13232
rect 3068 12646 3096 13223
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3160 12442 3188 13398
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3068 12170 3096 12242
rect 3252 12170 3280 12378
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 3240 12164 3292 12170
rect 3240 12106 3292 12112
rect 2884 11852 3004 11880
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2778 11656 2834 11665
rect 2700 11529 2728 11630
rect 2778 11591 2834 11600
rect 2686 11520 2742 11529
rect 2686 11455 2742 11464
rect 2686 11384 2742 11393
rect 2686 11319 2688 11328
rect 2740 11319 2742 11328
rect 2688 11290 2740 11296
rect 2792 11200 2820 11591
rect 2700 11172 2820 11200
rect 2700 10810 2728 11172
rect 2884 11121 2912 11852
rect 3344 11642 3372 13126
rect 3421 13084 3717 13104
rect 3477 13082 3501 13084
rect 3557 13082 3581 13084
rect 3637 13082 3661 13084
rect 3499 13030 3501 13082
rect 3563 13030 3575 13082
rect 3637 13030 3639 13082
rect 3477 13028 3501 13030
rect 3557 13028 3581 13030
rect 3637 13028 3661 13030
rect 3421 13008 3717 13028
rect 3804 12850 3832 13688
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3620 12617 3648 12786
rect 3792 12708 3844 12714
rect 3792 12650 3844 12656
rect 3606 12608 3662 12617
rect 3606 12543 3662 12552
rect 3421 11996 3717 12016
rect 3477 11994 3501 11996
rect 3557 11994 3581 11996
rect 3637 11994 3661 11996
rect 3499 11942 3501 11994
rect 3563 11942 3575 11994
rect 3637 11942 3639 11994
rect 3477 11940 3501 11942
rect 3557 11940 3581 11942
rect 3637 11940 3661 11942
rect 3421 11920 3717 11940
rect 3804 11914 3832 12650
rect 3896 12050 3924 14486
rect 3974 14447 4030 14456
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 3974 14104 4030 14113
rect 3974 14039 4030 14048
rect 3988 12714 4016 14039
rect 4158 13968 4214 13977
rect 4158 13903 4214 13912
rect 4172 13258 4200 13903
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 4158 13016 4214 13025
rect 4158 12951 4214 12960
rect 4172 12866 4200 12951
rect 4080 12838 4200 12866
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 4080 12481 4108 12838
rect 4160 12708 4212 12714
rect 4160 12650 4212 12656
rect 4066 12472 4122 12481
rect 4066 12407 4122 12416
rect 4066 12200 4122 12209
rect 4066 12135 4122 12144
rect 3896 12022 4016 12050
rect 3804 11886 3924 11914
rect 3344 11626 3464 11642
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 3344 11620 3476 11626
rect 3344 11614 3424 11620
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 3068 11150 3096 11290
rect 3056 11144 3108 11150
rect 2870 11112 2926 11121
rect 3056 11086 3108 11092
rect 2870 11047 2926 11056
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 3068 10674 3096 10950
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2700 10266 2728 10610
rect 2884 10577 2912 10610
rect 2870 10568 2926 10577
rect 2870 10503 2926 10512
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 3068 10130 3096 10406
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2792 9625 2820 10066
rect 3160 10062 3188 11562
rect 3344 11150 3372 11614
rect 3424 11562 3476 11568
rect 3792 11552 3844 11558
rect 3422 11520 3478 11529
rect 3792 11494 3844 11500
rect 3422 11455 3478 11464
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3148 10056 3200 10062
rect 3068 10004 3148 10010
rect 3068 9998 3200 10004
rect 3068 9982 3188 9998
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2778 9616 2834 9625
rect 2778 9551 2834 9560
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2700 8634 2728 9386
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2870 8800 2926 8809
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2792 8090 2820 8774
rect 2870 8735 2926 8744
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2700 6866 2728 7822
rect 2792 7449 2820 7890
rect 2778 7440 2834 7449
rect 2778 7375 2834 7384
rect 2780 7268 2832 7274
rect 2780 7210 2832 7216
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2700 5914 2728 6802
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2792 5817 2820 7210
rect 2594 5808 2650 5817
rect 2594 5743 2650 5752
rect 2778 5808 2834 5817
rect 2778 5743 2834 5752
rect 2608 4282 2636 5743
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2792 5148 2820 5306
rect 2884 5302 2912 8735
rect 2976 8430 3004 9862
rect 3068 9722 3096 9982
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 3160 9518 3188 9862
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 3068 8906 3096 9046
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2964 8288 3016 8294
rect 2962 8256 2964 8265
rect 3016 8256 3018 8265
rect 2962 8191 3018 8200
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 7478 3004 7890
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 3068 7324 3096 8842
rect 3160 8634 3188 9318
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 2976 7296 3096 7324
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2792 5120 2912 5148
rect 2686 4856 2742 4865
rect 2686 4791 2742 4800
rect 2596 4276 2648 4282
rect 2596 4218 2648 4224
rect 2700 3942 2728 4791
rect 2884 4282 2912 5120
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2516 3726 2728 3754
rect 2412 2032 2464 2038
rect 2412 1974 2464 1980
rect 2700 480 2728 3726
rect 2792 2825 2820 4218
rect 2870 3904 2926 3913
rect 2870 3839 2926 3848
rect 2884 3398 2912 3839
rect 2976 3670 3004 7296
rect 3160 7274 3188 7822
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2778 2816 2834 2825
rect 2778 2751 2834 2760
rect 2778 2680 2834 2689
rect 2884 2650 2912 3334
rect 2778 2615 2780 2624
rect 2832 2615 2834 2624
rect 2872 2644 2924 2650
rect 2780 2586 2832 2592
rect 2872 2586 2924 2592
rect 3068 2582 3096 6938
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 3160 5710 3188 6122
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3160 4434 3188 5510
rect 3252 4536 3280 11086
rect 3436 10996 3464 11455
rect 3344 10968 3464 10996
rect 3344 10792 3372 10968
rect 3421 10908 3717 10928
rect 3477 10906 3501 10908
rect 3557 10906 3581 10908
rect 3637 10906 3661 10908
rect 3499 10854 3501 10906
rect 3563 10854 3575 10906
rect 3637 10854 3639 10906
rect 3477 10852 3501 10854
rect 3557 10852 3581 10854
rect 3637 10852 3661 10854
rect 3421 10832 3717 10852
rect 3804 10810 3832 11494
rect 3792 10804 3844 10810
rect 3344 10764 3464 10792
rect 3330 10704 3386 10713
rect 3330 10639 3386 10648
rect 3344 8498 3372 10639
rect 3436 10130 3464 10764
rect 3792 10746 3844 10752
rect 3606 10704 3662 10713
rect 3606 10639 3662 10648
rect 3620 10606 3648 10639
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3421 9820 3717 9840
rect 3477 9818 3501 9820
rect 3557 9818 3581 9820
rect 3637 9818 3661 9820
rect 3499 9766 3501 9818
rect 3563 9766 3575 9818
rect 3637 9766 3639 9818
rect 3477 9764 3501 9766
rect 3557 9764 3581 9766
rect 3637 9764 3661 9766
rect 3421 9744 3717 9764
rect 3608 9648 3660 9654
rect 3608 9590 3660 9596
rect 3620 9217 3648 9590
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3606 9208 3662 9217
rect 3606 9143 3662 9152
rect 3712 8820 3740 9522
rect 3804 9382 3832 10746
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3792 8832 3844 8838
rect 3712 8792 3792 8820
rect 3792 8774 3844 8780
rect 3421 8732 3717 8752
rect 3477 8730 3501 8732
rect 3557 8730 3581 8732
rect 3637 8730 3661 8732
rect 3499 8678 3501 8730
rect 3563 8678 3575 8730
rect 3637 8678 3639 8730
rect 3477 8676 3501 8678
rect 3557 8676 3581 8678
rect 3637 8676 3661 8678
rect 3421 8656 3717 8676
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3330 8392 3386 8401
rect 3330 8327 3386 8336
rect 3344 7750 3372 8327
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7954 3464 8230
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3421 7644 3717 7664
rect 3477 7642 3501 7644
rect 3557 7642 3581 7644
rect 3637 7642 3661 7644
rect 3499 7590 3501 7642
rect 3563 7590 3575 7642
rect 3637 7590 3639 7642
rect 3477 7588 3501 7590
rect 3557 7588 3581 7590
rect 3637 7588 3661 7590
rect 3421 7568 3717 7588
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 3804 6458 3832 7890
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3344 5370 3372 5646
rect 3436 5642 3464 6122
rect 3896 5930 3924 11886
rect 3988 8129 4016 12022
rect 4080 11354 4108 12135
rect 4172 12102 4200 12650
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4066 10568 4122 10577
rect 4066 10503 4122 10512
rect 4080 9518 4108 10503
rect 4059 9512 4111 9518
rect 4059 9454 4111 9460
rect 4172 8906 4200 11154
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3974 8120 4030 8129
rect 3974 8055 4030 8064
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3804 5902 3924 5930
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3436 4690 3464 4762
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3804 4554 3832 5902
rect 3882 5672 3938 5681
rect 3882 5607 3938 5616
rect 3896 5574 3924 5607
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3988 5098 4016 7686
rect 4080 7585 4108 8774
rect 4066 7576 4122 7585
rect 4066 7511 4122 7520
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 4080 6458 4108 7142
rect 4158 6896 4214 6905
rect 4158 6831 4214 6840
rect 4172 6633 4200 6831
rect 4158 6624 4214 6633
rect 4158 6559 4214 6568
rect 4158 6488 4214 6497
rect 4068 6452 4120 6458
rect 4158 6423 4214 6432
rect 4068 6394 4120 6400
rect 4172 6254 4200 6423
rect 4160 6248 4212 6254
rect 4066 6216 4122 6225
rect 4160 6190 4212 6196
rect 4066 6151 4122 6160
rect 4080 6118 4108 6151
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4158 6080 4214 6089
rect 4264 6066 4292 14418
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4356 13308 4384 14350
rect 4448 13977 4476 17520
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 4434 13968 4490 13977
rect 4434 13903 4490 13912
rect 4540 13802 4568 15302
rect 4618 13968 4674 13977
rect 4618 13903 4620 13912
rect 4672 13903 4674 13912
rect 4620 13874 4672 13880
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4526 13696 4582 13705
rect 4526 13631 4582 13640
rect 4436 13320 4488 13326
rect 4356 13280 4436 13308
rect 4436 13262 4488 13268
rect 4448 12850 4476 13262
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 4342 12744 4398 12753
rect 4342 12679 4398 12688
rect 4356 12646 4384 12679
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4448 12306 4476 12582
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4344 12164 4396 12170
rect 4344 12106 4396 12112
rect 4356 11354 4384 12106
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4540 10690 4568 13631
rect 4618 13560 4674 13569
rect 4618 13495 4674 13504
rect 4632 13462 4660 13495
rect 4620 13456 4672 13462
rect 4620 13398 4672 13404
rect 4724 13025 4752 15506
rect 4816 14958 4844 17520
rect 4988 16312 5040 16318
rect 4988 16254 5040 16260
rect 5000 15638 5028 16254
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4896 15020 4948 15026
rect 4896 14962 4948 14968
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4710 13016 4766 13025
rect 4710 12951 4766 12960
rect 4816 12918 4844 13874
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 4620 12844 4672 12850
rect 4672 12804 4752 12832
rect 4620 12786 4672 12792
rect 4724 12458 4752 12804
rect 4724 12430 4844 12458
rect 4712 12300 4764 12306
rect 4816 12288 4844 12430
rect 4764 12260 4844 12288
rect 4712 12242 4764 12248
rect 4712 12164 4764 12170
rect 4908 12152 4936 14962
rect 4712 12106 4764 12112
rect 4816 12124 4936 12152
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4448 10662 4568 10690
rect 4342 10160 4398 10169
rect 4342 10095 4398 10104
rect 4356 8362 4384 10095
rect 4448 10062 4476 10662
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4448 8634 4476 8910
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4540 8498 4568 10134
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4632 8294 4660 12038
rect 4724 10538 4752 12106
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 4816 10418 4844 12124
rect 4894 12064 4950 12073
rect 4894 11999 4950 12008
rect 4908 11694 4936 11999
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4908 11014 4936 11630
rect 5000 11150 5028 15438
rect 5276 15162 5304 17520
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 5264 15156 5316 15162
rect 5552 15144 5580 15370
rect 5264 15098 5316 15104
rect 5368 15116 5580 15144
rect 5630 15192 5686 15201
rect 5630 15127 5686 15136
rect 5184 15042 5212 15098
rect 5368 15042 5396 15116
rect 5184 15014 5396 15042
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5460 14793 5488 14962
rect 5644 14890 5672 15127
rect 5736 15094 5764 17520
rect 6104 16046 6132 17520
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6092 16040 6144 16046
rect 6092 15982 6144 15988
rect 5886 15804 6182 15824
rect 5942 15802 5966 15804
rect 6022 15802 6046 15804
rect 6102 15802 6126 15804
rect 5964 15750 5966 15802
rect 6028 15750 6040 15802
rect 6102 15750 6104 15802
rect 5942 15748 5966 15750
rect 6022 15748 6046 15750
rect 6102 15748 6126 15750
rect 5886 15728 6182 15748
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5632 14884 5684 14890
rect 5632 14826 5684 14832
rect 5724 14816 5776 14822
rect 5446 14784 5502 14793
rect 5776 14793 6316 14804
rect 5776 14784 6330 14793
rect 5776 14776 6274 14784
rect 5724 14758 5776 14764
rect 5446 14719 5502 14728
rect 5886 14716 6182 14736
rect 6274 14719 6330 14728
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6126 14716
rect 5964 14662 5966 14714
rect 6028 14662 6040 14714
rect 6102 14662 6104 14714
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6126 14662
rect 5886 14640 6182 14660
rect 6380 14618 6408 16050
rect 6564 15706 6592 17520
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 5184 14006 5212 14554
rect 6460 14544 6512 14550
rect 6460 14486 6512 14492
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5276 13297 5304 13398
rect 5262 13288 5318 13297
rect 5184 13246 5262 13274
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5092 11529 5120 12786
rect 5078 11520 5134 11529
rect 5078 11455 5134 11464
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4896 11008 4948 11014
rect 5000 10985 5028 11086
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 4896 10950 4948 10956
rect 4986 10976 5042 10985
rect 4908 10674 4936 10950
rect 4986 10911 5042 10920
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4816 10390 5028 10418
rect 4802 10296 4858 10305
rect 4802 10231 4858 10240
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4356 7478 4384 7822
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4356 7177 4384 7414
rect 4540 7313 4568 7822
rect 4526 7304 4582 7313
rect 4526 7239 4582 7248
rect 4724 7206 4752 8434
rect 4712 7200 4764 7206
rect 4342 7168 4398 7177
rect 4712 7142 4764 7148
rect 4342 7103 4398 7112
rect 4434 7032 4490 7041
rect 4434 6967 4436 6976
rect 4488 6967 4490 6976
rect 4436 6938 4488 6944
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 4436 6792 4488 6798
rect 4434 6760 4436 6769
rect 4488 6760 4490 6769
rect 4434 6695 4490 6704
rect 4264 6038 4384 6066
rect 4158 6015 4214 6024
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4080 5545 4108 5782
rect 4066 5536 4122 5545
rect 4066 5471 4122 5480
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4080 5137 4108 5306
rect 4066 5128 4122 5137
rect 3976 5092 4028 5098
rect 4066 5063 4122 5072
rect 3976 5034 4028 5040
rect 3988 4622 4016 5034
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3976 4616 4028 4622
rect 3882 4584 3938 4593
rect 3792 4548 3844 4554
rect 3252 4508 3372 4536
rect 3160 4406 3280 4434
rect 3056 2576 3108 2582
rect 3056 2518 3108 2524
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 513 2820 2450
rect 3148 2100 3200 2106
rect 3148 2042 3200 2048
rect 2778 504 2834 513
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1398 0 1454 480
rect 1858 0 1914 480
rect 2318 0 2374 480
rect 2686 0 2742 480
rect 3160 480 3188 2042
rect 3252 1442 3280 4406
rect 3344 2582 3372 4508
rect 3976 4558 4028 4564
rect 3882 4519 3938 4528
rect 3792 4490 3844 4496
rect 3896 4486 3924 4519
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3882 4312 3938 4321
rect 3882 4247 3938 4256
rect 3790 4040 3846 4049
rect 3790 3975 3792 3984
rect 3844 3975 3846 3984
rect 3792 3946 3844 3952
rect 3896 3670 3924 4247
rect 3988 4146 4016 4558
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3988 3942 4016 4082
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3988 3602 4016 3878
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3792 3528 3844 3534
rect 4080 3482 4108 4966
rect 4172 3534 4200 6015
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4264 5030 4292 5578
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 3792 3470 3844 3476
rect 3421 3292 3717 3312
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3804 3210 3832 3470
rect 3896 3454 4108 3482
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 3896 3398 3924 3454
rect 3884 3392 3936 3398
rect 4160 3392 4212 3398
rect 3884 3334 3936 3340
rect 3988 3352 4160 3380
rect 3804 3182 3924 3210
rect 3332 2576 3384 2582
rect 3332 2518 3384 2524
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3421 2128 3717 2148
rect 3804 1630 3832 2450
rect 3896 2310 3924 3182
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3896 1902 3924 2246
rect 3884 1896 3936 1902
rect 3884 1838 3936 1844
rect 3792 1624 3844 1630
rect 3792 1566 3844 1572
rect 3252 1414 3648 1442
rect 3620 480 3648 1414
rect 3988 480 4016 3352
rect 4160 3334 4212 3340
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4066 2544 4122 2553
rect 4066 2479 4122 2488
rect 4080 1766 4108 2479
rect 4068 1760 4120 1766
rect 4068 1702 4120 1708
rect 4172 1562 4200 2790
rect 4264 1873 4292 4966
rect 4356 2854 4384 6038
rect 4448 3466 4476 6695
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 4865 4568 6598
rect 4632 5409 4660 6870
rect 4710 6352 4766 6361
rect 4710 6287 4766 6296
rect 4724 5681 4752 6287
rect 4710 5672 4766 5681
rect 4710 5607 4766 5616
rect 4618 5400 4674 5409
rect 4618 5335 4674 5344
rect 4526 4856 4582 4865
rect 4816 4826 4844 10231
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4908 8906 4936 9114
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4908 8294 4936 8366
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4908 7410 4936 8230
rect 5000 7721 5028 10390
rect 5092 9518 5120 11018
rect 5184 10062 5212 13246
rect 5262 13223 5318 13232
rect 5368 12986 5396 14350
rect 6092 14340 6144 14346
rect 6092 14282 6144 14288
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 5906 14240 5962 14249
rect 5906 14175 5962 14184
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5446 13560 5502 13569
rect 5552 13530 5580 13874
rect 5446 13495 5502 13504
rect 5540 13524 5592 13530
rect 5460 12986 5488 13495
rect 5540 13466 5592 13472
rect 5644 13462 5672 14010
rect 5920 13938 5948 14175
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 6104 13716 6132 14282
rect 6196 13870 6224 14282
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6380 13977 6408 14010
rect 6366 13968 6422 13977
rect 6366 13903 6422 13912
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 5722 13696 5778 13705
rect 6104 13688 6316 13716
rect 5722 13631 5778 13640
rect 5736 13530 5764 13631
rect 5886 13628 6182 13648
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6126 13628
rect 5964 13574 5966 13626
rect 6028 13574 6040 13626
rect 6102 13574 6104 13626
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6126 13574
rect 5886 13552 6182 13572
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5632 13456 5684 13462
rect 5632 13398 5684 13404
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5736 12940 5948 12968
rect 5264 12912 5316 12918
rect 5264 12854 5316 12860
rect 5354 12880 5410 12889
rect 5276 12306 5304 12854
rect 5354 12815 5410 12824
rect 5538 12880 5594 12889
rect 5538 12815 5594 12824
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5276 11626 5304 12242
rect 5368 12209 5396 12815
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5354 12200 5410 12209
rect 5354 12135 5410 12144
rect 5460 12102 5488 12650
rect 5552 12481 5580 12815
rect 5736 12696 5764 12940
rect 5920 12850 5948 12940
rect 6104 12889 6132 13126
rect 6090 12880 6146 12889
rect 5908 12844 5960 12850
rect 6090 12815 6092 12824
rect 5908 12786 5960 12792
rect 6144 12815 6146 12824
rect 6092 12786 6144 12792
rect 5644 12668 5764 12696
rect 5538 12472 5594 12481
rect 5538 12407 5594 12416
rect 5448 12096 5500 12102
rect 5354 12064 5410 12073
rect 5448 12038 5500 12044
rect 5354 11999 5410 12008
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5368 11150 5396 11999
rect 5448 11212 5500 11218
rect 5500 11172 5580 11200
rect 5448 11154 5500 11160
rect 5356 11144 5408 11150
rect 5552 11121 5580 11172
rect 5356 11086 5408 11092
rect 5538 11112 5594 11121
rect 5368 10520 5396 11086
rect 5538 11047 5594 11056
rect 5368 10492 5488 10520
rect 5460 10062 5488 10492
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5184 9761 5212 9998
rect 5170 9752 5226 9761
rect 5460 9722 5488 9998
rect 5552 9722 5580 10066
rect 5644 9994 5672 12668
rect 5816 12640 5868 12646
rect 5722 12608 5778 12617
rect 5816 12582 5868 12588
rect 5722 12543 5778 12552
rect 5736 12170 5764 12543
rect 5819 12356 5847 12582
rect 5886 12540 6182 12560
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6126 12540
rect 5964 12486 5966 12538
rect 6028 12486 6040 12538
rect 6102 12486 6104 12538
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6126 12486
rect 5886 12464 6182 12484
rect 5819 12328 5856 12356
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5828 11778 5856 12328
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 6012 11898 6040 12174
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6104 11898 6132 12038
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6196 11830 6224 12106
rect 6184 11824 6236 11830
rect 5828 11762 5948 11778
rect 6184 11766 6236 11772
rect 5828 11756 5960 11762
rect 5828 11750 5908 11756
rect 5908 11698 5960 11704
rect 6288 11694 6316 13688
rect 6472 13274 6500 14486
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6380 13246 6500 13274
rect 6380 12481 6408 13246
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6366 12472 6422 12481
rect 6366 12407 6422 12416
rect 6472 12084 6500 13126
rect 6564 12889 6592 14214
rect 6656 13977 6684 16458
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6748 14657 6776 15438
rect 6826 15328 6882 15337
rect 6826 15263 6882 15272
rect 6734 14648 6790 14657
rect 6734 14583 6790 14592
rect 6748 14414 6776 14583
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6840 14006 6868 15263
rect 6932 14074 6960 15982
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6828 14000 6880 14006
rect 6642 13968 6698 13977
rect 6828 13942 6880 13948
rect 6642 13903 6698 13912
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6550 12880 6606 12889
rect 6550 12815 6606 12824
rect 6656 12696 6684 13806
rect 7024 13705 7052 17520
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7102 15192 7158 15201
rect 7102 15127 7158 15136
rect 7116 14550 7144 15127
rect 7208 14657 7236 15506
rect 7392 15162 7420 17520
rect 7470 16008 7526 16017
rect 7470 15943 7526 15952
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7194 14648 7250 14657
rect 7194 14583 7250 14592
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7010 13696 7066 13705
rect 7010 13631 7066 13640
rect 7208 13394 7236 13874
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7024 12986 7052 13330
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6564 12668 6684 12696
rect 6564 12152 6592 12668
rect 6748 12617 6776 12854
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 6734 12608 6790 12617
rect 6734 12543 6790 12552
rect 6644 12368 6696 12374
rect 6920 12368 6972 12374
rect 6696 12328 6920 12356
rect 6644 12310 6696 12316
rect 6920 12310 6972 12316
rect 6564 12124 6684 12152
rect 6380 12056 6500 12084
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 5722 11520 5778 11529
rect 5778 11478 5856 11506
rect 5722 11455 5778 11464
rect 5722 11384 5778 11393
rect 5722 11319 5778 11328
rect 5736 11014 5764 11319
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5828 10792 5856 11478
rect 5886 11452 6182 11472
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6126 11452
rect 5964 11398 5966 11450
rect 6028 11398 6040 11450
rect 6102 11398 6104 11450
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6126 11398
rect 5886 11376 6182 11396
rect 5908 10804 5960 10810
rect 5828 10764 5908 10792
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5736 10198 5764 10542
rect 5828 10198 5856 10764
rect 5908 10746 5960 10752
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 5886 10364 6182 10384
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6126 10364
rect 5964 10310 5966 10362
rect 6028 10310 6040 10362
rect 6102 10310 6104 10362
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6126 10310
rect 5886 10288 6182 10308
rect 6288 10198 6316 10406
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 6092 9920 6144 9926
rect 6144 9880 6316 9908
rect 6092 9862 6144 9868
rect 5170 9687 5226 9696
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5078 9208 5134 9217
rect 5078 9143 5080 9152
rect 5132 9143 5134 9152
rect 5080 9114 5132 9120
rect 5460 8106 5488 9658
rect 5552 9450 5580 9658
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5886 9276 6182 9296
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6126 9276
rect 5964 9222 5966 9274
rect 6028 9222 6040 9274
rect 6102 9222 6104 9274
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6126 9222
rect 5886 9200 6182 9220
rect 6288 9042 6316 9880
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5552 8265 5580 8366
rect 5644 8362 5672 8978
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5538 8256 5594 8265
rect 5538 8191 5594 8200
rect 5460 8078 5672 8106
rect 5644 7954 5672 8078
rect 5828 8004 5856 8978
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6196 8809 6224 8842
rect 6182 8800 6238 8809
rect 6182 8735 6238 8744
rect 6288 8634 6316 8978
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 5886 8188 6182 8208
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6126 8188
rect 5964 8134 5966 8186
rect 6028 8134 6040 8186
rect 6102 8134 6104 8186
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6126 8134
rect 5886 8112 6182 8132
rect 6274 8120 6330 8129
rect 6274 8055 6330 8064
rect 5828 7976 6132 8004
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 4986 7712 5042 7721
rect 4986 7647 5042 7656
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 6322 4936 6734
rect 4986 6352 5042 6361
rect 4896 6316 4948 6322
rect 4986 6287 5042 6296
rect 4896 6258 4948 6264
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4908 5914 4936 6054
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4526 4791 4582 4800
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4816 4434 4844 4762
rect 4724 4406 4844 4434
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4526 3632 4582 3641
rect 4526 3567 4582 3576
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4434 3360 4490 3369
rect 4434 3295 4490 3304
rect 4448 2922 4476 3295
rect 4540 2961 4568 3567
rect 4632 3534 4660 3674
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4526 2952 4582 2961
rect 4436 2916 4488 2922
rect 4526 2887 4582 2896
rect 4436 2858 4488 2864
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4434 2816 4490 2825
rect 4250 1864 4306 1873
rect 4250 1799 4306 1808
rect 4356 1698 4384 2790
rect 4434 2751 4490 2760
rect 4448 2582 4476 2751
rect 4436 2576 4488 2582
rect 4436 2518 4488 2524
rect 4724 2310 4752 4406
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4816 4078 4844 4218
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4816 3233 4844 3606
rect 4802 3224 4858 3233
rect 4802 3159 4858 3168
rect 4802 2952 4858 2961
rect 4802 2887 4858 2896
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 4434 2000 4490 2009
rect 4434 1935 4490 1944
rect 4344 1692 4396 1698
rect 4344 1634 4396 1640
rect 4160 1556 4212 1562
rect 4160 1498 4212 1504
rect 4448 480 4476 1935
rect 4816 480 4844 2887
rect 4908 1562 4936 4966
rect 5000 4729 5028 6287
rect 5092 5658 5120 7890
rect 5264 7880 5316 7886
rect 5316 7840 5396 7868
rect 5264 7822 5316 7828
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 5184 7002 5212 7210
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5184 5778 5212 6734
rect 5276 6497 5304 7686
rect 5368 7206 5396 7840
rect 5446 7848 5502 7857
rect 5446 7783 5448 7792
rect 5500 7783 5502 7792
rect 5448 7754 5500 7760
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5908 7472 5960 7478
rect 5736 7432 5908 7460
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5356 7200 5408 7206
rect 5460 7177 5488 7210
rect 5356 7142 5408 7148
rect 5446 7168 5502 7177
rect 5446 7103 5502 7112
rect 5736 7041 5764 7432
rect 5908 7414 5960 7420
rect 6012 7342 6040 7482
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6104 7188 6132 7976
rect 6288 7698 6316 8055
rect 6196 7670 6316 7698
rect 6196 7478 6224 7670
rect 6274 7576 6330 7585
rect 6274 7511 6276 7520
rect 6328 7511 6330 7520
rect 6276 7482 6328 7488
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 5828 7160 6132 7188
rect 6276 7200 6328 7206
rect 5722 7032 5778 7041
rect 5722 6967 5778 6976
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5262 6488 5318 6497
rect 5262 6423 5318 6432
rect 5276 5846 5304 6423
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5092 5630 5304 5658
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4986 4720 5042 4729
rect 4986 4655 5042 4664
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 5000 2417 5028 3946
rect 5092 3534 5120 5510
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5184 3398 5212 4490
rect 5276 3398 5304 5630
rect 5368 5137 5396 6870
rect 5828 6644 5856 7160
rect 6276 7142 6328 7148
rect 5886 7100 6182 7120
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6126 7100
rect 5964 7046 5966 7098
rect 6028 7046 6040 7098
rect 6102 7046 6104 7098
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6126 7046
rect 5886 7024 6182 7044
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 5828 6616 5948 6644
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5460 6089 5488 6190
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5446 6080 5502 6089
rect 5446 6015 5502 6024
rect 5552 5778 5580 6122
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5354 5128 5410 5137
rect 5354 5063 5410 5072
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5262 3224 5318 3233
rect 5262 3159 5318 3168
rect 5170 3088 5226 3097
rect 5170 3023 5226 3032
rect 5184 2990 5212 3023
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5276 2666 5304 3159
rect 5368 3126 5396 5063
rect 5460 4826 5488 5510
rect 5552 4826 5580 5578
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5552 4282 5580 4626
rect 5644 4536 5672 6190
rect 5816 6180 5868 6186
rect 5816 6122 5868 6128
rect 5828 5896 5856 6122
rect 5920 6100 5948 6616
rect 6104 6254 6132 6802
rect 6288 6798 6316 7142
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 5920 6072 6316 6100
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 5828 5868 5948 5896
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5828 5273 5856 5510
rect 5814 5264 5870 5273
rect 5814 5199 5870 5208
rect 5722 4856 5778 4865
rect 5722 4791 5778 4800
rect 5736 4604 5764 4791
rect 5828 4729 5856 5199
rect 5920 5166 5948 5868
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6012 5166 6040 5646
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 6196 5098 6224 5714
rect 6288 5302 6316 6072
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 6288 4826 6316 4966
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6000 4752 6052 4758
rect 5814 4720 5870 4729
rect 6000 4694 6052 4700
rect 5814 4655 5870 4664
rect 5736 4576 5948 4604
rect 5644 4508 5764 4536
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5460 3738 5488 3946
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5552 3233 5580 3878
rect 5630 3768 5686 3777
rect 5630 3703 5686 3712
rect 5538 3224 5594 3233
rect 5538 3159 5594 3168
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 5644 3058 5672 3703
rect 5736 3670 5764 4508
rect 5814 4448 5870 4457
rect 5814 4383 5870 4392
rect 5724 3664 5776 3670
rect 5724 3606 5776 3612
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5828 2938 5856 4383
rect 5920 4214 5948 4576
rect 5908 4208 5960 4214
rect 5908 4150 5960 4156
rect 6012 4146 6040 4694
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5886 3836 6182 3856
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 5736 2910 5856 2938
rect 5630 2680 5686 2689
rect 5276 2650 5488 2666
rect 5276 2644 5500 2650
rect 5276 2638 5448 2644
rect 5630 2615 5632 2624
rect 5448 2586 5500 2592
rect 5684 2615 5686 2624
rect 5632 2586 5684 2592
rect 5262 2544 5318 2553
rect 5262 2479 5318 2488
rect 4986 2408 5042 2417
rect 4986 2343 5042 2352
rect 4896 1556 4948 1562
rect 4896 1498 4948 1504
rect 5276 480 5304 2479
rect 5736 480 5764 2910
rect 6288 2854 6316 4762
rect 6380 2922 6408 12056
rect 6656 11880 6684 12124
rect 6564 11852 6684 11880
rect 6458 11520 6514 11529
rect 6458 11455 6514 11464
rect 6472 11200 6500 11455
rect 6564 11354 6592 11852
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6552 11212 6604 11218
rect 6472 11172 6552 11200
rect 6552 11154 6604 11160
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6472 10606 6500 10746
rect 6460 10600 6512 10606
rect 6564 10577 6592 11018
rect 6460 10542 6512 10548
rect 6550 10568 6606 10577
rect 6550 10503 6606 10512
rect 6458 10432 6514 10441
rect 6458 10367 6514 10376
rect 6472 2990 6500 10367
rect 6564 9654 6592 10503
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6564 6322 6592 8026
rect 6656 6746 6684 11698
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6748 11354 6776 11562
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6840 11014 6868 11766
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6932 11218 6960 11562
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6748 9926 6776 10950
rect 6826 10840 6882 10849
rect 6826 10775 6882 10784
rect 6840 10577 6868 10775
rect 6932 10606 6960 11154
rect 6920 10600 6972 10606
rect 6826 10568 6882 10577
rect 6920 10542 6972 10548
rect 6826 10503 6882 10512
rect 6932 10062 6960 10542
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6932 9518 6960 9998
rect 7024 9738 7052 12650
rect 7102 11520 7158 11529
rect 7102 11455 7158 11464
rect 7116 11082 7144 11455
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7102 10976 7158 10985
rect 7102 10911 7158 10920
rect 7116 10606 7144 10911
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7208 10266 7236 13126
rect 7300 12782 7328 14894
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7392 13326 7420 14758
rect 7484 14618 7512 15943
rect 7656 15564 7708 15570
rect 7576 15524 7656 15552
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7576 14074 7604 15524
rect 7656 15506 7708 15512
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7654 14784 7710 14793
rect 7654 14719 7710 14728
rect 7668 14618 7696 14719
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7760 14498 7788 14962
rect 7852 14600 7880 17520
rect 8220 16454 8248 17520
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8680 16368 8708 17520
rect 8680 16340 9076 16368
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8300 15632 8352 15638
rect 8668 15632 8720 15638
rect 8300 15574 8352 15580
rect 8404 15592 8668 15620
rect 8312 15348 8340 15574
rect 8404 15502 8432 15592
rect 8668 15574 8720 15580
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8206 15328 8262 15337
rect 8312 15320 8708 15348
rect 8206 15263 8262 15272
rect 7932 14612 7984 14618
rect 7852 14572 7932 14600
rect 7932 14554 7984 14560
rect 8116 14544 8168 14550
rect 7760 14492 8116 14498
rect 7760 14486 8168 14492
rect 7760 14470 8156 14486
rect 8220 14482 8248 15263
rect 8352 15260 8648 15280
rect 8408 15258 8432 15260
rect 8488 15258 8512 15260
rect 8568 15258 8592 15260
rect 8430 15206 8432 15258
rect 8494 15206 8506 15258
rect 8568 15206 8570 15258
rect 8408 15204 8432 15206
rect 8488 15204 8512 15206
rect 8568 15204 8592 15206
rect 8352 15184 8648 15204
rect 8680 15162 8708 15320
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8666 14512 8722 14521
rect 8208 14476 8260 14482
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7484 13172 7512 13942
rect 7564 13864 7616 13870
rect 7668 13852 7696 14010
rect 7760 13938 7788 14470
rect 8666 14447 8722 14456
rect 8208 14418 8260 14424
rect 8300 14408 8352 14414
rect 7838 14376 7894 14385
rect 7838 14311 7894 14320
rect 7944 14356 8300 14362
rect 7944 14350 8352 14356
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 7944 14334 8340 14350
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7852 13870 7880 14311
rect 7616 13824 7696 13852
rect 7840 13864 7892 13870
rect 7564 13806 7616 13812
rect 7840 13806 7892 13812
rect 7564 13728 7616 13734
rect 7748 13728 7800 13734
rect 7564 13670 7616 13676
rect 7746 13696 7748 13705
rect 7800 13696 7802 13705
rect 7392 13144 7512 13172
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7392 12628 7420 13144
rect 7576 12714 7604 13670
rect 7746 13631 7802 13640
rect 7760 13394 7788 13631
rect 7748 13388 7800 13394
rect 7668 13348 7748 13376
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7300 12600 7420 12628
rect 7300 12102 7328 12600
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7378 12336 7434 12345
rect 7378 12271 7434 12280
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7392 11540 7420 12271
rect 7484 11694 7512 12378
rect 7576 12345 7604 12378
rect 7562 12336 7618 12345
rect 7562 12271 7618 12280
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7392 11512 7512 11540
rect 7576 11529 7604 12174
rect 7378 10432 7434 10441
rect 7378 10367 7434 10376
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7024 9710 7236 9738
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6748 8537 6776 9318
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 6932 8838 6960 9046
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6734 8528 6790 8537
rect 6734 8463 6790 8472
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6748 8090 6776 8298
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 7392 6776 7822
rect 6840 7546 6868 8774
rect 6918 8528 6974 8537
rect 6918 8463 6974 8472
rect 6932 8430 6960 8463
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 7024 8022 7052 9046
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7116 8634 7144 8978
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7102 8256 7158 8265
rect 7102 8191 7158 8200
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6828 7404 6880 7410
rect 6748 7364 6828 7392
rect 6828 7346 6880 7352
rect 6840 6934 6868 7346
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6656 6718 6868 6746
rect 6736 6656 6788 6662
rect 6656 6616 6736 6644
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6656 5386 6684 6616
rect 6736 6598 6788 6604
rect 6734 6352 6790 6361
rect 6734 6287 6790 6296
rect 6564 5358 6684 5386
rect 6748 5370 6776 6287
rect 6736 5364 6788 5370
rect 6564 4690 6592 5358
rect 6736 5306 6788 5312
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6656 5001 6684 5238
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6642 4992 6698 5001
rect 6642 4927 6698 4936
rect 6748 4842 6776 5034
rect 6656 4814 6776 4842
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6656 4570 6684 4814
rect 6736 4752 6788 4758
rect 6736 4694 6788 4700
rect 6564 4542 6684 4570
rect 6564 4049 6592 4542
rect 6748 4185 6776 4694
rect 6734 4176 6790 4185
rect 6644 4140 6696 4146
rect 6734 4111 6790 4120
rect 6644 4082 6696 4088
rect 6550 4040 6606 4049
rect 6550 3975 6606 3984
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6564 2990 6592 3606
rect 6656 3058 6684 4082
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6368 2916 6420 2922
rect 6368 2858 6420 2864
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 6276 2848 6328 2854
rect 6276 2790 6328 2796
rect 6644 2848 6696 2854
rect 6748 2825 6776 3130
rect 6644 2790 6696 2796
rect 6734 2816 6790 2825
rect 5828 1834 5856 2790
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 6550 2680 6606 2689
rect 6550 2615 6606 2624
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 5816 1828 5868 1834
rect 5816 1770 5868 1776
rect 5920 1630 5948 2450
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 6012 1902 6040 2314
rect 6000 1896 6052 1902
rect 6000 1838 6052 1844
rect 5908 1624 5960 1630
rect 6012 1601 6040 1838
rect 5908 1566 5960 1572
rect 5998 1592 6054 1601
rect 5998 1527 6054 1536
rect 6472 1494 6500 2450
rect 6564 2378 6592 2615
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 6460 1488 6512 1494
rect 6656 1442 6684 2790
rect 6734 2751 6790 2760
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6748 1834 6776 2450
rect 6840 2378 6868 6718
rect 6932 6186 6960 7686
rect 7116 7392 7144 8191
rect 7024 7364 7144 7392
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6932 5370 6960 5782
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 7024 5234 7052 7364
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7010 5128 7066 5137
rect 7010 5063 7012 5072
rect 7064 5063 7066 5072
rect 7012 5034 7064 5040
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 4826 6960 4966
rect 7010 4856 7066 4865
rect 6920 4820 6972 4826
rect 7010 4791 7066 4800
rect 6920 4762 6972 4768
rect 6920 4616 6972 4622
rect 7024 4593 7052 4791
rect 6920 4558 6972 4564
rect 7010 4584 7066 4593
rect 6932 4078 6960 4558
rect 7010 4519 7066 4528
rect 7116 4298 7144 7210
rect 7208 6497 7236 9710
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7300 7206 7328 7958
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7392 6610 7420 10367
rect 7484 8673 7512 11512
rect 7562 11520 7618 11529
rect 7668 11506 7696 13348
rect 7748 13330 7800 13336
rect 7944 13326 7972 14334
rect 8496 14260 8524 14350
rect 8036 14232 8524 14260
rect 8036 14006 8064 14232
rect 8352 14172 8648 14192
rect 8408 14170 8432 14172
rect 8488 14170 8512 14172
rect 8568 14170 8592 14172
rect 8430 14118 8432 14170
rect 8494 14118 8506 14170
rect 8568 14118 8570 14170
rect 8408 14116 8432 14118
rect 8488 14116 8512 14118
rect 8568 14116 8592 14118
rect 8206 14104 8262 14113
rect 8352 14096 8648 14116
rect 8206 14039 8262 14048
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 8220 13920 8248 14039
rect 8220 13892 8432 13920
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 8220 13258 8248 13738
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8312 13433 8340 13670
rect 8298 13424 8354 13433
rect 8298 13359 8354 13368
rect 8404 13326 8432 13892
rect 8680 13462 8708 14447
rect 8668 13456 8720 13462
rect 8668 13398 8720 13404
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 7748 13252 7800 13258
rect 7748 13194 7800 13200
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 7760 12889 7788 13194
rect 8024 13184 8076 13190
rect 8772 13161 8800 14826
rect 8864 14550 8892 16186
rect 8942 15600 8998 15609
rect 8942 15535 8998 15544
rect 8956 15094 8984 15535
rect 8944 15088 8996 15094
rect 8944 15030 8996 15036
rect 8942 14648 8998 14657
rect 8942 14583 8998 14592
rect 8852 14544 8904 14550
rect 8852 14486 8904 14492
rect 8850 14104 8906 14113
rect 8850 14039 8906 14048
rect 8864 13802 8892 14039
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8864 13326 8892 13738
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8024 13126 8076 13132
rect 8206 13152 8262 13161
rect 8036 13025 8064 13126
rect 8758 13152 8814 13161
rect 8206 13087 8262 13096
rect 8022 13016 8078 13025
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7932 12980 7984 12986
rect 8022 12951 8078 12960
rect 7932 12922 7984 12928
rect 7746 12880 7802 12889
rect 7746 12815 7802 12824
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7562 11455 7618 11464
rect 7659 11478 7696 11506
rect 7659 11370 7687 11478
rect 7576 11342 7687 11370
rect 7576 10810 7604 11342
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7668 10606 7696 11222
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7668 10266 7696 10542
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7576 9042 7604 9998
rect 7654 9752 7710 9761
rect 7654 9687 7710 9696
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7470 8664 7526 8673
rect 7576 8634 7604 8842
rect 7470 8599 7526 8608
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7576 8022 7604 8570
rect 7564 8016 7616 8022
rect 7564 7958 7616 7964
rect 7668 7868 7696 9687
rect 7576 7840 7696 7868
rect 7470 7712 7526 7721
rect 7470 7647 7526 7656
rect 7484 7342 7512 7647
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7300 6582 7420 6610
rect 7194 6488 7250 6497
rect 7194 6423 7250 6432
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7208 5370 7236 6190
rect 7300 6089 7328 6582
rect 7484 6440 7512 7142
rect 7392 6412 7512 6440
rect 7286 6080 7342 6089
rect 7286 6015 7342 6024
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7300 5574 7328 5782
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7286 5400 7342 5409
rect 7196 5364 7248 5370
rect 7286 5335 7342 5344
rect 7196 5306 7248 5312
rect 7208 5234 7236 5306
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7300 4690 7328 5335
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7208 4457 7236 4626
rect 7392 4593 7420 6412
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7484 4622 7512 6258
rect 7472 4616 7524 4622
rect 7378 4584 7434 4593
rect 7472 4558 7524 4564
rect 7378 4519 7434 4528
rect 7194 4448 7250 4457
rect 7194 4383 7250 4392
rect 7116 4270 7236 4298
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 7208 3924 7236 4270
rect 7288 3936 7340 3942
rect 6918 3904 6974 3913
rect 7208 3896 7288 3924
rect 7288 3878 7340 3884
rect 6918 3839 6974 3848
rect 6932 3738 6960 3839
rect 7194 3768 7250 3777
rect 6920 3732 6972 3738
rect 7194 3703 7196 3712
rect 6920 3674 6972 3680
rect 7248 3703 7250 3712
rect 7196 3674 7248 3680
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6932 3369 6960 3470
rect 7392 3448 7420 4519
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7484 3738 7512 4218
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7392 3420 7512 3448
rect 6918 3360 6974 3369
rect 6918 3295 6974 3304
rect 7102 3360 7158 3369
rect 7102 3295 7158 3304
rect 7378 3360 7434 3369
rect 7378 3295 7434 3304
rect 7116 3074 7144 3295
rect 7024 3046 7144 3074
rect 7024 2854 7052 3046
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7010 2680 7066 2689
rect 7010 2615 7066 2624
rect 7196 2644 7248 2650
rect 6828 2372 6880 2378
rect 6828 2314 6880 2320
rect 6736 1828 6788 1834
rect 6736 1770 6788 1776
rect 6460 1430 6512 1436
rect 6564 1414 6684 1442
rect 6092 1352 6144 1358
rect 6092 1294 6144 1300
rect 6104 480 6132 1294
rect 6564 480 6592 1414
rect 7024 480 7052 2615
rect 7196 2586 7248 2592
rect 7208 1834 7236 2586
rect 7196 1828 7248 1834
rect 7196 1770 7248 1776
rect 7392 480 7420 3295
rect 7484 3194 7512 3420
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7576 2514 7604 7840
rect 7760 7528 7788 12582
rect 7852 10656 7880 12922
rect 7944 12850 7972 12922
rect 8114 12880 8170 12889
rect 7932 12844 7984 12850
rect 8114 12815 8170 12824
rect 8220 12866 8248 13087
rect 8352 13084 8648 13104
rect 8758 13087 8814 13096
rect 8408 13082 8432 13084
rect 8488 13082 8512 13084
rect 8568 13082 8592 13084
rect 8430 13030 8432 13082
rect 8494 13030 8506 13082
rect 8568 13030 8570 13082
rect 8408 13028 8432 13030
rect 8488 13028 8512 13030
rect 8568 13028 8592 13030
rect 8352 13008 8648 13028
rect 8956 13025 8984 14583
rect 9048 13734 9076 16340
rect 9140 14793 9168 17520
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9218 15464 9274 15473
rect 9218 15399 9274 15408
rect 9312 15428 9364 15434
rect 9232 15026 9260 15399
rect 9312 15370 9364 15376
rect 9324 15201 9352 15370
rect 9310 15192 9366 15201
rect 9310 15127 9366 15136
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9232 14822 9260 14962
rect 9220 14816 9272 14822
rect 9126 14784 9182 14793
rect 9220 14758 9272 14764
rect 9126 14719 9182 14728
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 13569 9076 13670
rect 9034 13560 9090 13569
rect 9140 13530 9168 13738
rect 9034 13495 9090 13504
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9036 13456 9088 13462
rect 9036 13398 9088 13404
rect 8942 13016 8998 13025
rect 8760 12980 8812 12986
rect 9048 12986 9076 13398
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 8942 12951 8998 12960
rect 9036 12980 9088 12986
rect 8760 12922 8812 12928
rect 8220 12850 8432 12866
rect 8220 12844 8444 12850
rect 8220 12838 8392 12844
rect 7932 12786 7984 12792
rect 8128 12782 8156 12815
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7944 10792 7972 12582
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 8036 10985 8064 12378
rect 8114 11928 8170 11937
rect 8114 11863 8170 11872
rect 8128 11354 8156 11863
rect 8220 11642 8248 12838
rect 8392 12786 8444 12792
rect 8772 12782 8800 12922
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8864 12458 8892 12786
rect 8956 12646 8984 12951
rect 9036 12922 9088 12928
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8864 12430 8984 12458
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8404 12170 8432 12242
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8392 12164 8444 12170
rect 8392 12106 8444 12112
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8352 11996 8648 12016
rect 8408 11994 8432 11996
rect 8488 11994 8512 11996
rect 8568 11994 8592 11996
rect 8430 11942 8432 11994
rect 8494 11942 8506 11994
rect 8568 11942 8570 11994
rect 8408 11940 8432 11942
rect 8488 11940 8512 11942
rect 8568 11940 8592 11942
rect 8352 11920 8648 11940
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8220 11614 8432 11642
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 8022 10976 8078 10985
rect 8022 10911 8078 10920
rect 8114 10840 8170 10849
rect 8024 10804 8076 10810
rect 7944 10764 8024 10792
rect 8114 10775 8170 10784
rect 8024 10746 8076 10752
rect 8128 10674 8156 10775
rect 8116 10668 8168 10674
rect 7852 10628 7972 10656
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7852 9874 7880 10474
rect 7944 10266 7972 10628
rect 8116 10610 8168 10616
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7852 9846 7972 9874
rect 7838 9752 7894 9761
rect 7838 9687 7894 9696
rect 7852 9586 7880 9687
rect 7944 9654 7972 9846
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7852 8378 7880 9318
rect 8036 9110 8064 10474
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 8024 8832 8076 8838
rect 7930 8800 7986 8809
rect 8024 8774 8076 8780
rect 7930 8735 7986 8744
rect 7944 8498 7972 8735
rect 8036 8537 8064 8774
rect 8128 8673 8156 10066
rect 8114 8664 8170 8673
rect 8114 8599 8170 8608
rect 8022 8528 8078 8537
rect 7932 8492 7984 8498
rect 8220 8480 8248 11494
rect 8404 11082 8432 11614
rect 8496 11218 8524 11698
rect 8680 11694 8708 12106
rect 8772 12073 8800 12174
rect 8852 12096 8904 12102
rect 8758 12064 8814 12073
rect 8852 12038 8904 12044
rect 8758 11999 8814 12008
rect 8864 11694 8892 12038
rect 8956 11898 8984 12430
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8944 11552 8996 11558
rect 8588 11512 8944 11540
rect 8588 11286 8616 11512
rect 8944 11494 8996 11500
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8352 10908 8648 10928
rect 8408 10906 8432 10908
rect 8488 10906 8512 10908
rect 8568 10906 8592 10908
rect 8430 10854 8432 10906
rect 8494 10854 8506 10906
rect 8568 10854 8570 10906
rect 8408 10852 8432 10854
rect 8488 10852 8512 10854
rect 8568 10852 8592 10854
rect 8352 10832 8648 10852
rect 8680 10538 8708 11086
rect 8850 10976 8906 10985
rect 8850 10911 8906 10920
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 10130 8340 10406
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8404 10130 8432 10202
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8352 9820 8648 9840
rect 8408 9818 8432 9820
rect 8488 9818 8512 9820
rect 8568 9818 8592 9820
rect 8430 9766 8432 9818
rect 8494 9766 8506 9818
rect 8568 9766 8570 9818
rect 8408 9764 8432 9766
rect 8488 9764 8512 9766
rect 8568 9764 8592 9766
rect 8352 9744 8648 9764
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8312 9110 8340 9590
rect 8588 9518 8616 9590
rect 8680 9518 8708 10202
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8312 8820 8340 9046
rect 8760 8968 8812 8974
rect 8758 8936 8760 8945
rect 8812 8936 8814 8945
rect 8758 8871 8814 8880
rect 8288 8792 8340 8820
rect 8760 8832 8812 8838
rect 8288 8566 8316 8792
rect 8760 8774 8812 8780
rect 8763 8758 8800 8774
rect 8352 8732 8648 8752
rect 8408 8730 8432 8732
rect 8488 8730 8512 8732
rect 8568 8730 8592 8732
rect 8430 8678 8432 8730
rect 8494 8678 8506 8730
rect 8568 8678 8570 8730
rect 8408 8676 8432 8678
rect 8488 8676 8512 8678
rect 8568 8676 8592 8678
rect 8352 8656 8648 8676
rect 8288 8560 8352 8566
rect 8288 8520 8300 8560
rect 8763 8514 8791 8758
rect 8300 8502 8352 8508
rect 8022 8463 8078 8472
rect 7932 8434 7984 8440
rect 8128 8452 8248 8480
rect 8588 8486 8791 8514
rect 7852 8350 7972 8378
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7852 8022 7880 8230
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 7944 7528 7972 8350
rect 8022 7712 8078 7721
rect 8022 7647 8078 7656
rect 7729 7500 7788 7528
rect 7852 7500 7972 7528
rect 7729 7290 7757 7500
rect 7729 7262 7788 7290
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7668 6390 7696 6870
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7668 3670 7696 6190
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7760 2650 7788 7262
rect 7852 6254 7880 7500
rect 8036 7460 8064 7647
rect 8128 7528 8156 8452
rect 8484 8424 8536 8430
rect 8588 8412 8616 8486
rect 8536 8384 8616 8412
rect 8668 8424 8720 8430
rect 8484 8366 8536 8372
rect 8668 8366 8720 8372
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8220 7721 8248 8298
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8588 7886 8616 7958
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8206 7712 8262 7721
rect 8206 7647 8262 7656
rect 8352 7644 8648 7664
rect 8408 7642 8432 7644
rect 8488 7642 8512 7644
rect 8568 7642 8592 7644
rect 8430 7590 8432 7642
rect 8494 7590 8506 7642
rect 8568 7590 8570 7642
rect 8408 7588 8432 7590
rect 8488 7588 8512 7590
rect 8568 7588 8592 7590
rect 8352 7568 8648 7588
rect 8128 7500 8340 7528
rect 8036 7432 8156 7460
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7935 7262 7972 7278
rect 7944 7177 7972 7262
rect 7930 7168 7986 7177
rect 7930 7103 7986 7112
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7838 6080 7894 6089
rect 7838 6015 7894 6024
rect 7852 5846 7880 6015
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7944 5710 7972 6802
rect 8036 6322 8064 7278
rect 8128 7206 8156 7432
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8312 7018 8340 7500
rect 8680 7342 8708 8366
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8390 7168 8446 7177
rect 8390 7103 8446 7112
rect 8666 7168 8722 7177
rect 8666 7103 8722 7112
rect 8128 6990 8340 7018
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8128 6202 8156 6990
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8312 6769 8340 6870
rect 8404 6798 8432 7103
rect 8392 6792 8444 6798
rect 8298 6760 8354 6769
rect 8392 6734 8444 6740
rect 8482 6760 8538 6769
rect 8298 6695 8354 6704
rect 8482 6695 8538 6704
rect 8496 6644 8524 6695
rect 8220 6616 8524 6644
rect 8220 6497 8248 6616
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8206 6488 8262 6497
rect 8352 6480 8648 6500
rect 8680 6440 8708 7103
rect 8206 6423 8262 6432
rect 8036 6174 8156 6202
rect 8496 6412 8708 6440
rect 8300 6180 8352 6186
rect 8036 6066 8064 6174
rect 8300 6122 8352 6128
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8116 6112 8168 6118
rect 8027 6038 8064 6066
rect 8097 6060 8116 6066
rect 8208 6112 8260 6118
rect 8097 6054 8168 6060
rect 8206 6080 8208 6089
rect 8260 6080 8262 6089
rect 8097 6038 8156 6054
rect 8027 5828 8055 6038
rect 8097 5846 8125 6038
rect 8206 6015 8262 6024
rect 8097 5840 8168 5846
rect 8027 5800 8064 5828
rect 8097 5800 8116 5840
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7852 4060 7880 5510
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7944 4214 7972 4422
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7932 4072 7984 4078
rect 7852 4032 7932 4060
rect 7932 4014 7984 4020
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 7852 3126 7880 3538
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7838 2816 7894 2825
rect 7838 2751 7894 2760
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7576 2281 7604 2314
rect 7562 2272 7618 2281
rect 7562 2207 7618 2216
rect 7852 480 7880 2751
rect 7944 2417 7972 2994
rect 7930 2408 7986 2417
rect 7930 2343 7986 2352
rect 8036 1358 8064 5800
rect 8116 5782 8168 5788
rect 8312 5760 8340 6122
rect 8404 5914 8432 6122
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8392 5772 8444 5778
rect 8312 5732 8392 5760
rect 8392 5714 8444 5720
rect 8496 5658 8524 6412
rect 8574 6080 8630 6089
rect 8574 6015 8630 6024
rect 8588 5914 8616 6015
rect 8576 5908 8628 5914
rect 8772 5896 8800 7686
rect 8576 5850 8628 5856
rect 8680 5868 8800 5896
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8128 5630 8524 5658
rect 8128 5409 8156 5630
rect 8208 5568 8260 5574
rect 8588 5556 8616 5714
rect 8260 5528 8616 5556
rect 8208 5510 8260 5516
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8114 5400 8170 5409
rect 8352 5392 8648 5412
rect 8114 5335 8170 5344
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 8116 4480 8168 4486
rect 8114 4448 8116 4457
rect 8168 4448 8170 4457
rect 8114 4383 8170 4392
rect 8114 4312 8170 4321
rect 8114 4247 8170 4256
rect 8128 3602 8156 4247
rect 8220 4146 8248 5034
rect 8352 4380 8648 4400
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 8680 4282 8708 5868
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8772 4622 8800 5714
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 8772 4214 8800 4422
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8128 1426 8156 3538
rect 8220 3516 8248 4082
rect 8760 3936 8812 3942
rect 8588 3896 8760 3924
rect 8392 3528 8444 3534
rect 8220 3488 8392 3516
rect 8392 3470 8444 3476
rect 8588 3466 8616 3896
rect 8760 3878 8812 3884
rect 8864 3482 8892 10911
rect 8944 9988 8996 9994
rect 8944 9930 8996 9936
rect 8956 8956 8984 9930
rect 9048 9518 9076 12650
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8925 8928 8984 8956
rect 8925 8786 8953 8928
rect 8925 8758 8984 8786
rect 8956 7750 8984 8758
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 9034 7712 9090 7721
rect 9034 7647 9090 7656
rect 8942 7576 8998 7585
rect 8942 7511 8998 7520
rect 8956 6934 8984 7511
rect 9048 6934 9076 7647
rect 9140 7426 9168 13194
rect 9232 11898 9260 14282
rect 9324 14113 9352 15127
rect 9310 14104 9366 14113
rect 9310 14039 9366 14048
rect 9310 13424 9366 13433
rect 9310 13359 9366 13368
rect 9324 12850 9352 13359
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9310 12472 9366 12481
rect 9310 12407 9366 12416
rect 9324 12102 9352 12407
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9232 11354 9260 11834
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9324 11286 9352 11698
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10266 9260 10950
rect 9310 10840 9366 10849
rect 9310 10775 9366 10784
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9218 9208 9274 9217
rect 9218 9143 9274 9152
rect 9232 8945 9260 9143
rect 9218 8936 9274 8945
rect 9218 8871 9274 8880
rect 9324 8265 9352 10775
rect 9310 8256 9366 8265
rect 9310 8191 9366 8200
rect 9140 7398 9352 7426
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 9036 6928 9088 6934
rect 9036 6870 9088 6876
rect 8942 6488 8998 6497
rect 8942 6423 8998 6432
rect 8956 6089 8984 6423
rect 9048 6322 9076 6870
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8942 6080 8998 6089
rect 8942 6015 8998 6024
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8956 4554 8984 5646
rect 9048 5574 9076 5714
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 8944 4548 8996 4554
rect 8944 4490 8996 4496
rect 8942 4448 8998 4457
rect 8942 4383 8998 4392
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8680 3454 8892 3482
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8206 3224 8262 3233
rect 8352 3216 8648 3236
rect 8206 3159 8262 3168
rect 8220 3074 8248 3159
rect 8220 3046 8524 3074
rect 8496 2990 8524 3046
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8206 2680 8262 2689
rect 8206 2615 8262 2624
rect 8116 1420 8168 1426
rect 8116 1362 8168 1368
rect 8024 1352 8076 1358
rect 8024 1294 8076 1300
rect 8220 480 8248 2615
rect 8404 2378 8432 2926
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8588 2689 8616 2790
rect 8574 2680 8630 2689
rect 8574 2615 8630 2624
rect 8680 2582 8708 3454
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8864 2650 8892 3334
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 8668 2576 8720 2582
rect 8772 2553 8800 2586
rect 8668 2518 8720 2524
rect 8758 2544 8814 2553
rect 8956 2514 8984 4383
rect 9034 4312 9090 4321
rect 9034 4247 9090 4256
rect 9048 3738 9076 4247
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9140 3194 9168 6326
rect 9232 5250 9260 6734
rect 9324 6390 9352 7398
rect 9416 6905 9444 15982
rect 9508 14657 9536 17520
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9494 14648 9550 14657
rect 9494 14583 9550 14592
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9508 12714 9536 13466
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9508 8888 9536 12650
rect 9600 11098 9628 15574
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 14521 9720 15506
rect 9968 14600 9996 17520
rect 10324 16380 10376 16386
rect 10324 16322 10376 16328
rect 10140 16312 10192 16318
rect 10140 16254 10192 16260
rect 9876 14572 9996 14600
rect 9678 14512 9734 14521
rect 9678 14447 9734 14456
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9692 13462 9720 14350
rect 9876 14249 9904 14572
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9862 14240 9918 14249
rect 9862 14175 9918 14184
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 9692 12238 9720 13398
rect 9784 12306 9812 13874
rect 9876 13569 9904 13942
rect 9862 13560 9918 13569
rect 9862 13495 9918 13504
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9876 13326 9904 13398
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9876 13025 9904 13126
rect 9862 13016 9918 13025
rect 9968 12986 9996 14418
rect 9862 12951 9918 12960
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9772 12300 9824 12306
rect 9968 12288 9996 12922
rect 10060 12850 10088 14486
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 9772 12242 9824 12248
rect 9876 12260 9996 12288
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 11694 9720 12038
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 11354 9720 11494
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9876 11218 9904 12260
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9600 11082 9812 11098
rect 9600 11076 9824 11082
rect 9600 11070 9772 11076
rect 9772 11018 9824 11024
rect 9770 10976 9826 10985
rect 9770 10911 9826 10920
rect 9586 10840 9642 10849
rect 9586 10775 9642 10784
rect 9600 8956 9628 10775
rect 9680 10736 9732 10742
rect 9678 10704 9680 10713
rect 9732 10704 9734 10713
rect 9678 10639 9734 10648
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9692 10062 9720 10474
rect 9784 10418 9812 10911
rect 9876 10674 9904 11154
rect 9968 10810 9996 11494
rect 10060 11286 10088 12582
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 10152 10606 10180 16254
rect 10336 15706 10364 16322
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10244 13258 10272 14418
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10336 12594 10364 14894
rect 10428 14793 10456 17520
rect 10796 15892 10824 17520
rect 11256 16318 11284 17520
rect 11244 16312 11296 16318
rect 11244 16254 11296 16260
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11518 16008 11574 16017
rect 10612 15864 10824 15892
rect 10508 14952 10560 14958
rect 10508 14894 10560 14900
rect 10414 14784 10470 14793
rect 10414 14719 10470 14728
rect 10414 14648 10470 14657
rect 10414 14583 10470 14592
rect 10428 12646 10456 14583
rect 10520 14482 10548 14894
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10520 13569 10548 14010
rect 10506 13560 10562 13569
rect 10506 13495 10562 13504
rect 10506 13424 10562 13433
rect 10506 13359 10508 13368
rect 10560 13359 10562 13368
rect 10508 13330 10560 13336
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10244 12566 10364 12594
rect 10416 12640 10468 12646
rect 10520 12617 10548 12718
rect 10416 12582 10468 12588
rect 10506 12608 10562 12617
rect 10244 10810 10272 12566
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10336 11626 10364 11834
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10428 10690 10456 12582
rect 10506 12543 10562 12552
rect 10612 11778 10640 15864
rect 10817 15804 11113 15824
rect 10873 15802 10897 15804
rect 10953 15802 10977 15804
rect 11033 15802 11057 15804
rect 10895 15750 10897 15802
rect 10959 15750 10971 15802
rect 11033 15750 11035 15802
rect 10873 15748 10897 15750
rect 10953 15748 10977 15750
rect 11033 15748 11057 15750
rect 10817 15728 11113 15748
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 11164 14890 11192 15098
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10704 14278 10732 14758
rect 10817 14716 11113 14736
rect 10873 14714 10897 14716
rect 10953 14714 10977 14716
rect 11033 14714 11057 14716
rect 10895 14662 10897 14714
rect 10959 14662 10971 14714
rect 11033 14662 11035 14714
rect 10873 14660 10897 14662
rect 10953 14660 10977 14662
rect 11033 14660 11057 14662
rect 10817 14640 11113 14660
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 11256 13938 11284 15302
rect 11348 14498 11376 15982
rect 11518 15943 11574 15952
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11440 14618 11468 14758
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11348 14470 11468 14498
rect 11440 14278 11468 14470
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 11244 13728 11296 13734
rect 11242 13696 11244 13705
rect 11296 13696 11298 13705
rect 10817 13628 11113 13648
rect 11242 13631 11298 13640
rect 10873 13626 10897 13628
rect 10953 13626 10977 13628
rect 11033 13626 11057 13628
rect 10895 13574 10897 13626
rect 10959 13574 10971 13626
rect 11033 13574 11035 13626
rect 10873 13572 10897 13574
rect 10953 13572 10977 13574
rect 11033 13572 11057 13574
rect 10817 13552 11113 13572
rect 11256 13025 11284 13631
rect 11348 13308 11376 14214
rect 11428 13320 11480 13326
rect 11348 13280 11428 13308
rect 11428 13262 11480 13268
rect 11532 13172 11560 15943
rect 11624 13569 11652 17520
rect 12084 15688 12112 17520
rect 11900 15660 12112 15688
rect 11702 15192 11758 15201
rect 11702 15127 11758 15136
rect 11716 15026 11744 15127
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11796 14816 11848 14822
rect 11794 14784 11796 14793
rect 11848 14784 11850 14793
rect 11794 14719 11850 14728
rect 11808 14550 11836 14719
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11900 13818 11928 15660
rect 12164 15632 12216 15638
rect 12164 15574 12216 15580
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 11992 14346 12020 15506
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 12084 14482 12112 14826
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 12070 14240 12126 14249
rect 12070 14175 12126 14184
rect 11808 13790 11928 13818
rect 11610 13560 11666 13569
rect 11610 13495 11666 13504
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11440 13144 11560 13172
rect 11242 13016 11298 13025
rect 11242 12951 11298 12960
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 10817 12540 11113 12560
rect 10873 12538 10897 12540
rect 10953 12538 10977 12540
rect 11033 12538 11057 12540
rect 10895 12486 10897 12538
rect 10959 12486 10971 12538
rect 11033 12486 11035 12538
rect 10873 12484 10897 12486
rect 10953 12484 10977 12486
rect 11033 12484 11057 12486
rect 10817 12464 11113 12484
rect 10968 12232 11020 12238
rect 10782 12200 10838 12209
rect 10968 12174 11020 12180
rect 10782 12135 10838 12144
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10336 10662 10456 10690
rect 10520 11750 10640 11778
rect 10140 10600 10192 10606
rect 9968 10560 10140 10588
rect 9784 10390 9904 10418
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9784 9761 9812 10134
rect 9770 9752 9826 9761
rect 9770 9687 9826 9696
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9692 9382 9720 9590
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9784 9110 9812 9386
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9600 8928 9812 8956
rect 9508 8860 9720 8888
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9600 7954 9628 8230
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9692 7834 9720 8860
rect 9784 8265 9812 8928
rect 9770 8256 9826 8265
rect 9770 8191 9826 8200
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9600 7806 9720 7834
rect 9508 7342 9536 7754
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9402 6896 9458 6905
rect 9402 6831 9458 6840
rect 9416 6497 9444 6831
rect 9508 6798 9536 7278
rect 9600 7177 9628 7806
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9586 7168 9642 7177
rect 9586 7103 9642 7112
rect 9586 7032 9642 7041
rect 9692 7018 9720 7414
rect 9784 7206 9812 8026
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9642 6990 9720 7018
rect 9784 7002 9812 7142
rect 9876 7041 9904 10390
rect 9862 7032 9918 7041
rect 9772 6996 9824 7002
rect 9586 6967 9642 6976
rect 9862 6967 9918 6976
rect 9772 6938 9824 6944
rect 9968 6916 9996 10560
rect 10140 10542 10192 10548
rect 10336 10198 10364 10662
rect 10416 10600 10468 10606
rect 10414 10568 10416 10577
rect 10468 10568 10470 10577
rect 10414 10503 10470 10512
rect 10520 10266 10548 11750
rect 10704 11608 10732 12038
rect 10612 11580 10732 11608
rect 10612 11529 10640 11580
rect 10796 11540 10824 12135
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10888 11830 10916 12038
rect 10876 11824 10928 11830
rect 10876 11766 10928 11772
rect 10980 11694 11008 12174
rect 11256 12170 11284 12718
rect 11348 12442 11376 12786
rect 11440 12442 11468 13144
rect 11624 12986 11652 13398
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11532 12714 11560 12854
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11716 12594 11744 13330
rect 11624 12566 11744 12594
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11624 12238 11652 12566
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11334 12064 11390 12073
rect 11334 11999 11390 12008
rect 11152 11824 11204 11830
rect 11072 11772 11152 11778
rect 11072 11766 11204 11772
rect 11072 11762 11192 11766
rect 11060 11756 11192 11762
rect 11112 11750 11192 11756
rect 11060 11698 11112 11704
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10598 11520 10654 11529
rect 10598 11455 10654 11464
rect 10704 11512 10824 11540
rect 10704 11121 10732 11512
rect 10817 11452 11113 11472
rect 10873 11450 10897 11452
rect 10953 11450 10977 11452
rect 11033 11450 11057 11452
rect 10895 11398 10897 11450
rect 10959 11398 10971 11450
rect 11033 11398 11035 11450
rect 10873 11396 10897 11398
rect 10953 11396 10977 11398
rect 11033 11396 11057 11398
rect 10817 11376 11113 11396
rect 10690 11112 10746 11121
rect 10690 11047 10746 11056
rect 10598 10976 10654 10985
rect 10598 10911 10654 10920
rect 10612 10305 10640 10911
rect 11164 10826 11192 11630
rect 11348 11626 11376 11999
rect 11624 11898 11652 12174
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11520 11824 11572 11830
rect 11520 11766 11572 11772
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 11532 11286 11560 11766
rect 11612 11756 11664 11762
rect 11808 11744 11836 13790
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11612 11698 11664 11704
rect 11716 11716 11836 11744
rect 11624 11354 11652 11698
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11520 11280 11572 11286
rect 11242 11248 11298 11257
rect 11716 11234 11744 11716
rect 11900 11676 11928 13670
rect 11978 13288 12034 13297
rect 11978 13223 11980 13232
rect 12032 13223 12034 13232
rect 11980 13194 12032 13200
rect 12084 12628 12112 14175
rect 12176 13705 12204 15574
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12268 13734 12296 15370
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12360 14521 12388 14894
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12346 14512 12402 14521
rect 12346 14447 12402 14456
rect 12346 14104 12402 14113
rect 12346 14039 12402 14048
rect 12256 13728 12308 13734
rect 12162 13696 12218 13705
rect 12256 13670 12308 13676
rect 12162 13631 12218 13640
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 11520 11222 11572 11228
rect 11242 11183 11298 11192
rect 11336 11212 11388 11218
rect 11256 11082 11284 11183
rect 11336 11154 11388 11160
rect 11624 11206 11744 11234
rect 11808 11648 11928 11676
rect 11992 12600 12112 12628
rect 12164 12640 12216 12646
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 10692 10804 10744 10810
rect 11164 10798 11284 10826
rect 10692 10746 10744 10752
rect 10598 10296 10654 10305
rect 10508 10260 10560 10266
rect 10598 10231 10654 10240
rect 10508 10202 10560 10208
rect 10324 10192 10376 10198
rect 10324 10134 10376 10140
rect 10414 10160 10470 10169
rect 10048 10124 10100 10130
rect 10520 10130 10548 10202
rect 10598 10160 10654 10169
rect 10414 10095 10470 10104
rect 10508 10124 10560 10130
rect 10048 10066 10100 10072
rect 10060 9926 10088 10066
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 10428 9874 10456 10095
rect 10704 10130 10732 10746
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10796 10538 10824 10610
rect 10784 10532 10836 10538
rect 10784 10474 10836 10480
rect 10817 10364 11113 10384
rect 10873 10362 10897 10364
rect 10953 10362 10977 10364
rect 11033 10362 11057 10364
rect 10895 10310 10897 10362
rect 10959 10310 10971 10362
rect 11033 10310 11035 10362
rect 10873 10308 10897 10310
rect 10953 10308 10977 10310
rect 11033 10308 11057 10310
rect 10817 10288 11113 10308
rect 10598 10095 10654 10104
rect 10692 10124 10744 10130
rect 10508 10066 10560 10072
rect 10612 9994 10640 10095
rect 10692 10066 10744 10072
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10428 9846 10640 9874
rect 10138 9752 10194 9761
rect 10138 9687 10194 9696
rect 10322 9752 10378 9761
rect 10322 9687 10378 9696
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 10060 8430 10088 9454
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 9959 6888 9996 6916
rect 10060 6916 10088 7278
rect 10152 7206 10180 9687
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10244 8090 10272 9522
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10244 7313 10272 7346
rect 10230 7304 10286 7313
rect 10230 7239 10286 7248
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10060 6888 10272 6916
rect 9772 6860 9824 6866
rect 9959 6848 9987 6888
rect 9959 6820 10088 6848
rect 9772 6802 9824 6808
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9402 6488 9458 6497
rect 9402 6423 9458 6432
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9310 5808 9366 5817
rect 9310 5743 9366 5752
rect 9324 5409 9352 5743
rect 9310 5400 9366 5409
rect 9310 5335 9366 5344
rect 9232 5222 9352 5250
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9232 3534 9260 5102
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9218 3360 9274 3369
rect 9218 3295 9274 3304
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8758 2479 8814 2488
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 8668 1828 8720 1834
rect 8668 1770 8720 1776
rect 8680 480 8708 1770
rect 8772 1698 8800 2382
rect 8760 1692 8812 1698
rect 8760 1634 8812 1640
rect 9048 1601 9076 2994
rect 9232 2990 9260 3295
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9324 2922 9352 5222
rect 9312 2916 9364 2922
rect 9312 2858 9364 2864
rect 9324 2281 9352 2858
rect 9310 2272 9366 2281
rect 9310 2207 9366 2216
rect 9034 1592 9090 1601
rect 9034 1527 9090 1536
rect 9416 1408 9444 6258
rect 9508 5710 9536 6734
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9600 6458 9628 6598
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9508 5250 9536 5646
rect 9600 5370 9628 6394
rect 9784 6390 9812 6802
rect 10060 6769 10088 6820
rect 10046 6760 10102 6769
rect 10046 6695 10102 6704
rect 9954 6624 10010 6633
rect 9954 6559 10010 6568
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9968 6186 9996 6559
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 9968 5778 9996 6122
rect 10060 5953 10088 6695
rect 10244 6458 10272 6888
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10046 5944 10102 5953
rect 10046 5879 10102 5888
rect 10152 5846 10180 6054
rect 10230 5944 10286 5953
rect 10230 5879 10286 5888
rect 10140 5840 10192 5846
rect 10046 5808 10102 5817
rect 9772 5772 9824 5778
rect 9956 5772 10008 5778
rect 9824 5732 9904 5760
rect 9772 5714 9824 5720
rect 9770 5536 9826 5545
rect 9770 5471 9826 5480
rect 9678 5400 9734 5409
rect 9588 5364 9640 5370
rect 9678 5335 9680 5344
rect 9588 5306 9640 5312
rect 9732 5335 9734 5344
rect 9680 5306 9732 5312
rect 9508 5222 9628 5250
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9508 4282 9536 4966
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9508 3602 9536 4014
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9508 2310 9536 3402
rect 9600 3194 9628 5222
rect 9784 5137 9812 5471
rect 9770 5128 9826 5137
rect 9770 5063 9826 5072
rect 9678 4856 9734 4865
rect 9678 4791 9734 4800
rect 9692 4690 9720 4791
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9784 4486 9812 4558
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9692 3670 9720 4422
rect 9876 4078 9904 5732
rect 10140 5782 10192 5788
rect 10046 5743 10102 5752
rect 9956 5714 10008 5720
rect 9954 5400 10010 5409
rect 9954 5335 10010 5344
rect 9968 5234 9996 5335
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9968 4554 9996 5170
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9692 1630 9720 3470
rect 9784 3466 9812 3538
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9876 2990 9904 4014
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9968 3505 9996 3946
rect 9954 3496 10010 3505
rect 9954 3431 10010 3440
rect 10060 3380 10088 5743
rect 10138 4312 10194 4321
rect 10138 4247 10194 4256
rect 9968 3352 10088 3380
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9876 2650 9904 2790
rect 9968 2689 9996 3352
rect 10152 2922 10180 4247
rect 10244 3942 10272 5879
rect 10336 5234 10364 9687
rect 10414 9616 10470 9625
rect 10470 9574 10548 9602
rect 10612 9586 10640 9846
rect 10414 9551 10470 9560
rect 10416 9376 10468 9382
rect 10520 9364 10548 9574
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10600 9376 10652 9382
rect 10520 9336 10600 9364
rect 10416 9318 10468 9324
rect 10600 9318 10652 9324
rect 10428 9024 10456 9318
rect 10508 9036 10560 9042
rect 10428 8996 10508 9024
rect 10508 8978 10560 8984
rect 10598 8936 10654 8945
rect 10416 8900 10468 8906
rect 10598 8871 10654 8880
rect 10416 8842 10468 8848
rect 10428 8634 10456 8842
rect 10612 8634 10640 8871
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10704 8514 10732 10066
rect 11164 10062 11192 10678
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 10817 9276 11113 9296
rect 10873 9274 10897 9276
rect 10953 9274 10977 9276
rect 11033 9274 11057 9276
rect 10895 9222 10897 9274
rect 10959 9222 10971 9274
rect 11033 9222 11035 9274
rect 10873 9220 10897 9222
rect 10953 9220 10977 9222
rect 11033 9220 11057 9222
rect 10817 9200 11113 9220
rect 11164 9160 11192 9590
rect 10980 9132 11192 9160
rect 10980 8566 11008 9132
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11072 8945 11100 8978
rect 11058 8936 11114 8945
rect 11058 8871 11114 8880
rect 10612 8486 10732 8514
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10784 8492 10836 8498
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10428 7342 10456 8298
rect 10612 8090 10640 8486
rect 10784 8434 10836 8440
rect 10692 8288 10744 8294
rect 10796 8276 10824 8434
rect 11058 8392 11114 8401
rect 11058 8327 11060 8336
rect 11112 8327 11114 8336
rect 11060 8298 11112 8304
rect 10744 8248 10824 8276
rect 10692 8230 10744 8236
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10508 7948 10560 7954
rect 10560 7908 10640 7936
rect 10508 7890 10560 7896
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10428 6866 10456 7142
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10428 4758 10456 6802
rect 10520 6458 10548 7346
rect 10612 7002 10640 7908
rect 10704 7886 10732 8230
rect 10817 8188 11113 8208
rect 10873 8186 10897 8188
rect 10953 8186 10977 8188
rect 11033 8186 11057 8188
rect 10895 8134 10897 8186
rect 10959 8134 10971 8186
rect 11033 8134 11035 8186
rect 10873 8132 10897 8134
rect 10953 8132 10977 8134
rect 11033 8132 11057 8134
rect 10817 8112 11113 8132
rect 11164 8090 11192 8978
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 7410 10732 7822
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11072 7449 11100 7482
rect 11058 7440 11114 7449
rect 10692 7404 10744 7410
rect 11058 7375 11114 7384
rect 10692 7346 10744 7352
rect 11164 7274 11192 7686
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 10817 7100 11113 7120
rect 10873 7098 10897 7100
rect 10953 7098 10977 7100
rect 11033 7098 11057 7100
rect 10895 7046 10897 7098
rect 10959 7046 10971 7098
rect 11033 7046 11035 7098
rect 10873 7044 10897 7046
rect 10953 7044 10977 7046
rect 11033 7044 11057 7046
rect 10817 7024 11113 7044
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 11164 6866 11192 7210
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10598 6488 10654 6497
rect 10508 6452 10560 6458
rect 10598 6423 10654 6432
rect 10508 6394 10560 6400
rect 10612 6186 10640 6423
rect 10704 6322 10732 6734
rect 11072 6440 11100 6802
rect 11152 6452 11204 6458
rect 11072 6412 11152 6440
rect 11152 6394 11204 6400
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10796 6202 10824 6258
rect 10600 6180 10652 6186
rect 10600 6122 10652 6128
rect 10704 6174 10824 6202
rect 11152 6180 11204 6186
rect 10508 6112 10560 6118
rect 10506 6080 10508 6089
rect 10560 6080 10562 6089
rect 10704 6066 10732 6174
rect 11152 6122 11204 6128
rect 10506 6015 10562 6024
rect 10612 6038 10732 6066
rect 10506 5672 10562 5681
rect 10506 5607 10562 5616
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10336 4214 10364 4626
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10428 3777 10456 4218
rect 10520 4146 10548 5607
rect 10612 4865 10640 6038
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 11164 5896 11192 6122
rect 11256 6089 11284 10798
rect 11348 10248 11376 11154
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11532 10577 11560 10610
rect 11518 10568 11574 10577
rect 11518 10503 11574 10512
rect 11428 10464 11480 10470
rect 11426 10432 11428 10441
rect 11480 10432 11482 10441
rect 11426 10367 11482 10376
rect 11348 10220 11560 10248
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11440 9722 11468 9998
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11428 9376 11480 9382
rect 11334 9344 11390 9353
rect 11428 9318 11480 9324
rect 11334 9279 11390 9288
rect 11348 9042 11376 9279
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11440 8922 11468 9318
rect 11348 8906 11468 8922
rect 11336 8900 11468 8906
rect 11388 8894 11468 8900
rect 11336 8842 11388 8848
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11334 8392 11390 8401
rect 11334 8327 11390 8336
rect 11242 6080 11298 6089
rect 11242 6015 11298 6024
rect 11164 5868 11284 5896
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11072 5681 11100 5782
rect 11058 5672 11114 5681
rect 11058 5607 11114 5616
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 11152 5568 11204 5574
rect 11256 5556 11284 5868
rect 11204 5528 11284 5556
rect 11152 5510 11204 5516
rect 10874 5400 10930 5409
rect 10874 5335 10876 5344
rect 10928 5335 10930 5344
rect 10876 5306 10928 5312
rect 10980 5234 11008 5510
rect 11150 5400 11206 5409
rect 11150 5335 11206 5344
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10598 4856 10654 4865
rect 10817 4848 11113 4868
rect 10598 4791 10654 4800
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10508 3936 10560 3942
rect 10506 3904 10508 3913
rect 10560 3904 10562 3913
rect 10506 3839 10562 3848
rect 10414 3768 10470 3777
rect 10324 3732 10376 3738
rect 10414 3703 10470 3712
rect 10324 3674 10376 3680
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10244 3194 10272 3470
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10140 2916 10192 2922
rect 10140 2858 10192 2864
rect 10046 2816 10102 2825
rect 10046 2751 10102 2760
rect 9954 2680 10010 2689
rect 9864 2644 9916 2650
rect 9954 2615 10010 2624
rect 9864 2586 9916 2592
rect 10060 2564 10088 2751
rect 9968 2536 10088 2564
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9784 1902 9812 2246
rect 9772 1896 9824 1902
rect 9772 1838 9824 1844
rect 9680 1624 9732 1630
rect 9680 1566 9732 1572
rect 9496 1420 9548 1426
rect 9416 1380 9496 1408
rect 9496 1362 9548 1368
rect 9128 876 9180 882
rect 9128 818 9180 824
rect 9140 480 9168 818
rect 9508 480 9536 1362
rect 9968 480 9996 2536
rect 10152 2310 10180 2858
rect 10244 2825 10272 3130
rect 10336 2922 10364 3674
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10230 2816 10286 2825
rect 10230 2751 10286 2760
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10336 1902 10364 2858
rect 10428 2446 10456 3606
rect 10612 3398 10640 4791
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10704 3058 10732 4422
rect 10888 4010 10916 4490
rect 10980 4010 11008 4694
rect 11164 4690 11192 5335
rect 11242 4992 11298 5001
rect 11242 4927 11298 4936
rect 11256 4826 11284 4927
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11150 4312 11206 4321
rect 11150 4247 11206 4256
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 11164 3641 11192 4247
rect 11256 4214 11284 4558
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11348 3942 11376 8327
rect 11440 6662 11468 8570
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11440 5409 11468 6190
rect 11426 5400 11482 5409
rect 11426 5335 11482 5344
rect 11428 5296 11480 5302
rect 11428 5238 11480 5244
rect 11440 4593 11468 5238
rect 11426 4584 11482 4593
rect 11426 4519 11482 4528
rect 11532 4264 11560 10220
rect 11624 9908 11652 11206
rect 11624 9880 11744 9908
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11624 8498 11652 9114
rect 11716 9110 11744 9880
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11610 8256 11666 8265
rect 11610 8191 11666 8200
rect 11624 8090 11652 8191
rect 11702 8120 11758 8129
rect 11612 8084 11664 8090
rect 11702 8055 11758 8064
rect 11612 8026 11664 8032
rect 11610 7848 11666 7857
rect 11610 7783 11666 7792
rect 11624 7750 11652 7783
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11612 7336 11664 7342
rect 11610 7304 11612 7313
rect 11664 7304 11666 7313
rect 11610 7239 11666 7248
rect 11716 7154 11744 8055
rect 11624 7126 11744 7154
rect 11624 4282 11652 7126
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11716 5234 11744 6666
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11808 5098 11836 11648
rect 11886 11248 11942 11257
rect 11886 11183 11942 11192
rect 11900 9450 11928 11183
rect 11992 11150 12020 12600
rect 12164 12582 12216 12588
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11978 10840 12034 10849
rect 11978 10775 12034 10784
rect 11992 10470 12020 10775
rect 12084 10742 12112 12038
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11992 9897 12020 10202
rect 11978 9888 12034 9897
rect 11978 9823 12034 9832
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11900 8809 11928 9386
rect 11978 9208 12034 9217
rect 12084 9194 12112 10474
rect 12176 9518 12204 12582
rect 12268 12306 12296 13262
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12268 11218 12296 12242
rect 12360 11257 12388 14039
rect 12452 13705 12480 14758
rect 12438 13696 12494 13705
rect 12438 13631 12494 13640
rect 12544 13530 12572 17520
rect 12912 16153 12940 17520
rect 12898 16144 12954 16153
rect 12624 16108 12676 16114
rect 12898 16079 12954 16088
rect 12624 16050 12676 16056
rect 12636 15570 12664 16050
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12912 15638 12940 15914
rect 12900 15632 12952 15638
rect 12900 15574 12952 15580
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 13372 15348 13400 17520
rect 13728 16176 13780 16182
rect 13728 16118 13780 16124
rect 13740 15706 13768 16118
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13634 15600 13690 15609
rect 13634 15535 13690 15544
rect 13648 15366 13676 15535
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13188 15320 13400 15348
rect 13636 15360 13688 15366
rect 13188 15065 13216 15320
rect 13636 15302 13688 15308
rect 13282 15260 13578 15280
rect 13338 15258 13362 15260
rect 13418 15258 13442 15260
rect 13498 15258 13522 15260
rect 13360 15206 13362 15258
rect 13424 15206 13436 15258
rect 13498 15206 13500 15258
rect 13338 15204 13362 15206
rect 13418 15204 13442 15206
rect 13498 15204 13522 15206
rect 13282 15184 13578 15204
rect 13544 15088 13596 15094
rect 13174 15056 13230 15065
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 13084 15020 13136 15026
rect 13544 15030 13596 15036
rect 13174 14991 13230 15000
rect 13084 14962 13136 14968
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12544 13297 12572 13466
rect 12530 13288 12586 13297
rect 12530 13223 12586 13232
rect 12438 13152 12494 13161
rect 12438 13087 12494 13096
rect 12452 12442 12480 13087
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12544 12782 12572 12854
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12452 12073 12480 12378
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12438 12064 12494 12073
rect 12438 11999 12494 12008
rect 12438 11656 12494 11665
rect 12544 11626 12572 12174
rect 12438 11591 12494 11600
rect 12532 11620 12584 11626
rect 12452 11558 12480 11591
rect 12532 11562 12584 11568
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12346 11248 12402 11257
rect 12256 11212 12308 11218
rect 12636 11234 12664 14758
rect 12806 14512 12862 14521
rect 12806 14447 12862 14456
rect 12820 14414 12848 14447
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12728 14006 12756 14350
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12728 11937 12756 13670
rect 12820 13394 12848 14214
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12912 13258 12940 14962
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12714 11928 12770 11937
rect 12714 11863 12770 11872
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 12728 11354 12756 11562
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12636 11206 12756 11234
rect 12346 11183 12402 11192
rect 12256 11154 12308 11160
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12360 10470 12388 11086
rect 12438 10704 12494 10713
rect 12636 10674 12664 11086
rect 12438 10639 12494 10648
rect 12624 10668 12676 10674
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12034 9166 12112 9194
rect 12162 9208 12218 9217
rect 11978 9143 12034 9152
rect 12162 9143 12218 9152
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11886 8800 11942 8809
rect 11886 8735 11942 8744
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 11992 8022 12020 8502
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11900 5846 11928 7890
rect 11978 7848 12034 7857
rect 11978 7783 12034 7792
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11900 5370 11928 5646
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11796 5092 11848 5098
rect 11796 5034 11848 5040
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11440 4236 11560 4264
rect 11612 4276 11664 4282
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11244 3664 11296 3670
rect 11150 3632 11206 3641
rect 11060 3596 11112 3602
rect 10980 3556 11060 3584
rect 10980 3194 11008 3556
rect 11440 3652 11468 4236
rect 11612 4218 11664 4224
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11296 3624 11468 3652
rect 11244 3606 11296 3612
rect 11150 3567 11206 3576
rect 11060 3538 11112 3544
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10692 3052 10744 3058
rect 11256 3040 11284 3606
rect 11532 3534 11560 4082
rect 11716 4078 11744 4966
rect 11886 4856 11942 4865
rect 11886 4791 11942 4800
rect 11900 4758 11928 4791
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11808 4146 11836 4694
rect 11886 4584 11942 4593
rect 11886 4519 11942 4528
rect 11900 4486 11928 4519
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11702 3904 11758 3913
rect 11624 3738 11652 3878
rect 11702 3839 11758 3848
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11426 3360 11482 3369
rect 11426 3295 11482 3304
rect 10692 2994 10744 3000
rect 11164 3012 11284 3040
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 10612 2689 10640 2858
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10598 2680 10654 2689
rect 10817 2672 11113 2692
rect 10598 2615 10654 2624
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10324 1896 10376 1902
rect 10324 1838 10376 1844
rect 10336 1748 10364 1838
rect 10336 1720 10456 1748
rect 10428 480 10456 1720
rect 10612 882 10640 2615
rect 11164 1834 11192 3012
rect 11440 2854 11468 3295
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11334 2680 11390 2689
rect 11624 2632 11652 2790
rect 11390 2624 11652 2632
rect 11334 2615 11652 2624
rect 11348 2604 11652 2615
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11242 2136 11298 2145
rect 11242 2071 11298 2080
rect 11152 1828 11204 1834
rect 11152 1770 11204 1776
rect 11164 1494 11192 1770
rect 11152 1488 11204 1494
rect 11152 1430 11204 1436
rect 10782 1320 10838 1329
rect 10782 1255 10838 1264
rect 10600 876 10652 882
rect 10600 818 10652 824
rect 10796 480 10824 1255
rect 11256 480 11284 2071
rect 11348 1970 11376 2450
rect 11336 1964 11388 1970
rect 11336 1906 11388 1912
rect 11624 480 11652 2604
rect 11716 2582 11744 3839
rect 11886 3768 11942 3777
rect 11886 3703 11888 3712
rect 11940 3703 11942 3712
rect 11888 3674 11940 3680
rect 11992 3482 12020 7783
rect 12084 7528 12112 8978
rect 12176 8265 12204 9143
rect 12268 9042 12296 10406
rect 12452 9738 12480 10639
rect 12624 10610 12676 10616
rect 12636 10198 12664 10610
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12360 9710 12480 9738
rect 12360 9042 12388 9710
rect 12438 9208 12494 9217
rect 12438 9143 12494 9152
rect 12452 9110 12480 9143
rect 12440 9104 12492 9110
rect 12544 9081 12572 9998
rect 12636 9586 12664 9998
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12440 9046 12492 9052
rect 12530 9072 12586 9081
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12348 9036 12400 9042
rect 12530 9007 12586 9016
rect 12348 8978 12400 8984
rect 12360 8922 12388 8978
rect 12360 8894 12572 8922
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8634 12480 8774
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12162 8256 12218 8265
rect 12218 8214 12296 8242
rect 12162 8191 12218 8200
rect 12084 7500 12204 7528
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 5098 12112 7346
rect 12176 7177 12204 7500
rect 12268 7206 12296 8214
rect 12348 8084 12400 8090
rect 12544 8072 12572 8894
rect 12348 8026 12400 8032
rect 12452 8044 12572 8072
rect 12360 7857 12388 8026
rect 12346 7848 12402 7857
rect 12346 7783 12402 7792
rect 12452 7410 12480 8044
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12256 7200 12308 7206
rect 12162 7168 12218 7177
rect 12256 7142 12308 7148
rect 12162 7103 12218 7112
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 12072 5092 12124 5098
rect 12072 5034 12124 5040
rect 11900 3454 12020 3482
rect 11794 3224 11850 3233
rect 11794 3159 11850 3168
rect 11808 2938 11836 3159
rect 11900 3058 11928 3454
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 11808 2910 11928 2938
rect 11794 2816 11850 2825
rect 11794 2751 11850 2760
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 11704 2440 11756 2446
rect 11808 2417 11836 2751
rect 11900 2514 11928 2910
rect 11992 2689 12020 3334
rect 11978 2680 12034 2689
rect 11978 2615 12034 2624
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 11704 2382 11756 2388
rect 11794 2408 11850 2417
rect 11716 1562 11744 2382
rect 11794 2343 11850 2352
rect 11704 1556 11756 1562
rect 11704 1498 11756 1504
rect 12084 480 12112 5034
rect 12176 3670 12204 6734
rect 12268 6662 12296 6802
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12452 6458 12480 6870
rect 12544 6662 12572 7890
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12636 7002 12664 7346
rect 12728 7342 12756 11206
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12820 10985 12848 11154
rect 12806 10976 12862 10985
rect 12806 10911 12862 10920
rect 12808 10192 12860 10198
rect 12808 10134 12860 10140
rect 12820 9654 12848 10134
rect 12912 10130 12940 11494
rect 13004 10810 13032 14894
rect 13096 14770 13124 14962
rect 13096 14742 13216 14770
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13096 13530 13124 14554
rect 13188 13938 13216 14742
rect 13556 14550 13584 15030
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13280 14385 13308 14418
rect 13266 14376 13322 14385
rect 13266 14311 13322 14320
rect 13282 14172 13578 14192
rect 13338 14170 13362 14172
rect 13418 14170 13442 14172
rect 13498 14170 13522 14172
rect 13360 14118 13362 14170
rect 13424 14118 13436 14170
rect 13498 14118 13500 14170
rect 13338 14116 13362 14118
rect 13418 14116 13442 14118
rect 13498 14116 13522 14118
rect 13282 14096 13578 14116
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 13188 13240 13216 13874
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13096 13212 13216 13240
rect 13096 12102 13124 13212
rect 13280 13172 13308 13398
rect 13188 13144 13308 13172
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13082 11928 13138 11937
rect 13082 11863 13138 11872
rect 13096 11098 13124 11863
rect 13188 11694 13216 13144
rect 13282 13084 13578 13104
rect 13338 13082 13362 13084
rect 13418 13082 13442 13084
rect 13498 13082 13522 13084
rect 13360 13030 13362 13082
rect 13424 13030 13436 13082
rect 13498 13030 13500 13082
rect 13338 13028 13362 13030
rect 13418 13028 13442 13030
rect 13498 13028 13522 13030
rect 13282 13008 13578 13028
rect 13648 12714 13676 15302
rect 13740 13569 13768 15438
rect 13726 13560 13782 13569
rect 13726 13495 13782 13504
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13740 13297 13768 13398
rect 13726 13288 13782 13297
rect 13726 13223 13782 13232
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13450 12336 13506 12345
rect 13268 12300 13320 12306
rect 13450 12271 13506 12280
rect 13268 12242 13320 12248
rect 13280 12209 13308 12242
rect 13464 12238 13492 12271
rect 13452 12232 13504 12238
rect 13266 12200 13322 12209
rect 13544 12232 13596 12238
rect 13452 12174 13504 12180
rect 13542 12200 13544 12209
rect 13596 12200 13598 12209
rect 13266 12135 13322 12144
rect 13542 12135 13598 12144
rect 13282 11996 13578 12016
rect 13338 11994 13362 11996
rect 13418 11994 13442 11996
rect 13498 11994 13522 11996
rect 13360 11942 13362 11994
rect 13424 11942 13436 11994
rect 13498 11942 13500 11994
rect 13338 11940 13362 11942
rect 13418 11940 13442 11942
rect 13498 11940 13522 11942
rect 13282 11920 13578 11940
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13188 11529 13216 11630
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13174 11520 13230 11529
rect 13174 11455 13230 11464
rect 13280 11218 13308 11562
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13266 11112 13322 11121
rect 13096 11070 13216 11098
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12820 8537 12848 8978
rect 12806 8528 12862 8537
rect 12806 8463 12862 8472
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12636 6866 12664 6938
rect 12820 6934 12848 8230
rect 12912 7342 12940 9862
rect 13004 9217 13032 10474
rect 13096 10305 13124 10950
rect 13188 10441 13216 11070
rect 13266 11047 13268 11056
rect 13320 11047 13322 11056
rect 13268 11018 13320 11024
rect 13556 10996 13584 11494
rect 13648 11354 13676 12650
rect 13832 11830 13860 17520
rect 14200 15042 14228 17520
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14476 15706 14504 15846
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14200 15014 14320 15042
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 14016 13802 14044 14894
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14004 13796 14056 13802
rect 14004 13738 14056 13744
rect 14016 13410 14044 13738
rect 14108 13530 14136 14350
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14186 13424 14242 13433
rect 13924 13382 14136 13410
rect 13924 12782 13952 13382
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13820 11824 13872 11830
rect 13740 11784 13820 11812
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13634 11248 13690 11257
rect 13634 11183 13636 11192
rect 13688 11183 13690 11192
rect 13636 11154 13688 11160
rect 13556 10968 13676 10996
rect 13282 10908 13578 10928
rect 13338 10906 13362 10908
rect 13418 10906 13442 10908
rect 13498 10906 13522 10908
rect 13360 10854 13362 10906
rect 13424 10854 13436 10906
rect 13498 10854 13500 10906
rect 13338 10852 13362 10854
rect 13418 10852 13442 10854
rect 13498 10852 13522 10854
rect 13282 10832 13578 10852
rect 13648 10792 13676 10968
rect 13556 10764 13676 10792
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13174 10432 13230 10441
rect 13174 10367 13230 10376
rect 13082 10296 13138 10305
rect 13082 10231 13138 10240
rect 13188 10198 13216 10367
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13280 10044 13308 10542
rect 13556 10130 13584 10764
rect 13740 10690 13768 11784
rect 13820 11766 13872 11772
rect 13924 11218 13952 12582
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13912 11076 13964 11082
rect 13648 10662 13768 10690
rect 13832 11036 13912 11064
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13188 10016 13308 10044
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 13096 9586 13124 9930
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12990 9208 13046 9217
rect 12990 9143 13046 9152
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 13004 7546 13032 8910
rect 13096 8906 13124 9522
rect 13188 9364 13216 10016
rect 13282 9820 13578 9840
rect 13338 9818 13362 9820
rect 13418 9818 13442 9820
rect 13498 9818 13522 9820
rect 13360 9766 13362 9818
rect 13424 9766 13436 9818
rect 13498 9766 13500 9818
rect 13338 9764 13362 9766
rect 13418 9764 13442 9766
rect 13498 9764 13522 9766
rect 13282 9744 13578 9764
rect 13648 9654 13676 10662
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13740 10169 13768 10542
rect 13726 10160 13782 10169
rect 13726 10095 13782 10104
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13268 9376 13320 9382
rect 13188 9336 13268 9364
rect 13268 9318 13320 9324
rect 13280 8906 13308 9318
rect 13372 9110 13400 9522
rect 13634 9480 13690 9489
rect 13634 9415 13690 9424
rect 13648 9382 13676 9415
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13740 9178 13768 9998
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13360 9104 13412 9110
rect 13360 9046 13412 9052
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13082 8664 13138 8673
rect 13082 8599 13138 8608
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12808 6928 12860 6934
rect 12808 6870 12860 6876
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12268 6186 12296 6394
rect 12544 6322 12572 6598
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12912 6202 12940 7278
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13004 6322 13032 6734
rect 13096 6440 13124 8599
rect 13188 8090 13216 8774
rect 13282 8732 13578 8752
rect 13338 8730 13362 8732
rect 13418 8730 13442 8732
rect 13498 8730 13522 8732
rect 13360 8678 13362 8730
rect 13424 8678 13436 8730
rect 13498 8678 13500 8730
rect 13338 8676 13362 8678
rect 13418 8676 13442 8678
rect 13498 8676 13522 8678
rect 13282 8656 13578 8676
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13464 8294 13492 8434
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13188 7546 13216 7822
rect 13282 7644 13578 7664
rect 13338 7642 13362 7644
rect 13418 7642 13442 7644
rect 13498 7642 13522 7644
rect 13360 7590 13362 7642
rect 13424 7590 13436 7642
rect 13498 7590 13500 7642
rect 13338 7588 13362 7590
rect 13418 7588 13442 7590
rect 13498 7588 13522 7590
rect 13282 7568 13578 7588
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13268 7472 13320 7478
rect 13266 7440 13268 7449
rect 13320 7440 13322 7449
rect 13266 7375 13322 7384
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13266 7304 13322 7313
rect 13188 7177 13216 7278
rect 13266 7239 13322 7248
rect 13280 7206 13308 7239
rect 13268 7200 13320 7206
rect 13174 7168 13230 7177
rect 13268 7142 13320 7148
rect 13174 7103 13230 7112
rect 13188 6798 13216 7103
rect 13372 7041 13400 7346
rect 13358 7032 13414 7041
rect 13358 6967 13414 6976
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13176 6452 13228 6458
rect 13096 6412 13176 6440
rect 13176 6394 13228 6400
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12256 6180 12308 6186
rect 12912 6174 13032 6202
rect 12256 6122 12308 6128
rect 12440 6112 12492 6118
rect 12438 6080 12440 6089
rect 12532 6112 12584 6118
rect 12492 6080 12494 6089
rect 12532 6054 12584 6060
rect 12806 6080 12862 6089
rect 12438 6015 12494 6024
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12346 5672 12402 5681
rect 12256 5636 12308 5642
rect 12346 5607 12402 5616
rect 12256 5578 12308 5584
rect 12268 5409 12296 5578
rect 12254 5400 12310 5409
rect 12254 5335 12310 5344
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12164 3664 12216 3670
rect 12164 3606 12216 3612
rect 12268 1970 12296 4762
rect 12360 4554 12388 5607
rect 12452 4826 12480 5782
rect 12544 5030 12572 6054
rect 12806 6015 12862 6024
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12530 4856 12586 4865
rect 12440 4820 12492 4826
rect 12530 4791 12586 4800
rect 12440 4762 12492 4768
rect 12544 4622 12572 4791
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12440 4208 12492 4214
rect 12438 4176 12440 4185
rect 12492 4176 12494 4185
rect 12438 4111 12494 4120
rect 12544 4049 12572 4558
rect 12530 4040 12586 4049
rect 12530 3975 12586 3984
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 12346 3496 12402 3505
rect 12346 3431 12402 3440
rect 12256 1964 12308 1970
rect 12256 1906 12308 1912
rect 12360 1902 12388 3431
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12452 2310 12480 3334
rect 12544 3194 12572 3606
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12636 2990 12664 5714
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12728 5545 12756 5646
rect 12714 5536 12770 5545
rect 12714 5471 12770 5480
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12728 3534 12756 4490
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12714 3224 12770 3233
rect 12714 3159 12770 3168
rect 12728 2990 12756 3159
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12820 2582 12848 6015
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12912 3738 12940 4966
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 13004 3618 13032 6174
rect 13648 5914 13676 7822
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12912 3590 13032 3618
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 12728 2310 12756 2450
rect 12912 2378 12940 3590
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 2446 13032 3470
rect 13096 3466 13124 4762
rect 13282 4380 13578 4400
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 13648 4282 13676 5714
rect 13740 5710 13768 8434
rect 13832 8401 13860 11036
rect 13912 11018 13964 11024
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13924 9761 13952 10474
rect 13910 9752 13966 9761
rect 13910 9687 13966 9696
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13818 8392 13874 8401
rect 13818 8327 13874 8336
rect 13818 7984 13874 7993
rect 13818 7919 13874 7928
rect 13832 6730 13860 7919
rect 13924 7834 13952 9454
rect 14016 8129 14044 13126
rect 14108 9382 14136 13382
rect 14186 13359 14242 13368
rect 14200 12850 14228 13359
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14186 12744 14242 12753
rect 14186 12679 14242 12688
rect 14200 12306 14228 12679
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 14292 11286 14320 15014
rect 14554 14920 14610 14929
rect 14554 14855 14610 14864
rect 14568 14822 14596 14855
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 13841 14412 14214
rect 14370 13832 14426 13841
rect 14370 13767 14426 13776
rect 14660 12374 14688 17520
rect 15028 14600 15056 17520
rect 15488 15162 15516 17520
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15108 14884 15160 14890
rect 15108 14826 15160 14832
rect 14844 14572 15056 14600
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14660 11778 14688 12310
rect 14384 11750 14688 11778
rect 14280 11280 14332 11286
rect 14280 11222 14332 11228
rect 14292 10130 14320 11222
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14096 9376 14148 9382
rect 14292 9353 14320 9590
rect 14096 9318 14148 9324
rect 14278 9344 14334 9353
rect 14002 8120 14058 8129
rect 14002 8055 14058 8064
rect 14108 7993 14136 9318
rect 14278 9279 14334 9288
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14200 8809 14228 8978
rect 14186 8800 14242 8809
rect 14186 8735 14242 8744
rect 14292 8650 14320 9279
rect 14200 8622 14320 8650
rect 14094 7984 14150 7993
rect 14094 7919 14150 7928
rect 13924 7806 14136 7834
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13740 5302 13768 5646
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 13832 5148 13860 5782
rect 13740 5120 13860 5148
rect 13740 4826 13768 5120
rect 13818 4992 13874 5001
rect 13818 4927 13874 4936
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13648 4146 13676 4218
rect 13832 4214 13860 4927
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 13280 3738 13308 3946
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13084 3460 13136 3466
rect 13084 3402 13136 3408
rect 13082 3360 13138 3369
rect 13082 3295 13138 3304
rect 13096 3194 13124 3295
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 13096 2689 13124 2994
rect 13082 2680 13138 2689
rect 13082 2615 13138 2624
rect 13084 2508 13136 2514
rect 13084 2450 13136 2456
rect 12992 2440 13044 2446
rect 13096 2417 13124 2450
rect 12992 2382 13044 2388
rect 13082 2408 13138 2417
rect 12900 2372 12952 2378
rect 13082 2343 13138 2352
rect 12900 2314 12952 2320
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 12636 2038 12664 2246
rect 12624 2032 12676 2038
rect 12624 1974 12676 1980
rect 12348 1896 12400 1902
rect 12348 1838 12400 1844
rect 12530 1592 12586 1601
rect 12530 1527 12586 1536
rect 12544 480 12572 1527
rect 12912 480 12940 2314
rect 13082 2272 13138 2281
rect 13188 2258 13216 3470
rect 13280 3466 13308 3674
rect 13360 3664 13412 3670
rect 13452 3664 13504 3670
rect 13360 3606 13412 3612
rect 13450 3632 13452 3641
rect 13504 3632 13506 3641
rect 13372 3505 13400 3606
rect 13450 3567 13506 3576
rect 13358 3496 13414 3505
rect 13268 3460 13320 3466
rect 13358 3431 13414 3440
rect 13268 3402 13320 3408
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13372 2514 13400 2926
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13556 2378 13584 2926
rect 13648 2650 13676 3878
rect 13832 3777 13860 3878
rect 13818 3768 13874 3777
rect 13728 3732 13780 3738
rect 13818 3703 13874 3712
rect 13728 3674 13780 3680
rect 13740 3097 13768 3674
rect 13818 3496 13874 3505
rect 13818 3431 13874 3440
rect 13726 3088 13782 3097
rect 13726 3023 13782 3032
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 13138 2230 13216 2258
rect 13082 2207 13138 2216
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 13358 2000 13414 2009
rect 13358 1935 13414 1944
rect 13372 480 13400 1935
rect 13832 480 13860 3431
rect 13924 2922 13952 7686
rect 14016 6202 14044 7686
rect 14108 7274 14136 7806
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 14016 6174 14136 6202
rect 14108 5522 14136 6174
rect 14200 6118 14228 8622
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14292 8090 14320 8502
rect 14384 8430 14412 11750
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14476 8634 14504 11630
rect 14752 10826 14780 13466
rect 14844 13394 14872 14572
rect 14922 14512 14978 14521
rect 14922 14447 14978 14456
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14568 10798 14780 10826
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14384 7750 14412 8366
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 14476 7410 14504 8230
rect 14568 7410 14596 10798
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14752 10577 14780 10610
rect 14738 10568 14794 10577
rect 14738 10503 14794 10512
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 14646 10024 14702 10033
rect 14646 9959 14648 9968
rect 14700 9959 14702 9968
rect 14648 9930 14700 9936
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14660 9518 14688 9658
rect 14648 9512 14700 9518
rect 14752 9500 14780 10066
rect 14844 9654 14872 12718
rect 14832 9648 14884 9654
rect 14832 9590 14884 9596
rect 14752 9472 14872 9500
rect 14648 9454 14700 9460
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14648 8288 14700 8294
rect 14752 8265 14780 8366
rect 14648 8230 14700 8236
rect 14738 8256 14794 8265
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14292 5914 14320 6802
rect 14372 6792 14424 6798
rect 14476 6769 14504 7346
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 14372 6734 14424 6740
rect 14462 6760 14518 6769
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14016 5494 14136 5522
rect 14016 4690 14044 5494
rect 14094 5264 14150 5273
rect 14094 5199 14096 5208
rect 14148 5199 14150 5208
rect 14096 5170 14148 5176
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14016 4078 14044 4422
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 14108 3602 14136 5034
rect 14200 4593 14228 5714
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14186 4584 14242 4593
rect 14186 4519 14242 4528
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14016 3126 14044 3470
rect 14108 3194 14136 3538
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 14108 2650 14136 2994
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14200 2582 14228 4218
rect 14292 2650 14320 4966
rect 14384 3194 14412 6734
rect 14462 6695 14518 6704
rect 14476 5710 14504 6695
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14476 4282 14504 5306
rect 14568 4690 14596 7210
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14660 4570 14688 8230
rect 14738 8191 14794 8200
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14568 4542 14688 4570
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14462 4040 14518 4049
rect 14462 3975 14518 3984
rect 14476 3602 14504 3975
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14476 2854 14504 3402
rect 14464 2848 14516 2854
rect 14568 2825 14596 4542
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14660 4185 14688 4422
rect 14646 4176 14702 4185
rect 14646 4111 14702 4120
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14464 2790 14516 2796
rect 14554 2816 14610 2825
rect 14554 2751 14610 2760
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 14188 1964 14240 1970
rect 14188 1906 14240 1912
rect 14200 480 14228 1906
rect 14660 480 14688 4014
rect 14752 626 14780 7482
rect 14844 7426 14872 9472
rect 14936 7546 14964 14447
rect 15016 14000 15068 14006
rect 15014 13968 15016 13977
rect 15068 13968 15070 13977
rect 15014 13903 15070 13912
rect 15120 12782 15148 14826
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15488 11218 15516 15098
rect 15948 11694 15976 17520
rect 16316 14890 16344 17520
rect 16304 14884 16356 14890
rect 16304 14826 16356 14832
rect 16776 14482 16804 17520
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15016 9648 15068 9654
rect 15014 9616 15016 9625
rect 15068 9616 15070 9625
rect 15014 9551 15070 9560
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14844 7398 14964 7426
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14844 3058 14872 5646
rect 14936 5642 14964 7398
rect 15016 6384 15068 6390
rect 15014 6352 15016 6361
rect 15068 6352 15070 6361
rect 15014 6287 15070 6296
rect 14924 5636 14976 5642
rect 14924 5578 14976 5584
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 15028 4554 15056 4966
rect 15016 4548 15068 4554
rect 15016 4490 15068 4496
rect 14922 4176 14978 4185
rect 14922 4111 14978 4120
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14936 2446 14964 4111
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 15028 2961 15056 3878
rect 15014 2952 15070 2961
rect 15014 2887 15070 2896
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 15028 2106 15056 2246
rect 15016 2100 15068 2106
rect 15016 2042 15068 2048
rect 15120 1766 15148 8910
rect 15212 6186 15240 10406
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 15304 6934 15332 8842
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15292 6928 15344 6934
rect 15292 6870 15344 6876
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 15212 5914 15240 6122
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15396 4185 15424 7822
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15382 4176 15438 4185
rect 15382 4111 15438 4120
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15304 2990 15332 3334
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 15476 1828 15528 1834
rect 15476 1770 15528 1776
rect 15108 1760 15160 1766
rect 15108 1702 15160 1708
rect 14752 598 15056 626
rect 15028 480 15056 598
rect 15488 480 15516 1770
rect 15948 480 15976 7142
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16762 6896 16818 6905
rect 16316 480 16344 6870
rect 16762 6831 16818 6840
rect 16776 480 16804 6831
rect 2778 439 2834 448
rect 3146 0 3202 480
rect 3606 0 3662 480
rect 3974 0 4030 480
rect 4434 0 4490 480
rect 4802 0 4858 480
rect 5262 0 5318 480
rect 5722 0 5778 480
rect 6090 0 6146 480
rect 6550 0 6606 480
rect 7010 0 7066 480
rect 7378 0 7434 480
rect 7838 0 7894 480
rect 8206 0 8262 480
rect 8666 0 8722 480
rect 9126 0 9182 480
rect 9494 0 9550 480
rect 9954 0 10010 480
rect 10414 0 10470 480
rect 10782 0 10838 480
rect 11242 0 11298 480
rect 11610 0 11666 480
rect 12070 0 12126 480
rect 12530 0 12586 480
rect 12898 0 12954 480
rect 13358 0 13414 480
rect 13818 0 13874 480
rect 14186 0 14242 480
rect 14646 0 14702 480
rect 15014 0 15070 480
rect 15474 0 15530 480
rect 15934 0 15990 480
rect 16302 0 16358 480
rect 16762 0 16818 480
<< via2 >>
rect 1030 14864 1086 14920
rect 1490 14320 1546 14376
rect 1674 9832 1730 9888
rect 1582 9016 1638 9072
rect 1398 6860 1454 6896
rect 1398 6840 1400 6860
rect 1400 6840 1452 6860
rect 1452 6840 1454 6860
rect 570 3440 626 3496
rect 1030 2896 1086 2952
rect 1950 17312 2006 17368
rect 1858 13368 1914 13424
rect 1950 12416 2006 12472
rect 1858 9832 1914 9888
rect 2042 11228 2044 11248
rect 2044 11228 2096 11248
rect 2096 11228 2098 11248
rect 2042 11192 2098 11228
rect 1950 9444 2006 9480
rect 1950 9424 1952 9444
rect 1952 9424 2004 9444
rect 2004 9424 2006 9444
rect 1858 6432 1914 6488
rect 1858 5208 1914 5264
rect 2042 7948 2098 7984
rect 2042 7928 2044 7948
rect 2044 7928 2096 7948
rect 2096 7928 2098 7948
rect 2410 13776 2466 13832
rect 2226 12280 2282 12336
rect 2410 8916 2412 8936
rect 2412 8916 2464 8936
rect 2464 8916 2466 8936
rect 2410 8880 2466 8916
rect 2318 8472 2374 8528
rect 2502 7792 2558 7848
rect 2042 3712 2098 3768
rect 2870 12144 2926 12200
rect 3054 14048 3110 14104
rect 4066 16244 4122 16280
rect 4066 16224 4068 16244
rect 4068 16224 4120 16244
rect 4120 16224 4122 16244
rect 4066 15408 4122 15464
rect 3421 15258 3477 15260
rect 3501 15258 3557 15260
rect 3581 15258 3637 15260
rect 3661 15258 3717 15260
rect 3421 15206 3447 15258
rect 3447 15206 3477 15258
rect 3501 15206 3511 15258
rect 3511 15206 3557 15258
rect 3581 15206 3627 15258
rect 3627 15206 3637 15258
rect 3661 15206 3691 15258
rect 3691 15206 3717 15258
rect 3421 15204 3477 15206
rect 3501 15204 3557 15206
rect 3581 15204 3637 15206
rect 3661 15204 3717 15206
rect 4066 15020 4122 15056
rect 4066 15000 4068 15020
rect 4068 15000 4120 15020
rect 4120 15000 4122 15020
rect 4250 14592 4306 14648
rect 3421 14170 3477 14172
rect 3501 14170 3557 14172
rect 3581 14170 3637 14172
rect 3661 14170 3717 14172
rect 3421 14118 3447 14170
rect 3447 14118 3477 14170
rect 3501 14118 3511 14170
rect 3511 14118 3557 14170
rect 3581 14118 3627 14170
rect 3627 14118 3637 14170
rect 3661 14118 3691 14170
rect 3691 14118 3717 14170
rect 3421 14116 3477 14118
rect 3501 14116 3557 14118
rect 3581 14116 3637 14118
rect 3661 14116 3717 14118
rect 3054 13232 3110 13288
rect 2778 11600 2834 11656
rect 2686 11464 2742 11520
rect 2686 11348 2742 11384
rect 2686 11328 2688 11348
rect 2688 11328 2740 11348
rect 2740 11328 2742 11348
rect 3421 13082 3477 13084
rect 3501 13082 3557 13084
rect 3581 13082 3637 13084
rect 3661 13082 3717 13084
rect 3421 13030 3447 13082
rect 3447 13030 3477 13082
rect 3501 13030 3511 13082
rect 3511 13030 3557 13082
rect 3581 13030 3627 13082
rect 3627 13030 3637 13082
rect 3661 13030 3691 13082
rect 3691 13030 3717 13082
rect 3421 13028 3477 13030
rect 3501 13028 3557 13030
rect 3581 13028 3637 13030
rect 3661 13028 3717 13030
rect 3606 12552 3662 12608
rect 3421 11994 3477 11996
rect 3501 11994 3557 11996
rect 3581 11994 3637 11996
rect 3661 11994 3717 11996
rect 3421 11942 3447 11994
rect 3447 11942 3477 11994
rect 3501 11942 3511 11994
rect 3511 11942 3557 11994
rect 3581 11942 3627 11994
rect 3627 11942 3637 11994
rect 3661 11942 3691 11994
rect 3691 11942 3717 11994
rect 3421 11940 3477 11942
rect 3501 11940 3557 11942
rect 3581 11940 3637 11942
rect 3661 11940 3717 11942
rect 3974 14456 4030 14512
rect 3974 14048 4030 14104
rect 4158 13912 4214 13968
rect 4158 12960 4214 13016
rect 4066 12416 4122 12472
rect 4066 12144 4122 12200
rect 2870 11056 2926 11112
rect 2870 10512 2926 10568
rect 3422 11464 3478 11520
rect 2778 9560 2834 9616
rect 2870 8744 2926 8800
rect 2778 7384 2834 7440
rect 2594 5752 2650 5808
rect 2778 5752 2834 5808
rect 2962 8236 2964 8256
rect 2964 8236 3016 8256
rect 3016 8236 3018 8256
rect 2962 8200 3018 8236
rect 2686 4800 2742 4856
rect 2870 3848 2926 3904
rect 2778 2760 2834 2816
rect 2778 2644 2834 2680
rect 2778 2624 2780 2644
rect 2780 2624 2832 2644
rect 2832 2624 2834 2644
rect 3421 10906 3477 10908
rect 3501 10906 3557 10908
rect 3581 10906 3637 10908
rect 3661 10906 3717 10908
rect 3421 10854 3447 10906
rect 3447 10854 3477 10906
rect 3501 10854 3511 10906
rect 3511 10854 3557 10906
rect 3581 10854 3627 10906
rect 3627 10854 3637 10906
rect 3661 10854 3691 10906
rect 3691 10854 3717 10906
rect 3421 10852 3477 10854
rect 3501 10852 3557 10854
rect 3581 10852 3637 10854
rect 3661 10852 3717 10854
rect 3330 10648 3386 10704
rect 3606 10648 3662 10704
rect 3421 9818 3477 9820
rect 3501 9818 3557 9820
rect 3581 9818 3637 9820
rect 3661 9818 3717 9820
rect 3421 9766 3447 9818
rect 3447 9766 3477 9818
rect 3501 9766 3511 9818
rect 3511 9766 3557 9818
rect 3581 9766 3627 9818
rect 3627 9766 3637 9818
rect 3661 9766 3691 9818
rect 3691 9766 3717 9818
rect 3421 9764 3477 9766
rect 3501 9764 3557 9766
rect 3581 9764 3637 9766
rect 3661 9764 3717 9766
rect 3606 9152 3662 9208
rect 3421 8730 3477 8732
rect 3501 8730 3557 8732
rect 3581 8730 3637 8732
rect 3661 8730 3717 8732
rect 3421 8678 3447 8730
rect 3447 8678 3477 8730
rect 3501 8678 3511 8730
rect 3511 8678 3557 8730
rect 3581 8678 3627 8730
rect 3627 8678 3637 8730
rect 3661 8678 3691 8730
rect 3691 8678 3717 8730
rect 3421 8676 3477 8678
rect 3501 8676 3557 8678
rect 3581 8676 3637 8678
rect 3661 8676 3717 8678
rect 3330 8336 3386 8392
rect 3421 7642 3477 7644
rect 3501 7642 3557 7644
rect 3581 7642 3637 7644
rect 3661 7642 3717 7644
rect 3421 7590 3447 7642
rect 3447 7590 3477 7642
rect 3501 7590 3511 7642
rect 3511 7590 3557 7642
rect 3581 7590 3627 7642
rect 3627 7590 3637 7642
rect 3661 7590 3691 7642
rect 3691 7590 3717 7642
rect 3421 7588 3477 7590
rect 3501 7588 3557 7590
rect 3581 7588 3637 7590
rect 3661 7588 3717 7590
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 4066 10512 4122 10568
rect 3974 8064 4030 8120
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 3882 5616 3938 5672
rect 4066 7520 4122 7576
rect 4158 6840 4214 6896
rect 4158 6568 4214 6624
rect 4158 6432 4214 6488
rect 4066 6160 4122 6216
rect 4158 6024 4214 6080
rect 4434 13912 4490 13968
rect 4618 13932 4674 13968
rect 4618 13912 4620 13932
rect 4620 13912 4672 13932
rect 4672 13912 4674 13932
rect 4526 13640 4582 13696
rect 4342 12688 4398 12744
rect 4618 13504 4674 13560
rect 4710 12960 4766 13016
rect 4342 10104 4398 10160
rect 4894 12008 4950 12064
rect 5630 15136 5686 15192
rect 5886 15802 5942 15804
rect 5966 15802 6022 15804
rect 6046 15802 6102 15804
rect 6126 15802 6182 15804
rect 5886 15750 5912 15802
rect 5912 15750 5942 15802
rect 5966 15750 5976 15802
rect 5976 15750 6022 15802
rect 6046 15750 6092 15802
rect 6092 15750 6102 15802
rect 6126 15750 6156 15802
rect 6156 15750 6182 15802
rect 5886 15748 5942 15750
rect 5966 15748 6022 15750
rect 6046 15748 6102 15750
rect 6126 15748 6182 15750
rect 5446 14728 5502 14784
rect 6274 14728 6330 14784
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 6126 14714 6182 14716
rect 5886 14662 5912 14714
rect 5912 14662 5942 14714
rect 5966 14662 5976 14714
rect 5976 14662 6022 14714
rect 6046 14662 6092 14714
rect 6092 14662 6102 14714
rect 6126 14662 6156 14714
rect 6156 14662 6182 14714
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 6126 14660 6182 14662
rect 5078 11464 5134 11520
rect 4986 10920 5042 10976
rect 4802 10240 4858 10296
rect 4526 7248 4582 7304
rect 4342 7112 4398 7168
rect 4434 6996 4490 7032
rect 4434 6976 4436 6996
rect 4436 6976 4488 6996
rect 4488 6976 4490 6996
rect 4434 6740 4436 6760
rect 4436 6740 4488 6760
rect 4488 6740 4490 6760
rect 4434 6704 4490 6740
rect 4066 5480 4122 5536
rect 4066 5072 4122 5128
rect 2778 448 2834 504
rect 3882 4528 3938 4584
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 3882 4256 3938 4312
rect 3790 4004 3846 4040
rect 3790 3984 3792 4004
rect 3792 3984 3844 4004
rect 3844 3984 3846 4004
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 4066 2488 4122 2544
rect 4710 6296 4766 6352
rect 4710 5616 4766 5672
rect 4618 5344 4674 5400
rect 4526 4800 4582 4856
rect 5262 13232 5318 13288
rect 5906 14184 5962 14240
rect 5446 13504 5502 13560
rect 6366 13912 6422 13968
rect 5722 13640 5778 13696
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 6126 13626 6182 13628
rect 5886 13574 5912 13626
rect 5912 13574 5942 13626
rect 5966 13574 5976 13626
rect 5976 13574 6022 13626
rect 6046 13574 6092 13626
rect 6092 13574 6102 13626
rect 6126 13574 6156 13626
rect 6156 13574 6182 13626
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 6126 13572 6182 13574
rect 5354 12824 5410 12880
rect 5538 12824 5594 12880
rect 5354 12144 5410 12200
rect 6090 12844 6146 12880
rect 6090 12824 6092 12844
rect 6092 12824 6144 12844
rect 6144 12824 6146 12844
rect 5538 12416 5594 12472
rect 5354 12008 5410 12064
rect 5538 11056 5594 11112
rect 5170 9696 5226 9752
rect 5722 12552 5778 12608
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 6126 12538 6182 12540
rect 5886 12486 5912 12538
rect 5912 12486 5942 12538
rect 5966 12486 5976 12538
rect 5976 12486 6022 12538
rect 6046 12486 6092 12538
rect 6092 12486 6102 12538
rect 6126 12486 6156 12538
rect 6156 12486 6182 12538
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 6126 12484 6182 12486
rect 6366 12416 6422 12472
rect 6826 15272 6882 15328
rect 6734 14592 6790 14648
rect 6642 13912 6698 13968
rect 6550 12824 6606 12880
rect 7102 15136 7158 15192
rect 7470 15952 7526 16008
rect 7194 14592 7250 14648
rect 7010 13640 7066 13696
rect 6734 12552 6790 12608
rect 5722 11464 5778 11520
rect 5722 11328 5778 11384
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 6126 11450 6182 11452
rect 5886 11398 5912 11450
rect 5912 11398 5942 11450
rect 5966 11398 5976 11450
rect 5976 11398 6022 11450
rect 6046 11398 6092 11450
rect 6092 11398 6102 11450
rect 6126 11398 6156 11450
rect 6156 11398 6182 11450
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 6126 11396 6182 11398
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 6126 10362 6182 10364
rect 5886 10310 5912 10362
rect 5912 10310 5942 10362
rect 5966 10310 5976 10362
rect 5976 10310 6022 10362
rect 6046 10310 6092 10362
rect 6092 10310 6102 10362
rect 6126 10310 6156 10362
rect 6156 10310 6182 10362
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 6126 10308 6182 10310
rect 5078 9172 5134 9208
rect 5078 9152 5080 9172
rect 5080 9152 5132 9172
rect 5132 9152 5134 9172
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 6126 9274 6182 9276
rect 5886 9222 5912 9274
rect 5912 9222 5942 9274
rect 5966 9222 5976 9274
rect 5976 9222 6022 9274
rect 6046 9222 6092 9274
rect 6092 9222 6102 9274
rect 6126 9222 6156 9274
rect 6156 9222 6182 9274
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 6126 9220 6182 9222
rect 5538 8200 5594 8256
rect 6182 8744 6238 8800
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 6126 8186 6182 8188
rect 5886 8134 5912 8186
rect 5912 8134 5942 8186
rect 5966 8134 5976 8186
rect 5976 8134 6022 8186
rect 6046 8134 6092 8186
rect 6092 8134 6102 8186
rect 6126 8134 6156 8186
rect 6156 8134 6182 8186
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 6126 8132 6182 8134
rect 6274 8064 6330 8120
rect 4986 7656 5042 7712
rect 4986 6296 5042 6352
rect 4526 3576 4582 3632
rect 4434 3304 4490 3360
rect 4526 2896 4582 2952
rect 4250 1808 4306 1864
rect 4434 2760 4490 2816
rect 4802 3168 4858 3224
rect 4802 2896 4858 2952
rect 4434 1944 4490 2000
rect 5446 7812 5502 7848
rect 5446 7792 5448 7812
rect 5448 7792 5500 7812
rect 5500 7792 5502 7812
rect 5446 7112 5502 7168
rect 6274 7540 6330 7576
rect 6274 7520 6276 7540
rect 6276 7520 6328 7540
rect 6328 7520 6330 7540
rect 5722 6976 5778 7032
rect 5262 6432 5318 6488
rect 4986 4664 5042 4720
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 6126 7098 6182 7100
rect 5886 7046 5912 7098
rect 5912 7046 5942 7098
rect 5966 7046 5976 7098
rect 5976 7046 6022 7098
rect 6046 7046 6092 7098
rect 6092 7046 6102 7098
rect 6126 7046 6156 7098
rect 6156 7046 6182 7098
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 6126 7044 6182 7046
rect 5446 6024 5502 6080
rect 5354 5072 5410 5128
rect 5262 3168 5318 3224
rect 5170 3032 5226 3088
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 5814 5208 5870 5264
rect 5722 4800 5778 4856
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 5814 4664 5870 4720
rect 5630 3712 5686 3768
rect 5538 3168 5594 3224
rect 5814 4392 5870 4448
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 5630 2644 5686 2680
rect 5630 2624 5632 2644
rect 5632 2624 5684 2644
rect 5684 2624 5686 2644
rect 5262 2488 5318 2544
rect 4986 2352 5042 2408
rect 6458 11464 6514 11520
rect 6550 10512 6606 10568
rect 6458 10376 6514 10432
rect 6826 10784 6882 10840
rect 6826 10512 6882 10568
rect 7102 11464 7158 11520
rect 7102 10920 7158 10976
rect 7654 14728 7710 14784
rect 8206 15272 8262 15328
rect 8352 15258 8408 15260
rect 8432 15258 8488 15260
rect 8512 15258 8568 15260
rect 8592 15258 8648 15260
rect 8352 15206 8378 15258
rect 8378 15206 8408 15258
rect 8432 15206 8442 15258
rect 8442 15206 8488 15258
rect 8512 15206 8558 15258
rect 8558 15206 8568 15258
rect 8592 15206 8622 15258
rect 8622 15206 8648 15258
rect 8352 15204 8408 15206
rect 8432 15204 8488 15206
rect 8512 15204 8568 15206
rect 8592 15204 8648 15206
rect 8666 14456 8722 14512
rect 7838 14320 7894 14376
rect 7746 13676 7748 13696
rect 7748 13676 7800 13696
rect 7800 13676 7802 13696
rect 7746 13640 7802 13676
rect 7378 12280 7434 12336
rect 7562 12280 7618 12336
rect 7378 10376 7434 10432
rect 6734 8472 6790 8528
rect 6918 8472 6974 8528
rect 7102 8200 7158 8256
rect 6734 6296 6790 6352
rect 6642 4936 6698 4992
rect 6734 4120 6790 4176
rect 6550 3984 6606 4040
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 6550 2624 6606 2680
rect 5998 1536 6054 1592
rect 6734 2760 6790 2816
rect 7010 5092 7066 5128
rect 7010 5072 7012 5092
rect 7012 5072 7064 5092
rect 7064 5072 7066 5092
rect 7010 4800 7066 4856
rect 7010 4528 7066 4584
rect 7562 11464 7618 11520
rect 8352 14170 8408 14172
rect 8432 14170 8488 14172
rect 8512 14170 8568 14172
rect 8592 14170 8648 14172
rect 8352 14118 8378 14170
rect 8378 14118 8408 14170
rect 8432 14118 8442 14170
rect 8442 14118 8488 14170
rect 8512 14118 8558 14170
rect 8558 14118 8568 14170
rect 8592 14118 8622 14170
rect 8622 14118 8648 14170
rect 8352 14116 8408 14118
rect 8432 14116 8488 14118
rect 8512 14116 8568 14118
rect 8592 14116 8648 14118
rect 8206 14048 8262 14104
rect 8298 13368 8354 13424
rect 8942 15544 8998 15600
rect 8942 14592 8998 14648
rect 8850 14048 8906 14104
rect 8206 13096 8262 13152
rect 8022 12960 8078 13016
rect 7746 12824 7802 12880
rect 7654 9696 7710 9752
rect 7470 8608 7526 8664
rect 7470 7656 7526 7712
rect 7194 6432 7250 6488
rect 7286 6024 7342 6080
rect 7286 5344 7342 5400
rect 7378 4528 7434 4584
rect 7194 4392 7250 4448
rect 6918 3848 6974 3904
rect 7194 3732 7250 3768
rect 7194 3712 7196 3732
rect 7196 3712 7248 3732
rect 7248 3712 7250 3732
rect 6918 3304 6974 3360
rect 7102 3304 7158 3360
rect 7378 3304 7434 3360
rect 7010 2624 7066 2680
rect 8114 12824 8170 12880
rect 8758 13096 8814 13152
rect 8352 13082 8408 13084
rect 8432 13082 8488 13084
rect 8512 13082 8568 13084
rect 8592 13082 8648 13084
rect 8352 13030 8378 13082
rect 8378 13030 8408 13082
rect 8432 13030 8442 13082
rect 8442 13030 8488 13082
rect 8512 13030 8558 13082
rect 8558 13030 8568 13082
rect 8592 13030 8622 13082
rect 8622 13030 8648 13082
rect 8352 13028 8408 13030
rect 8432 13028 8488 13030
rect 8512 13028 8568 13030
rect 8592 13028 8648 13030
rect 9218 15408 9274 15464
rect 9310 15136 9366 15192
rect 9126 14728 9182 14784
rect 9034 13504 9090 13560
rect 8942 12960 8998 13016
rect 8114 11872 8170 11928
rect 8352 11994 8408 11996
rect 8432 11994 8488 11996
rect 8512 11994 8568 11996
rect 8592 11994 8648 11996
rect 8352 11942 8378 11994
rect 8378 11942 8408 11994
rect 8432 11942 8442 11994
rect 8442 11942 8488 11994
rect 8512 11942 8558 11994
rect 8558 11942 8568 11994
rect 8592 11942 8622 11994
rect 8622 11942 8648 11994
rect 8352 11940 8408 11942
rect 8432 11940 8488 11942
rect 8512 11940 8568 11942
rect 8592 11940 8648 11942
rect 8022 10920 8078 10976
rect 8114 10784 8170 10840
rect 7838 9696 7894 9752
rect 7930 8744 7986 8800
rect 8114 8608 8170 8664
rect 8022 8472 8078 8528
rect 8758 12008 8814 12064
rect 8352 10906 8408 10908
rect 8432 10906 8488 10908
rect 8512 10906 8568 10908
rect 8592 10906 8648 10908
rect 8352 10854 8378 10906
rect 8378 10854 8408 10906
rect 8432 10854 8442 10906
rect 8442 10854 8488 10906
rect 8512 10854 8558 10906
rect 8558 10854 8568 10906
rect 8592 10854 8622 10906
rect 8622 10854 8648 10906
rect 8352 10852 8408 10854
rect 8432 10852 8488 10854
rect 8512 10852 8568 10854
rect 8592 10852 8648 10854
rect 8850 10920 8906 10976
rect 8352 9818 8408 9820
rect 8432 9818 8488 9820
rect 8512 9818 8568 9820
rect 8592 9818 8648 9820
rect 8352 9766 8378 9818
rect 8378 9766 8408 9818
rect 8432 9766 8442 9818
rect 8442 9766 8488 9818
rect 8512 9766 8558 9818
rect 8558 9766 8568 9818
rect 8592 9766 8622 9818
rect 8622 9766 8648 9818
rect 8352 9764 8408 9766
rect 8432 9764 8488 9766
rect 8512 9764 8568 9766
rect 8592 9764 8648 9766
rect 8758 8916 8760 8936
rect 8760 8916 8812 8936
rect 8812 8916 8814 8936
rect 8758 8880 8814 8916
rect 8352 8730 8408 8732
rect 8432 8730 8488 8732
rect 8512 8730 8568 8732
rect 8592 8730 8648 8732
rect 8352 8678 8378 8730
rect 8378 8678 8408 8730
rect 8432 8678 8442 8730
rect 8442 8678 8488 8730
rect 8512 8678 8558 8730
rect 8558 8678 8568 8730
rect 8592 8678 8622 8730
rect 8622 8678 8648 8730
rect 8352 8676 8408 8678
rect 8432 8676 8488 8678
rect 8512 8676 8568 8678
rect 8592 8676 8648 8678
rect 8022 7656 8078 7712
rect 8206 7656 8262 7712
rect 8352 7642 8408 7644
rect 8432 7642 8488 7644
rect 8512 7642 8568 7644
rect 8592 7642 8648 7644
rect 8352 7590 8378 7642
rect 8378 7590 8408 7642
rect 8432 7590 8442 7642
rect 8442 7590 8488 7642
rect 8512 7590 8558 7642
rect 8558 7590 8568 7642
rect 8592 7590 8622 7642
rect 8622 7590 8648 7642
rect 8352 7588 8408 7590
rect 8432 7588 8488 7590
rect 8512 7588 8568 7590
rect 8592 7588 8648 7590
rect 7930 7112 7986 7168
rect 7838 6024 7894 6080
rect 8390 7112 8446 7168
rect 8666 7112 8722 7168
rect 8298 6704 8354 6760
rect 8482 6704 8538 6760
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 8206 6432 8262 6488
rect 8206 6060 8208 6080
rect 8208 6060 8260 6080
rect 8260 6060 8262 6080
rect 8206 6024 8262 6060
rect 7838 2760 7894 2816
rect 7562 2216 7618 2272
rect 7930 2352 7986 2408
rect 8574 6024 8630 6080
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 8114 5344 8170 5400
rect 8114 4428 8116 4448
rect 8116 4428 8168 4448
rect 8168 4428 8170 4448
rect 8114 4392 8170 4428
rect 8114 4256 8170 4312
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 9034 7656 9090 7712
rect 8942 7520 8998 7576
rect 9310 14048 9366 14104
rect 9310 13368 9366 13424
rect 9310 12416 9366 12472
rect 9310 10784 9366 10840
rect 9218 9152 9274 9208
rect 9218 8880 9274 8936
rect 9310 8200 9366 8256
rect 8942 6432 8998 6488
rect 8942 6024 8998 6080
rect 8942 4392 8998 4448
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 8206 3168 8262 3224
rect 8206 2624 8262 2680
rect 8574 2624 8630 2680
rect 8758 2488 8814 2544
rect 9034 4256 9090 4312
rect 9494 14592 9550 14648
rect 9678 14456 9734 14512
rect 9862 14184 9918 14240
rect 9862 13504 9918 13560
rect 9862 12960 9918 13016
rect 9770 10920 9826 10976
rect 9586 10784 9642 10840
rect 9678 10684 9680 10704
rect 9680 10684 9732 10704
rect 9732 10684 9734 10704
rect 9678 10648 9734 10684
rect 10414 14728 10470 14784
rect 10414 14592 10470 14648
rect 10506 13504 10562 13560
rect 10506 13388 10562 13424
rect 10506 13368 10508 13388
rect 10508 13368 10560 13388
rect 10560 13368 10562 13388
rect 10506 12552 10562 12608
rect 10817 15802 10873 15804
rect 10897 15802 10953 15804
rect 10977 15802 11033 15804
rect 11057 15802 11113 15804
rect 10817 15750 10843 15802
rect 10843 15750 10873 15802
rect 10897 15750 10907 15802
rect 10907 15750 10953 15802
rect 10977 15750 11023 15802
rect 11023 15750 11033 15802
rect 11057 15750 11087 15802
rect 11087 15750 11113 15802
rect 10817 15748 10873 15750
rect 10897 15748 10953 15750
rect 10977 15748 11033 15750
rect 11057 15748 11113 15750
rect 10817 14714 10873 14716
rect 10897 14714 10953 14716
rect 10977 14714 11033 14716
rect 11057 14714 11113 14716
rect 10817 14662 10843 14714
rect 10843 14662 10873 14714
rect 10897 14662 10907 14714
rect 10907 14662 10953 14714
rect 10977 14662 11023 14714
rect 11023 14662 11033 14714
rect 11057 14662 11087 14714
rect 11087 14662 11113 14714
rect 10817 14660 10873 14662
rect 10897 14660 10953 14662
rect 10977 14660 11033 14662
rect 11057 14660 11113 14662
rect 11518 15952 11574 16008
rect 11242 13676 11244 13696
rect 11244 13676 11296 13696
rect 11296 13676 11298 13696
rect 11242 13640 11298 13676
rect 10817 13626 10873 13628
rect 10897 13626 10953 13628
rect 10977 13626 11033 13628
rect 11057 13626 11113 13628
rect 10817 13574 10843 13626
rect 10843 13574 10873 13626
rect 10897 13574 10907 13626
rect 10907 13574 10953 13626
rect 10977 13574 11023 13626
rect 11023 13574 11033 13626
rect 11057 13574 11087 13626
rect 11087 13574 11113 13626
rect 10817 13572 10873 13574
rect 10897 13572 10953 13574
rect 10977 13572 11033 13574
rect 11057 13572 11113 13574
rect 11702 15136 11758 15192
rect 11794 14764 11796 14784
rect 11796 14764 11848 14784
rect 11848 14764 11850 14784
rect 11794 14728 11850 14764
rect 12070 14184 12126 14240
rect 11610 13504 11666 13560
rect 11242 12960 11298 13016
rect 10817 12538 10873 12540
rect 10897 12538 10953 12540
rect 10977 12538 11033 12540
rect 11057 12538 11113 12540
rect 10817 12486 10843 12538
rect 10843 12486 10873 12538
rect 10897 12486 10907 12538
rect 10907 12486 10953 12538
rect 10977 12486 11023 12538
rect 11023 12486 11033 12538
rect 11057 12486 11087 12538
rect 11087 12486 11113 12538
rect 10817 12484 10873 12486
rect 10897 12484 10953 12486
rect 10977 12484 11033 12486
rect 11057 12484 11113 12486
rect 10782 12144 10838 12200
rect 9770 9696 9826 9752
rect 9770 8200 9826 8256
rect 9402 6840 9458 6896
rect 9586 7112 9642 7168
rect 9586 6976 9642 7032
rect 9862 6976 9918 7032
rect 10414 10548 10416 10568
rect 10416 10548 10468 10568
rect 10468 10548 10470 10568
rect 10414 10512 10470 10548
rect 11334 12008 11390 12064
rect 10598 11464 10654 11520
rect 10817 11450 10873 11452
rect 10897 11450 10953 11452
rect 10977 11450 11033 11452
rect 11057 11450 11113 11452
rect 10817 11398 10843 11450
rect 10843 11398 10873 11450
rect 10897 11398 10907 11450
rect 10907 11398 10953 11450
rect 10977 11398 11023 11450
rect 11023 11398 11033 11450
rect 11057 11398 11087 11450
rect 11087 11398 11113 11450
rect 10817 11396 10873 11398
rect 10897 11396 10953 11398
rect 10977 11396 11033 11398
rect 11057 11396 11113 11398
rect 10690 11056 10746 11112
rect 10598 10920 10654 10976
rect 11242 11192 11298 11248
rect 11978 13252 12034 13288
rect 11978 13232 11980 13252
rect 11980 13232 12032 13252
rect 12032 13232 12034 13252
rect 12346 14456 12402 14512
rect 12346 14048 12402 14104
rect 12162 13640 12218 13696
rect 10598 10240 10654 10296
rect 10414 10104 10470 10160
rect 10598 10104 10654 10160
rect 10817 10362 10873 10364
rect 10897 10362 10953 10364
rect 10977 10362 11033 10364
rect 11057 10362 11113 10364
rect 10817 10310 10843 10362
rect 10843 10310 10873 10362
rect 10897 10310 10907 10362
rect 10907 10310 10953 10362
rect 10977 10310 11023 10362
rect 11023 10310 11033 10362
rect 11057 10310 11087 10362
rect 11087 10310 11113 10362
rect 10817 10308 10873 10310
rect 10897 10308 10953 10310
rect 10977 10308 11033 10310
rect 11057 10308 11113 10310
rect 10138 9696 10194 9752
rect 10322 9696 10378 9752
rect 10230 7248 10286 7304
rect 9402 6432 9458 6488
rect 9310 5752 9366 5808
rect 9310 5344 9366 5400
rect 9218 3304 9274 3360
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 9310 2216 9366 2272
rect 9034 1536 9090 1592
rect 10046 6704 10102 6760
rect 9954 6568 10010 6624
rect 10046 5888 10102 5944
rect 10230 5888 10286 5944
rect 9770 5480 9826 5536
rect 9678 5364 9734 5400
rect 9678 5344 9680 5364
rect 9680 5344 9732 5364
rect 9732 5344 9734 5364
rect 9770 5072 9826 5128
rect 9678 4800 9734 4856
rect 10046 5752 10102 5808
rect 9954 5344 10010 5400
rect 9954 3440 10010 3496
rect 10138 4256 10194 4312
rect 10414 9560 10470 9616
rect 10598 8880 10654 8936
rect 10817 9274 10873 9276
rect 10897 9274 10953 9276
rect 10977 9274 11033 9276
rect 11057 9274 11113 9276
rect 10817 9222 10843 9274
rect 10843 9222 10873 9274
rect 10897 9222 10907 9274
rect 10907 9222 10953 9274
rect 10977 9222 11023 9274
rect 11023 9222 11033 9274
rect 11057 9222 11087 9274
rect 11087 9222 11113 9274
rect 10817 9220 10873 9222
rect 10897 9220 10953 9222
rect 10977 9220 11033 9222
rect 11057 9220 11113 9222
rect 11058 8880 11114 8936
rect 11058 8356 11114 8392
rect 11058 8336 11060 8356
rect 11060 8336 11112 8356
rect 11112 8336 11114 8356
rect 10817 8186 10873 8188
rect 10897 8186 10953 8188
rect 10977 8186 11033 8188
rect 11057 8186 11113 8188
rect 10817 8134 10843 8186
rect 10843 8134 10873 8186
rect 10897 8134 10907 8186
rect 10907 8134 10953 8186
rect 10977 8134 11023 8186
rect 11023 8134 11033 8186
rect 11057 8134 11087 8186
rect 11087 8134 11113 8186
rect 10817 8132 10873 8134
rect 10897 8132 10953 8134
rect 10977 8132 11033 8134
rect 11057 8132 11113 8134
rect 11058 7384 11114 7440
rect 10817 7098 10873 7100
rect 10897 7098 10953 7100
rect 10977 7098 11033 7100
rect 11057 7098 11113 7100
rect 10817 7046 10843 7098
rect 10843 7046 10873 7098
rect 10897 7046 10907 7098
rect 10907 7046 10953 7098
rect 10977 7046 11023 7098
rect 11023 7046 11033 7098
rect 11057 7046 11087 7098
rect 11087 7046 11113 7098
rect 10817 7044 10873 7046
rect 10897 7044 10953 7046
rect 10977 7044 11033 7046
rect 11057 7044 11113 7046
rect 10598 6432 10654 6488
rect 10506 6060 10508 6080
rect 10508 6060 10560 6080
rect 10560 6060 10562 6080
rect 10506 6024 10562 6060
rect 10506 5616 10562 5672
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 11518 10512 11574 10568
rect 11426 10412 11428 10432
rect 11428 10412 11480 10432
rect 11480 10412 11482 10432
rect 11426 10376 11482 10412
rect 11334 9288 11390 9344
rect 11334 8336 11390 8392
rect 11242 6024 11298 6080
rect 11058 5616 11114 5672
rect 10874 5364 10930 5400
rect 10874 5344 10876 5364
rect 10876 5344 10928 5364
rect 10928 5344 10930 5364
rect 11150 5344 11206 5400
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 10598 4800 10654 4856
rect 10506 3884 10508 3904
rect 10508 3884 10560 3904
rect 10560 3884 10562 3904
rect 10506 3848 10562 3884
rect 10414 3712 10470 3768
rect 10046 2760 10102 2816
rect 9954 2624 10010 2680
rect 10230 2760 10286 2816
rect 11242 4936 11298 4992
rect 11150 4256 11206 4312
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 11426 5344 11482 5400
rect 11426 4528 11482 4584
rect 11610 8200 11666 8256
rect 11702 8064 11758 8120
rect 11610 7792 11666 7848
rect 11610 7284 11612 7304
rect 11612 7284 11664 7304
rect 11664 7284 11666 7304
rect 11610 7248 11666 7284
rect 11886 11192 11942 11248
rect 11978 10784 12034 10840
rect 11978 9832 12034 9888
rect 11978 9152 12034 9208
rect 12438 13640 12494 13696
rect 12898 16088 12954 16144
rect 13634 15544 13690 15600
rect 13282 15258 13338 15260
rect 13362 15258 13418 15260
rect 13442 15258 13498 15260
rect 13522 15258 13578 15260
rect 13282 15206 13308 15258
rect 13308 15206 13338 15258
rect 13362 15206 13372 15258
rect 13372 15206 13418 15258
rect 13442 15206 13488 15258
rect 13488 15206 13498 15258
rect 13522 15206 13552 15258
rect 13552 15206 13578 15258
rect 13282 15204 13338 15206
rect 13362 15204 13418 15206
rect 13442 15204 13498 15206
rect 13522 15204 13578 15206
rect 13174 15000 13230 15056
rect 12530 13232 12586 13288
rect 12438 13096 12494 13152
rect 12438 12008 12494 12064
rect 12438 11600 12494 11656
rect 12346 11192 12402 11248
rect 12806 14456 12862 14512
rect 12714 11872 12770 11928
rect 12438 10648 12494 10704
rect 12162 9152 12218 9208
rect 11886 8744 11942 8800
rect 11978 7792 12034 7848
rect 11150 3576 11206 3632
rect 11886 4800 11942 4856
rect 11886 4528 11942 4584
rect 11702 3848 11758 3904
rect 11426 3304 11482 3360
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 10598 2624 10654 2680
rect 11334 2624 11390 2680
rect 11242 2080 11298 2136
rect 10782 1264 10838 1320
rect 11886 3732 11942 3768
rect 11886 3712 11888 3732
rect 11888 3712 11940 3732
rect 11940 3712 11942 3732
rect 12438 9152 12494 9208
rect 12530 9016 12586 9072
rect 12162 8200 12218 8256
rect 12346 7792 12402 7848
rect 12162 7112 12218 7168
rect 11794 3168 11850 3224
rect 11794 2760 11850 2816
rect 11978 2624 12034 2680
rect 11794 2352 11850 2408
rect 12806 10920 12862 10976
rect 13266 14320 13322 14376
rect 13282 14170 13338 14172
rect 13362 14170 13418 14172
rect 13442 14170 13498 14172
rect 13522 14170 13578 14172
rect 13282 14118 13308 14170
rect 13308 14118 13338 14170
rect 13362 14118 13372 14170
rect 13372 14118 13418 14170
rect 13442 14118 13488 14170
rect 13488 14118 13498 14170
rect 13522 14118 13552 14170
rect 13552 14118 13578 14170
rect 13282 14116 13338 14118
rect 13362 14116 13418 14118
rect 13442 14116 13498 14118
rect 13522 14116 13578 14118
rect 13082 11872 13138 11928
rect 13282 13082 13338 13084
rect 13362 13082 13418 13084
rect 13442 13082 13498 13084
rect 13522 13082 13578 13084
rect 13282 13030 13308 13082
rect 13308 13030 13338 13082
rect 13362 13030 13372 13082
rect 13372 13030 13418 13082
rect 13442 13030 13488 13082
rect 13488 13030 13498 13082
rect 13522 13030 13552 13082
rect 13552 13030 13578 13082
rect 13282 13028 13338 13030
rect 13362 13028 13418 13030
rect 13442 13028 13498 13030
rect 13522 13028 13578 13030
rect 13726 13504 13782 13560
rect 13726 13232 13782 13288
rect 13450 12280 13506 12336
rect 13266 12144 13322 12200
rect 13542 12180 13544 12200
rect 13544 12180 13596 12200
rect 13596 12180 13598 12200
rect 13542 12144 13598 12180
rect 13282 11994 13338 11996
rect 13362 11994 13418 11996
rect 13442 11994 13498 11996
rect 13522 11994 13578 11996
rect 13282 11942 13308 11994
rect 13308 11942 13338 11994
rect 13362 11942 13372 11994
rect 13372 11942 13418 11994
rect 13442 11942 13488 11994
rect 13488 11942 13498 11994
rect 13522 11942 13552 11994
rect 13552 11942 13578 11994
rect 13282 11940 13338 11942
rect 13362 11940 13418 11942
rect 13442 11940 13498 11942
rect 13522 11940 13578 11942
rect 13174 11464 13230 11520
rect 12806 8472 12862 8528
rect 13266 11076 13322 11112
rect 13266 11056 13268 11076
rect 13268 11056 13320 11076
rect 13320 11056 13322 11076
rect 13634 11212 13690 11248
rect 13634 11192 13636 11212
rect 13636 11192 13688 11212
rect 13688 11192 13690 11212
rect 13282 10906 13338 10908
rect 13362 10906 13418 10908
rect 13442 10906 13498 10908
rect 13522 10906 13578 10908
rect 13282 10854 13308 10906
rect 13308 10854 13338 10906
rect 13362 10854 13372 10906
rect 13372 10854 13418 10906
rect 13442 10854 13488 10906
rect 13488 10854 13498 10906
rect 13522 10854 13552 10906
rect 13552 10854 13578 10906
rect 13282 10852 13338 10854
rect 13362 10852 13418 10854
rect 13442 10852 13498 10854
rect 13522 10852 13578 10854
rect 13174 10376 13230 10432
rect 13082 10240 13138 10296
rect 12990 9152 13046 9208
rect 13282 9818 13338 9820
rect 13362 9818 13418 9820
rect 13442 9818 13498 9820
rect 13522 9818 13578 9820
rect 13282 9766 13308 9818
rect 13308 9766 13338 9818
rect 13362 9766 13372 9818
rect 13372 9766 13418 9818
rect 13442 9766 13488 9818
rect 13488 9766 13498 9818
rect 13522 9766 13552 9818
rect 13552 9766 13578 9818
rect 13282 9764 13338 9766
rect 13362 9764 13418 9766
rect 13442 9764 13498 9766
rect 13522 9764 13578 9766
rect 13726 10104 13782 10160
rect 13634 9424 13690 9480
rect 13082 8608 13138 8664
rect 13282 8730 13338 8732
rect 13362 8730 13418 8732
rect 13442 8730 13498 8732
rect 13522 8730 13578 8732
rect 13282 8678 13308 8730
rect 13308 8678 13338 8730
rect 13362 8678 13372 8730
rect 13372 8678 13418 8730
rect 13442 8678 13488 8730
rect 13488 8678 13498 8730
rect 13522 8678 13552 8730
rect 13552 8678 13578 8730
rect 13282 8676 13338 8678
rect 13362 8676 13418 8678
rect 13442 8676 13498 8678
rect 13522 8676 13578 8678
rect 13282 7642 13338 7644
rect 13362 7642 13418 7644
rect 13442 7642 13498 7644
rect 13522 7642 13578 7644
rect 13282 7590 13308 7642
rect 13308 7590 13338 7642
rect 13362 7590 13372 7642
rect 13372 7590 13418 7642
rect 13442 7590 13488 7642
rect 13488 7590 13498 7642
rect 13522 7590 13552 7642
rect 13552 7590 13578 7642
rect 13282 7588 13338 7590
rect 13362 7588 13418 7590
rect 13442 7588 13498 7590
rect 13522 7588 13578 7590
rect 13266 7420 13268 7440
rect 13268 7420 13320 7440
rect 13320 7420 13322 7440
rect 13266 7384 13322 7420
rect 13266 7248 13322 7304
rect 13174 7112 13230 7168
rect 13358 6976 13414 7032
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 12438 6060 12440 6080
rect 12440 6060 12492 6080
rect 12492 6060 12494 6080
rect 12438 6024 12494 6060
rect 12346 5616 12402 5672
rect 12254 5344 12310 5400
rect 12806 6024 12862 6080
rect 12530 4800 12586 4856
rect 12438 4156 12440 4176
rect 12440 4156 12492 4176
rect 12492 4156 12494 4176
rect 12438 4120 12494 4156
rect 12530 3984 12586 4040
rect 12346 3440 12402 3496
rect 12714 5480 12770 5536
rect 12714 3168 12770 3224
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 13910 9696 13966 9752
rect 13818 8336 13874 8392
rect 13818 7928 13874 7984
rect 14186 13368 14242 13424
rect 14186 12688 14242 12744
rect 14554 14864 14610 14920
rect 14370 13776 14426 13832
rect 14002 8064 14058 8120
rect 14278 9288 14334 9344
rect 14186 8744 14242 8800
rect 14094 7928 14150 7984
rect 13818 4936 13874 4992
rect 13082 3304 13138 3360
rect 13082 2624 13138 2680
rect 13082 2352 13138 2408
rect 12530 1536 12586 1592
rect 13082 2216 13138 2272
rect 13450 3612 13452 3632
rect 13452 3612 13504 3632
rect 13504 3612 13506 3632
rect 13450 3576 13506 3612
rect 13358 3440 13414 3496
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 13818 3712 13874 3768
rect 13818 3440 13874 3496
rect 13726 3032 13782 3088
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
rect 13358 1944 13414 2000
rect 14922 14456 14978 14512
rect 14738 10512 14794 10568
rect 14646 9988 14702 10024
rect 14646 9968 14648 9988
rect 14648 9968 14700 9988
rect 14700 9968 14702 9988
rect 14094 5228 14150 5264
rect 14094 5208 14096 5228
rect 14096 5208 14148 5228
rect 14148 5208 14150 5228
rect 14186 4528 14242 4584
rect 14462 6704 14518 6760
rect 14738 8200 14794 8256
rect 14462 3984 14518 4040
rect 14646 4120 14702 4176
rect 14554 2760 14610 2816
rect 15014 13948 15016 13968
rect 15016 13948 15068 13968
rect 15068 13948 15070 13968
rect 15014 13912 15070 13948
rect 15014 9596 15016 9616
rect 15016 9596 15068 9616
rect 15068 9596 15070 9616
rect 15014 9560 15070 9596
rect 15014 6332 15016 6352
rect 15016 6332 15068 6352
rect 15068 6332 15070 6352
rect 15014 6296 15070 6332
rect 14922 4120 14978 4176
rect 15014 2896 15070 2952
rect 15382 4120 15438 4176
rect 16762 6840 16818 6896
<< metal3 >>
rect 0 17370 480 17400
rect 1945 17370 2011 17373
rect 0 17368 2011 17370
rect 0 17312 1950 17368
rect 2006 17312 2011 17368
rect 0 17310 2011 17312
rect 0 17280 480 17310
rect 1945 17307 2011 17310
rect 0 16282 480 16312
rect 4061 16282 4127 16285
rect 0 16280 4127 16282
rect 0 16224 4066 16280
rect 4122 16224 4127 16280
rect 0 16222 4127 16224
rect 0 16192 480 16222
rect 4061 16219 4127 16222
rect 12382 16084 12388 16148
rect 12452 16146 12458 16148
rect 12893 16146 12959 16149
rect 12452 16144 12959 16146
rect 12452 16088 12898 16144
rect 12954 16088 12959 16144
rect 12452 16086 12959 16088
rect 12452 16084 12458 16086
rect 12893 16083 12959 16086
rect 7465 16010 7531 16013
rect 11513 16010 11579 16013
rect 7465 16008 11579 16010
rect 7465 15952 7470 16008
rect 7526 15952 11518 16008
rect 11574 15952 11579 16008
rect 7465 15950 11579 15952
rect 7465 15947 7531 15950
rect 11513 15947 11579 15950
rect 5874 15808 6194 15809
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6194 15808
rect 5874 15743 6194 15744
rect 10805 15808 11125 15809
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 15743 11125 15744
rect 6862 15676 6868 15740
rect 6932 15738 6938 15740
rect 6932 15678 9138 15738
rect 6932 15676 6938 15678
rect 8937 15602 9003 15605
rect 3236 15600 9003 15602
rect 3236 15544 8942 15600
rect 8998 15544 9003 15600
rect 3236 15542 9003 15544
rect 9078 15602 9138 15678
rect 13629 15602 13695 15605
rect 9078 15600 13695 15602
rect 9078 15544 13634 15600
rect 13690 15544 13695 15600
rect 9078 15542 13695 15544
rect 0 15194 480 15224
rect 3236 15194 3296 15542
rect 8937 15539 9003 15542
rect 13629 15539 13695 15542
rect 4061 15466 4127 15469
rect 9213 15466 9279 15469
rect 4061 15464 9279 15466
rect 4061 15408 4066 15464
rect 4122 15408 9218 15464
rect 9274 15408 9279 15464
rect 4061 15406 9279 15408
rect 4061 15403 4127 15406
rect 9213 15403 9279 15406
rect 6821 15330 6887 15333
rect 8201 15330 8267 15333
rect 6821 15328 8267 15330
rect 6821 15272 6826 15328
rect 6882 15272 8206 15328
rect 8262 15272 8267 15328
rect 6821 15270 8267 15272
rect 6821 15267 6887 15270
rect 8201 15267 8267 15270
rect 3409 15264 3729 15265
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 15199 3729 15200
rect 8340 15264 8660 15265
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 15199 8660 15200
rect 13270 15264 13590 15265
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 15199 13590 15200
rect 0 15134 3296 15194
rect 5625 15194 5691 15197
rect 6862 15194 6868 15196
rect 5625 15192 6868 15194
rect 5625 15136 5630 15192
rect 5686 15136 6868 15192
rect 5625 15134 6868 15136
rect 0 15104 480 15134
rect 5625 15131 5691 15134
rect 6862 15132 6868 15134
rect 6932 15194 6938 15196
rect 7097 15194 7163 15197
rect 6932 15192 7163 15194
rect 6932 15136 7102 15192
rect 7158 15136 7163 15192
rect 6932 15134 7163 15136
rect 6932 15132 6938 15134
rect 7097 15131 7163 15134
rect 9305 15194 9371 15197
rect 11697 15194 11763 15197
rect 9305 15192 11763 15194
rect 9305 15136 9310 15192
rect 9366 15136 11702 15192
rect 11758 15136 11763 15192
rect 9305 15134 11763 15136
rect 9305 15131 9371 15134
rect 11697 15131 11763 15134
rect 4061 15058 4127 15061
rect 12198 15058 12204 15060
rect 4061 15056 12204 15058
rect 4061 15000 4066 15056
rect 4122 15000 12204 15056
rect 4061 14998 12204 15000
rect 4061 14995 4127 14998
rect 12198 14996 12204 14998
rect 12268 15058 12274 15060
rect 13169 15058 13235 15061
rect 12268 15056 13235 15058
rect 12268 15000 13174 15056
rect 13230 15000 13235 15056
rect 12268 14998 13235 15000
rect 12268 14996 12274 14998
rect 13169 14995 13235 14998
rect 1025 14922 1091 14925
rect 14549 14922 14615 14925
rect 1025 14920 14615 14922
rect 1025 14864 1030 14920
rect 1086 14864 14554 14920
rect 14610 14864 14615 14920
rect 1025 14862 14615 14864
rect 1025 14859 1091 14862
rect 14549 14859 14615 14862
rect 5206 14724 5212 14788
rect 5276 14786 5282 14788
rect 5441 14786 5507 14789
rect 5276 14784 5507 14786
rect 5276 14728 5446 14784
rect 5502 14728 5507 14784
rect 5276 14726 5507 14728
rect 5276 14724 5282 14726
rect 5441 14723 5507 14726
rect 6269 14786 6335 14789
rect 7649 14786 7715 14789
rect 9121 14786 9187 14789
rect 9622 14786 9628 14788
rect 6269 14784 9628 14786
rect 6269 14728 6274 14784
rect 6330 14728 7654 14784
rect 7710 14728 9126 14784
rect 9182 14728 9628 14784
rect 6269 14726 9628 14728
rect 6269 14723 6335 14726
rect 7649 14723 7715 14726
rect 9121 14723 9187 14726
rect 9622 14724 9628 14726
rect 9692 14724 9698 14788
rect 9990 14724 9996 14788
rect 10060 14786 10066 14788
rect 10409 14786 10475 14789
rect 10060 14784 10475 14786
rect 10060 14728 10414 14784
rect 10470 14728 10475 14784
rect 10060 14726 10475 14728
rect 10060 14724 10066 14726
rect 10409 14723 10475 14726
rect 11646 14724 11652 14788
rect 11716 14786 11722 14788
rect 11789 14786 11855 14789
rect 11716 14784 11855 14786
rect 11716 14728 11794 14784
rect 11850 14728 11855 14784
rect 11716 14726 11855 14728
rect 11716 14724 11722 14726
rect 11789 14723 11855 14726
rect 5874 14720 6194 14721
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6194 14720
rect 5874 14655 6194 14656
rect 10805 14720 11125 14721
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 14655 11125 14656
rect 4245 14650 4311 14653
rect 5574 14650 5580 14652
rect 4245 14648 5580 14650
rect 4245 14592 4250 14648
rect 4306 14592 5580 14648
rect 4245 14590 5580 14592
rect 4245 14587 4311 14590
rect 5574 14588 5580 14590
rect 5644 14588 5650 14652
rect 6310 14588 6316 14652
rect 6380 14650 6386 14652
rect 6729 14650 6795 14653
rect 6380 14648 6795 14650
rect 6380 14592 6734 14648
rect 6790 14592 6795 14648
rect 6380 14590 6795 14592
rect 6380 14588 6386 14590
rect 6729 14587 6795 14590
rect 7189 14650 7255 14653
rect 8937 14650 9003 14653
rect 7189 14648 9003 14650
rect 7189 14592 7194 14648
rect 7250 14592 8942 14648
rect 8998 14592 9003 14648
rect 7189 14590 9003 14592
rect 7189 14587 7255 14590
rect 8937 14587 9003 14590
rect 9489 14650 9555 14653
rect 10409 14650 10475 14653
rect 9489 14648 10475 14650
rect 9489 14592 9494 14648
rect 9550 14592 10414 14648
rect 10470 14592 10475 14648
rect 9489 14590 10475 14592
rect 9489 14587 9555 14590
rect 10409 14587 10475 14590
rect 3969 14514 4035 14517
rect 8661 14514 8727 14517
rect 9673 14514 9739 14517
rect 12341 14514 12407 14517
rect 12801 14514 12867 14517
rect 14917 14514 14983 14517
rect 3969 14512 9874 14514
rect 3969 14456 3974 14512
rect 4030 14456 8666 14512
rect 8722 14456 9678 14512
rect 9734 14456 9874 14512
rect 3969 14454 9874 14456
rect 3969 14451 4035 14454
rect 8661 14451 8727 14454
rect 9673 14451 9739 14454
rect 1485 14378 1551 14381
rect 7598 14378 7604 14380
rect 1485 14376 7604 14378
rect 1485 14320 1490 14376
rect 1546 14320 7604 14376
rect 1485 14318 7604 14320
rect 1485 14315 1551 14318
rect 7598 14316 7604 14318
rect 7668 14316 7674 14380
rect 7833 14378 7899 14381
rect 9814 14378 9874 14454
rect 12341 14512 12867 14514
rect 12341 14456 12346 14512
rect 12402 14456 12806 14512
rect 12862 14456 12867 14512
rect 12341 14454 12867 14456
rect 12341 14451 12407 14454
rect 12801 14451 12867 14454
rect 12942 14512 14983 14514
rect 12942 14456 14922 14512
rect 14978 14456 14983 14512
rect 12942 14454 14983 14456
rect 12942 14378 13002 14454
rect 14917 14451 14983 14454
rect 7833 14376 9736 14378
rect 7833 14320 7838 14376
rect 7894 14320 9736 14376
rect 7833 14318 9736 14320
rect 9814 14318 13002 14378
rect 7833 14315 7899 14318
rect 5390 14180 5396 14244
rect 5460 14242 5466 14244
rect 5901 14242 5967 14245
rect 5460 14240 5967 14242
rect 5460 14184 5906 14240
rect 5962 14184 5967 14240
rect 5460 14182 5967 14184
rect 9676 14242 9736 14318
rect 13118 14316 13124 14380
rect 13188 14378 13194 14380
rect 13261 14378 13327 14381
rect 13188 14376 13327 14378
rect 13188 14320 13266 14376
rect 13322 14320 13327 14376
rect 13188 14318 13327 14320
rect 13188 14316 13194 14318
rect 13261 14315 13327 14318
rect 9857 14242 9923 14245
rect 12065 14242 12131 14245
rect 9676 14240 12131 14242
rect 9676 14184 9862 14240
rect 9918 14184 12070 14240
rect 12126 14184 12131 14240
rect 9676 14182 12131 14184
rect 5460 14180 5466 14182
rect 5901 14179 5967 14182
rect 9857 14179 9923 14182
rect 12065 14179 12131 14182
rect 3409 14176 3729 14177
rect 0 14106 480 14136
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 14111 3729 14112
rect 8340 14176 8660 14177
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 14111 8660 14112
rect 13270 14176 13590 14177
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 14111 13590 14112
rect 3049 14106 3115 14109
rect 0 14104 3115 14106
rect 0 14048 3054 14104
rect 3110 14048 3115 14104
rect 0 14046 3115 14048
rect 0 14016 480 14046
rect 3049 14043 3115 14046
rect 3969 14106 4035 14109
rect 8201 14106 8267 14109
rect 3969 14104 8267 14106
rect 3969 14048 3974 14104
rect 4030 14048 8206 14104
rect 8262 14048 8267 14104
rect 3969 14046 8267 14048
rect 3969 14043 4035 14046
rect 8201 14043 8267 14046
rect 8845 14106 8911 14109
rect 9305 14106 9371 14109
rect 8845 14104 9371 14106
rect 8845 14048 8850 14104
rect 8906 14048 9310 14104
rect 9366 14048 9371 14104
rect 8845 14046 9371 14048
rect 8845 14043 8911 14046
rect 9305 14043 9371 14046
rect 9622 14044 9628 14108
rect 9692 14106 9698 14108
rect 12341 14106 12407 14109
rect 9692 14104 12407 14106
rect 9692 14048 12346 14104
rect 12402 14048 12407 14104
rect 9692 14046 12407 14048
rect 9692 14044 9698 14046
rect 12341 14043 12407 14046
rect 4153 13970 4219 13973
rect 4429 13970 4495 13973
rect 4153 13968 4495 13970
rect 4153 13912 4158 13968
rect 4214 13912 4434 13968
rect 4490 13912 4495 13968
rect 4153 13910 4495 13912
rect 4153 13907 4219 13910
rect 4429 13907 4495 13910
rect 4613 13970 4679 13973
rect 6361 13970 6427 13973
rect 4613 13968 6427 13970
rect 4613 13912 4618 13968
rect 4674 13912 6366 13968
rect 6422 13912 6427 13968
rect 4613 13910 6427 13912
rect 4613 13907 4679 13910
rect 6361 13907 6427 13910
rect 6637 13970 6703 13973
rect 15009 13970 15075 13973
rect 6637 13968 15075 13970
rect 6637 13912 6642 13968
rect 6698 13912 15014 13968
rect 15070 13912 15075 13968
rect 6637 13910 15075 13912
rect 6637 13907 6703 13910
rect 15009 13907 15075 13910
rect 2405 13834 2471 13837
rect 2405 13832 6378 13834
rect 2405 13776 2410 13832
rect 2466 13776 6378 13832
rect 2405 13774 6378 13776
rect 2405 13771 2471 13774
rect 4521 13698 4587 13701
rect 5717 13698 5783 13701
rect 4521 13696 5783 13698
rect 4521 13640 4526 13696
rect 4582 13640 5722 13696
rect 5778 13640 5783 13696
rect 4521 13638 5783 13640
rect 4521 13635 4587 13638
rect 5717 13635 5783 13638
rect 5874 13632 6194 13633
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6194 13632
rect 5874 13567 6194 13568
rect 4613 13562 4679 13565
rect 5441 13562 5507 13565
rect 4613 13560 5507 13562
rect 4613 13504 4618 13560
rect 4674 13504 5446 13560
rect 5502 13504 5507 13560
rect 4613 13502 5507 13504
rect 6318 13562 6378 13774
rect 8150 13772 8156 13836
rect 8220 13834 8226 13836
rect 14365 13834 14431 13837
rect 8220 13832 14431 13834
rect 8220 13776 14370 13832
rect 14426 13776 14431 13832
rect 8220 13774 14431 13776
rect 8220 13772 8226 13774
rect 14365 13771 14431 13774
rect 6678 13636 6684 13700
rect 6748 13698 6754 13700
rect 7005 13698 7071 13701
rect 6748 13696 7071 13698
rect 6748 13640 7010 13696
rect 7066 13640 7071 13696
rect 6748 13638 7071 13640
rect 6748 13636 6754 13638
rect 7005 13635 7071 13638
rect 7741 13698 7807 13701
rect 11237 13698 11303 13701
rect 12157 13698 12223 13701
rect 7741 13696 10564 13698
rect 7741 13640 7746 13696
rect 7802 13640 10564 13696
rect 7741 13638 10564 13640
rect 7741 13635 7807 13638
rect 10504 13565 10564 13638
rect 11237 13696 12223 13698
rect 11237 13640 11242 13696
rect 11298 13640 12162 13696
rect 12218 13640 12223 13696
rect 11237 13638 12223 13640
rect 11237 13635 11303 13638
rect 12157 13635 12223 13638
rect 12433 13698 12499 13701
rect 12566 13698 12572 13700
rect 12433 13696 12572 13698
rect 12433 13640 12438 13696
rect 12494 13640 12572 13696
rect 12433 13638 12572 13640
rect 12433 13635 12499 13638
rect 12566 13636 12572 13638
rect 12636 13636 12642 13700
rect 10805 13632 11125 13633
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 13567 11125 13568
rect 9029 13562 9095 13565
rect 9857 13564 9923 13565
rect 6318 13560 9095 13562
rect 6318 13504 9034 13560
rect 9090 13504 9095 13560
rect 6318 13502 9095 13504
rect 4613 13499 4679 13502
rect 5441 13499 5507 13502
rect 9029 13499 9095 13502
rect 9806 13500 9812 13564
rect 9876 13562 9923 13564
rect 10501 13564 10567 13565
rect 10501 13562 10548 13564
rect 9876 13560 9968 13562
rect 9918 13504 9968 13560
rect 9876 13502 9968 13504
rect 10456 13560 10548 13562
rect 10456 13504 10506 13560
rect 10456 13502 10548 13504
rect 9876 13500 9923 13502
rect 9857 13499 9923 13500
rect 10501 13500 10548 13502
rect 10612 13500 10618 13564
rect 11605 13562 11671 13565
rect 11830 13562 11836 13564
rect 11605 13560 11836 13562
rect 11605 13504 11610 13560
rect 11666 13504 11836 13560
rect 11605 13502 11836 13504
rect 10501 13499 10567 13500
rect 11605 13499 11671 13502
rect 11830 13500 11836 13502
rect 11900 13500 11906 13564
rect 12014 13500 12020 13564
rect 12084 13562 12090 13564
rect 13721 13562 13787 13565
rect 16520 13562 17000 13592
rect 12084 13560 17000 13562
rect 12084 13504 13726 13560
rect 13782 13504 17000 13560
rect 12084 13502 17000 13504
rect 12084 13500 12090 13502
rect 13721 13499 13787 13502
rect 16520 13472 17000 13502
rect 1853 13426 1919 13429
rect 8293 13426 8359 13429
rect 1853 13424 8359 13426
rect 1853 13368 1858 13424
rect 1914 13368 8298 13424
rect 8354 13368 8359 13424
rect 1853 13366 8359 13368
rect 1853 13363 1919 13366
rect 8293 13363 8359 13366
rect 9305 13426 9371 13429
rect 10501 13426 10567 13429
rect 14181 13426 14247 13429
rect 9305 13424 14247 13426
rect 9305 13368 9310 13424
rect 9366 13368 10506 13424
rect 10562 13368 14186 13424
rect 14242 13368 14247 13424
rect 9305 13366 14247 13368
rect 9305 13363 9371 13366
rect 10501 13363 10567 13366
rect 14181 13363 14247 13366
rect 3049 13290 3115 13293
rect 5257 13290 5323 13293
rect 11973 13290 12039 13293
rect 3049 13288 4906 13290
rect 3049 13232 3054 13288
rect 3110 13232 4906 13288
rect 3049 13230 4906 13232
rect 3049 13227 3115 13230
rect 0 13154 480 13184
rect 0 13094 3296 13154
rect 0 13064 480 13094
rect 3236 12882 3296 13094
rect 3409 13088 3729 13089
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 13023 3729 13024
rect 4153 13018 4219 13021
rect 4705 13018 4771 13021
rect 4153 13016 4771 13018
rect 4153 12960 4158 13016
rect 4214 12960 4710 13016
rect 4766 12960 4771 13016
rect 4153 12958 4771 12960
rect 4846 13018 4906 13230
rect 5257 13288 12039 13290
rect 5257 13232 5262 13288
rect 5318 13232 11978 13288
rect 12034 13232 12039 13288
rect 5257 13230 12039 13232
rect 5257 13227 5323 13230
rect 11973 13227 12039 13230
rect 12525 13290 12591 13293
rect 13721 13290 13787 13293
rect 12525 13288 13787 13290
rect 12525 13232 12530 13288
rect 12586 13232 13726 13288
rect 13782 13232 13787 13288
rect 12525 13230 13787 13232
rect 12525 13227 12591 13230
rect 13721 13227 13787 13230
rect 5574 13092 5580 13156
rect 5644 13154 5650 13156
rect 8201 13154 8267 13157
rect 5644 13152 8267 13154
rect 5644 13096 8206 13152
rect 8262 13096 8267 13152
rect 5644 13094 8267 13096
rect 5644 13092 5650 13094
rect 8201 13091 8267 13094
rect 8753 13154 8819 13157
rect 12433 13154 12499 13157
rect 8753 13152 12499 13154
rect 8753 13096 8758 13152
rect 8814 13096 12438 13152
rect 12494 13096 12499 13152
rect 8753 13094 12499 13096
rect 8753 13091 8819 13094
rect 12433 13091 12499 13094
rect 8340 13088 8660 13089
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 13023 8660 13024
rect 13270 13088 13590 13089
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 13023 13590 13024
rect 4846 12958 6792 13018
rect 4153 12955 4219 12958
rect 4705 12955 4771 12958
rect 5349 12882 5415 12885
rect 3236 12880 5415 12882
rect 3236 12824 5354 12880
rect 5410 12824 5415 12880
rect 3236 12822 5415 12824
rect 5349 12819 5415 12822
rect 5533 12882 5599 12885
rect 6085 12882 6151 12885
rect 6545 12884 6611 12885
rect 6494 12882 6500 12884
rect 5533 12880 6151 12882
rect 5533 12824 5538 12880
rect 5594 12824 6090 12880
rect 6146 12824 6151 12880
rect 5533 12822 6151 12824
rect 6454 12822 6500 12882
rect 6564 12880 6611 12884
rect 6606 12824 6611 12880
rect 5533 12819 5599 12822
rect 6085 12819 6151 12822
rect 6494 12820 6500 12822
rect 6564 12820 6611 12824
rect 6732 12882 6792 12958
rect 7414 12956 7420 13020
rect 7484 13018 7490 13020
rect 8017 13018 8083 13021
rect 7484 13016 8083 13018
rect 7484 12960 8022 13016
rect 8078 12960 8083 13016
rect 7484 12958 8083 12960
rect 7484 12956 7490 12958
rect 8017 12955 8083 12958
rect 8937 13018 9003 13021
rect 9254 13018 9260 13020
rect 8937 13016 9260 13018
rect 8937 12960 8942 13016
rect 8998 12960 9260 13016
rect 8937 12958 9260 12960
rect 8937 12955 9003 12958
rect 9254 12956 9260 12958
rect 9324 12956 9330 13020
rect 9857 13018 9923 13021
rect 10174 13018 10180 13020
rect 9857 13016 10180 13018
rect 9857 12960 9862 13016
rect 9918 12960 10180 13016
rect 9857 12958 10180 12960
rect 9857 12955 9923 12958
rect 10174 12956 10180 12958
rect 10244 13018 10250 13020
rect 11237 13018 11303 13021
rect 10244 13016 11303 13018
rect 10244 12960 11242 13016
rect 11298 12960 11303 13016
rect 10244 12958 11303 12960
rect 10244 12956 10250 12958
rect 11237 12955 11303 12958
rect 7741 12882 7807 12885
rect 6732 12880 7807 12882
rect 6732 12824 7746 12880
rect 7802 12824 7807 12880
rect 6732 12822 7807 12824
rect 6545 12819 6611 12820
rect 7741 12819 7807 12822
rect 8109 12882 8175 12885
rect 11278 12882 11284 12884
rect 8109 12880 11284 12882
rect 8109 12824 8114 12880
rect 8170 12824 11284 12880
rect 8109 12822 11284 12824
rect 8109 12819 8175 12822
rect 11278 12820 11284 12822
rect 11348 12820 11354 12884
rect 4337 12746 4403 12749
rect 14181 12746 14247 12749
rect 4337 12744 14247 12746
rect 4337 12688 4342 12744
rect 4398 12688 14186 12744
rect 14242 12688 14247 12744
rect 4337 12686 14247 12688
rect 4337 12683 4403 12686
rect 14181 12683 14247 12686
rect 3601 12610 3667 12613
rect 5717 12610 5783 12613
rect 3601 12608 5783 12610
rect 3601 12552 3606 12608
rect 3662 12552 5722 12608
rect 5778 12552 5783 12608
rect 3601 12550 5783 12552
rect 3601 12547 3667 12550
rect 5717 12547 5783 12550
rect 6729 12610 6795 12613
rect 9438 12610 9444 12612
rect 6729 12608 9444 12610
rect 6729 12552 6734 12608
rect 6790 12552 9444 12608
rect 6729 12550 9444 12552
rect 6729 12547 6795 12550
rect 9438 12548 9444 12550
rect 9508 12548 9514 12612
rect 10358 12548 10364 12612
rect 10428 12610 10434 12612
rect 10501 12610 10567 12613
rect 10428 12608 10567 12610
rect 10428 12552 10506 12608
rect 10562 12552 10567 12608
rect 10428 12550 10567 12552
rect 10428 12548 10434 12550
rect 10501 12547 10567 12550
rect 5874 12544 6194 12545
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6194 12544
rect 5874 12479 6194 12480
rect 10805 12544 11125 12545
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 12479 11125 12480
rect 1945 12474 2011 12477
rect 4061 12474 4127 12477
rect 1945 12472 4127 12474
rect 1945 12416 1950 12472
rect 2006 12416 4066 12472
rect 4122 12416 4127 12472
rect 1945 12414 4127 12416
rect 1945 12411 2011 12414
rect 4061 12411 4127 12414
rect 4838 12412 4844 12476
rect 4908 12474 4914 12476
rect 5533 12474 5599 12477
rect 4908 12472 5599 12474
rect 4908 12416 5538 12472
rect 5594 12416 5599 12472
rect 4908 12414 5599 12416
rect 4908 12412 4914 12414
rect 5533 12411 5599 12414
rect 6361 12474 6427 12477
rect 9305 12474 9371 12477
rect 6361 12472 9371 12474
rect 6361 12416 6366 12472
rect 6422 12416 9310 12472
rect 9366 12416 9371 12472
rect 6361 12414 9371 12416
rect 6361 12411 6427 12414
rect 9305 12411 9371 12414
rect 2221 12338 2287 12341
rect 4286 12338 4292 12340
rect 2221 12336 4292 12338
rect 2221 12280 2226 12336
rect 2282 12280 4292 12336
rect 2221 12278 4292 12280
rect 2221 12275 2287 12278
rect 4286 12276 4292 12278
rect 4356 12276 4362 12340
rect 7373 12338 7439 12341
rect 7557 12338 7623 12341
rect 13445 12338 13511 12341
rect 5214 12336 7623 12338
rect 5214 12280 7378 12336
rect 7434 12280 7562 12336
rect 7618 12280 7623 12336
rect 5214 12278 7623 12280
rect 2865 12202 2931 12205
rect 2998 12202 3004 12204
rect 2865 12200 3004 12202
rect 2865 12144 2870 12200
rect 2926 12144 3004 12200
rect 2865 12142 3004 12144
rect 2865 12139 2931 12142
rect 2998 12140 3004 12142
rect 3068 12202 3074 12204
rect 4061 12202 4127 12205
rect 5214 12202 5274 12278
rect 7373 12275 7439 12278
rect 7557 12275 7623 12278
rect 10136 12336 13511 12338
rect 10136 12280 13450 12336
rect 13506 12280 13511 12336
rect 10136 12278 13511 12280
rect 3068 12142 3986 12202
rect 3068 12140 3074 12142
rect 0 12066 480 12096
rect 0 12006 3296 12066
rect 0 11976 480 12006
rect 3236 11794 3296 12006
rect 3409 12000 3729 12001
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 11935 3729 11936
rect 3926 11930 3986 12142
rect 4061 12200 5274 12202
rect 4061 12144 4066 12200
rect 4122 12144 5274 12200
rect 4061 12142 5274 12144
rect 5349 12202 5415 12205
rect 8020 12202 8218 12236
rect 10136 12202 10196 12278
rect 13445 12275 13511 12278
rect 5349 12200 10196 12202
rect 5349 12144 5354 12200
rect 5410 12176 10196 12200
rect 5410 12144 8080 12176
rect 5349 12142 8080 12144
rect 8158 12142 10196 12176
rect 10777 12202 10843 12205
rect 13261 12202 13327 12205
rect 10777 12200 13327 12202
rect 10777 12144 10782 12200
rect 10838 12144 13266 12200
rect 13322 12144 13327 12200
rect 10777 12142 13327 12144
rect 4061 12139 4127 12142
rect 5349 12139 5415 12142
rect 10777 12139 10843 12142
rect 13261 12139 13327 12142
rect 13537 12202 13603 12205
rect 13537 12200 13738 12202
rect 13537 12144 13542 12200
rect 13598 12144 13738 12200
rect 13537 12142 13738 12144
rect 13537 12139 13603 12142
rect 4889 12066 4955 12069
rect 5349 12066 5415 12069
rect 7414 12066 7420 12068
rect 4889 12064 7420 12066
rect 4889 12008 4894 12064
rect 4950 12008 5354 12064
rect 5410 12008 7420 12064
rect 4889 12006 7420 12008
rect 4889 12003 4955 12006
rect 5349 12003 5415 12006
rect 7414 12004 7420 12006
rect 7484 12004 7490 12068
rect 8753 12066 8819 12069
rect 11329 12066 11395 12069
rect 8753 12064 11395 12066
rect 8753 12008 8758 12064
rect 8814 12008 11334 12064
rect 11390 12008 11395 12064
rect 8753 12006 11395 12008
rect 8753 12003 8819 12006
rect 11329 12003 11395 12006
rect 12433 12066 12499 12069
rect 12433 12064 13140 12066
rect 12433 12008 12438 12064
rect 12494 12008 13140 12064
rect 12433 12006 13140 12008
rect 12433 12003 12499 12006
rect 8340 12000 8660 12001
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 11935 8660 11936
rect 13080 11933 13140 12006
rect 13270 12000 13590 12001
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 11935 13590 11936
rect 8109 11930 8175 11933
rect 3926 11928 8175 11930
rect 3926 11872 8114 11928
rect 8170 11872 8175 11928
rect 3926 11870 8175 11872
rect 8109 11867 8175 11870
rect 9070 11868 9076 11932
rect 9140 11930 9146 11932
rect 12709 11930 12775 11933
rect 9140 11928 12775 11930
rect 9140 11872 12714 11928
rect 12770 11872 12775 11928
rect 9140 11870 12775 11872
rect 9140 11868 9146 11870
rect 12709 11867 12775 11870
rect 13077 11928 13143 11933
rect 13077 11872 13082 11928
rect 13138 11872 13143 11928
rect 13077 11867 13143 11872
rect 13678 11794 13738 12142
rect 3236 11734 13738 11794
rect 2773 11658 2839 11661
rect 12433 11658 12499 11661
rect 2773 11656 12499 11658
rect 2773 11600 2778 11656
rect 2834 11600 12438 11656
rect 12494 11600 12499 11656
rect 2773 11598 12499 11600
rect 2773 11595 2839 11598
rect 12433 11595 12499 11598
rect 2681 11522 2747 11525
rect 3417 11522 3483 11525
rect 2681 11520 3483 11522
rect 2681 11464 2686 11520
rect 2742 11464 3422 11520
rect 3478 11464 3483 11520
rect 2681 11462 3483 11464
rect 2681 11459 2747 11462
rect 3417 11459 3483 11462
rect 5073 11522 5139 11525
rect 5717 11522 5783 11525
rect 5073 11520 5783 11522
rect 5073 11464 5078 11520
rect 5134 11464 5722 11520
rect 5778 11464 5783 11520
rect 5073 11462 5783 11464
rect 5073 11459 5139 11462
rect 5717 11459 5783 11462
rect 6310 11460 6316 11524
rect 6380 11522 6386 11524
rect 6453 11522 6519 11525
rect 6380 11520 6519 11522
rect 6380 11464 6458 11520
rect 6514 11464 6519 11520
rect 6380 11462 6519 11464
rect 6380 11460 6386 11462
rect 6453 11459 6519 11462
rect 7097 11522 7163 11525
rect 7557 11522 7623 11525
rect 7097 11520 7623 11522
rect 7097 11464 7102 11520
rect 7158 11464 7562 11520
rect 7618 11464 7623 11520
rect 7097 11462 7623 11464
rect 7097 11459 7163 11462
rect 7557 11459 7623 11462
rect 7966 11460 7972 11524
rect 8036 11522 8042 11524
rect 10593 11522 10659 11525
rect 13169 11522 13235 11525
rect 8036 11520 10659 11522
rect 8036 11464 10598 11520
rect 10654 11464 10659 11520
rect 8036 11462 10659 11464
rect 8036 11460 8042 11462
rect 10593 11459 10659 11462
rect 11240 11520 13235 11522
rect 11240 11464 13174 11520
rect 13230 11464 13235 11520
rect 11240 11462 13235 11464
rect 5874 11456 6194 11457
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6194 11456
rect 5874 11391 6194 11392
rect 10805 11456 11125 11457
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 11391 11125 11392
rect 2681 11386 2747 11389
rect 5717 11386 5783 11389
rect 2681 11384 5783 11386
rect 2681 11328 2686 11384
rect 2742 11328 5722 11384
rect 5778 11328 5783 11384
rect 2681 11326 5783 11328
rect 2681 11323 2747 11326
rect 5717 11323 5783 11326
rect 6310 11324 6316 11388
rect 6380 11386 6386 11388
rect 6380 11326 9000 11386
rect 6380 11324 6386 11326
rect 2037 11250 2103 11253
rect 8748 11250 8754 11252
rect 2037 11248 8754 11250
rect 2037 11192 2042 11248
rect 2098 11192 8754 11248
rect 2037 11190 8754 11192
rect 2037 11187 2103 11190
rect 8748 11188 8754 11190
rect 8818 11188 8824 11252
rect 8940 11250 9000 11326
rect 11240 11253 11300 11462
rect 13169 11459 13235 11462
rect 8940 11190 10932 11250
rect 2865 11114 2931 11117
rect 5533 11114 5599 11117
rect 10685 11114 10751 11117
rect 2865 11112 3986 11114
rect 2865 11056 2870 11112
rect 2926 11056 3986 11112
rect 2865 11054 3986 11056
rect 2865 11051 2931 11054
rect 0 10978 480 11008
rect 0 10918 3112 10978
rect 0 10888 480 10918
rect 3052 10706 3112 10918
rect 3409 10912 3729 10913
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 10847 3729 10848
rect 3926 10842 3986 11054
rect 5533 11112 10751 11114
rect 5533 11056 5538 11112
rect 5594 11056 10690 11112
rect 10746 11056 10751 11112
rect 5533 11054 10751 11056
rect 10872 11114 10932 11190
rect 11237 11248 11303 11253
rect 11881 11252 11947 11253
rect 11237 11192 11242 11248
rect 11298 11192 11303 11248
rect 11237 11187 11303 11192
rect 11830 11188 11836 11252
rect 11900 11250 11947 11252
rect 12341 11250 12407 11253
rect 13629 11250 13695 11253
rect 11900 11248 11992 11250
rect 11942 11192 11992 11248
rect 11900 11190 11992 11192
rect 12341 11248 13695 11250
rect 12341 11192 12346 11248
rect 12402 11192 13634 11248
rect 13690 11192 13695 11248
rect 12341 11190 13695 11192
rect 11900 11188 11947 11190
rect 11881 11187 11947 11188
rect 12341 11187 12407 11190
rect 13629 11187 13695 11190
rect 13261 11114 13327 11117
rect 10872 11112 13327 11114
rect 10872 11056 13266 11112
rect 13322 11056 13327 11112
rect 10872 11054 13327 11056
rect 5533 11051 5599 11054
rect 10685 11051 10751 11054
rect 13261 11051 13327 11054
rect 4981 10978 5047 10981
rect 7097 10978 7163 10981
rect 8017 10978 8083 10981
rect 4981 10976 8083 10978
rect 4981 10920 4986 10976
rect 5042 10920 7102 10976
rect 7158 10920 8022 10976
rect 8078 10920 8083 10976
rect 4981 10918 8083 10920
rect 4981 10915 5047 10918
rect 7097 10915 7163 10918
rect 8017 10915 8083 10918
rect 8845 10978 8911 10981
rect 9765 10980 9831 10981
rect 9438 10978 9444 10980
rect 8845 10976 9444 10978
rect 8845 10920 8850 10976
rect 8906 10920 9444 10976
rect 8845 10918 9444 10920
rect 8845 10915 8911 10918
rect 9438 10916 9444 10918
rect 9508 10916 9514 10980
rect 9765 10976 9812 10980
rect 9876 10978 9882 10980
rect 10593 10978 10659 10981
rect 12801 10978 12867 10981
rect 9765 10920 9770 10976
rect 9765 10916 9812 10920
rect 9876 10918 9922 10978
rect 10593 10976 10978 10978
rect 10593 10920 10598 10976
rect 10654 10920 10978 10976
rect 10593 10918 10978 10920
rect 9876 10916 9882 10918
rect 9765 10915 9831 10916
rect 10593 10915 10659 10918
rect 8340 10912 8660 10913
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 10847 8660 10848
rect 6821 10842 6887 10845
rect 3926 10840 6887 10842
rect 3926 10784 6826 10840
rect 6882 10784 6887 10840
rect 3926 10782 6887 10784
rect 6821 10779 6887 10782
rect 7598 10780 7604 10844
rect 7668 10842 7674 10844
rect 8109 10842 8175 10845
rect 9305 10844 9371 10845
rect 7668 10840 8175 10842
rect 7668 10784 8114 10840
rect 8170 10784 8175 10840
rect 7668 10782 8175 10784
rect 7668 10780 7674 10782
rect 8109 10779 8175 10782
rect 9254 10780 9260 10844
rect 9324 10842 9371 10844
rect 9581 10842 9647 10845
rect 9990 10842 9996 10844
rect 9324 10840 9416 10842
rect 9366 10784 9416 10840
rect 9324 10782 9416 10784
rect 9581 10840 9996 10842
rect 9581 10784 9586 10840
rect 9642 10784 9996 10840
rect 9581 10782 9996 10784
rect 9324 10780 9371 10782
rect 9305 10779 9371 10780
rect 9581 10779 9647 10782
rect 9990 10780 9996 10782
rect 10060 10780 10066 10844
rect 10918 10842 10978 10918
rect 11608 10976 12867 10978
rect 11608 10920 12806 10976
rect 12862 10920 12867 10976
rect 11608 10918 12867 10920
rect 11608 10842 11668 10918
rect 12801 10915 12867 10918
rect 13270 10912 13590 10913
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 10847 13590 10848
rect 10918 10782 11668 10842
rect 11973 10842 12039 10845
rect 12382 10842 12388 10844
rect 11973 10840 12388 10842
rect 11973 10784 11978 10840
rect 12034 10784 12388 10840
rect 11973 10782 12388 10784
rect 11973 10779 12039 10782
rect 12382 10780 12388 10782
rect 12452 10780 12458 10844
rect 3325 10706 3391 10709
rect 3052 10704 3391 10706
rect 3052 10648 3330 10704
rect 3386 10648 3391 10704
rect 3052 10646 3391 10648
rect 3325 10643 3391 10646
rect 3601 10706 3667 10709
rect 9673 10706 9739 10709
rect 12433 10706 12499 10709
rect 3601 10704 9739 10706
rect 3601 10648 3606 10704
rect 3662 10648 9678 10704
rect 9734 10648 9739 10704
rect 3601 10646 9739 10648
rect 3601 10643 3667 10646
rect 9673 10643 9739 10646
rect 9814 10704 12499 10706
rect 9814 10648 12438 10704
rect 12494 10648 12499 10704
rect 9814 10646 12499 10648
rect 2865 10570 2931 10573
rect 4061 10570 4127 10573
rect 6545 10570 6611 10573
rect 2865 10568 6611 10570
rect 2865 10512 2870 10568
rect 2926 10512 4066 10568
rect 4122 10512 6550 10568
rect 6606 10512 6611 10568
rect 2865 10510 6611 10512
rect 2865 10507 2931 10510
rect 4061 10507 4127 10510
rect 6545 10507 6611 10510
rect 6821 10570 6887 10573
rect 9814 10570 9874 10646
rect 12433 10643 12499 10646
rect 10409 10572 10475 10573
rect 6821 10568 9874 10570
rect 6821 10512 6826 10568
rect 6882 10512 9874 10568
rect 6821 10510 9874 10512
rect 6821 10507 6887 10510
rect 10358 10508 10364 10572
rect 10428 10570 10475 10572
rect 11513 10570 11579 10573
rect 14733 10570 14799 10573
rect 10428 10568 10520 10570
rect 10470 10512 10520 10568
rect 10428 10510 10520 10512
rect 10596 10510 11300 10570
rect 10428 10508 10475 10510
rect 10409 10507 10475 10508
rect 6453 10436 6519 10437
rect 6453 10434 6500 10436
rect 6408 10432 6500 10434
rect 6408 10376 6458 10432
rect 6408 10374 6500 10376
rect 6453 10372 6500 10374
rect 6564 10372 6570 10436
rect 6678 10372 6684 10436
rect 6748 10434 6754 10436
rect 7373 10434 7439 10437
rect 6748 10432 7439 10434
rect 6748 10376 7378 10432
rect 7434 10376 7439 10432
rect 6748 10374 7439 10376
rect 6748 10372 6754 10374
rect 6453 10371 6519 10372
rect 7373 10371 7439 10374
rect 7782 10372 7788 10436
rect 7852 10434 7858 10436
rect 10596 10434 10656 10510
rect 7852 10374 10656 10434
rect 7852 10372 7858 10374
rect 5874 10368 6194 10369
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6194 10368
rect 5874 10303 6194 10304
rect 10805 10368 11125 10369
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 10303 11125 10304
rect 4797 10298 4863 10301
rect 5206 10298 5212 10300
rect 4797 10296 5212 10298
rect 4797 10240 4802 10296
rect 4858 10240 5212 10296
rect 4797 10238 5212 10240
rect 4797 10235 4863 10238
rect 5206 10236 5212 10238
rect 5276 10236 5282 10300
rect 7230 10298 7236 10300
rect 6318 10238 7236 10298
rect 4337 10162 4403 10165
rect 6318 10162 6378 10238
rect 7230 10236 7236 10238
rect 7300 10236 7306 10300
rect 7414 10236 7420 10300
rect 7484 10298 7490 10300
rect 10593 10298 10659 10301
rect 7484 10296 10659 10298
rect 7484 10240 10598 10296
rect 10654 10240 10659 10296
rect 7484 10238 10659 10240
rect 11240 10298 11300 10510
rect 11513 10568 14799 10570
rect 11513 10512 11518 10568
rect 11574 10512 14738 10568
rect 14794 10512 14799 10568
rect 11513 10510 14799 10512
rect 11513 10507 11579 10510
rect 14733 10507 14799 10510
rect 11421 10434 11487 10437
rect 11830 10434 11836 10436
rect 11421 10432 11836 10434
rect 11421 10376 11426 10432
rect 11482 10376 11836 10432
rect 11421 10374 11836 10376
rect 11421 10371 11487 10374
rect 11830 10372 11836 10374
rect 11900 10372 11906 10436
rect 13169 10434 13235 10437
rect 13854 10434 13860 10436
rect 13169 10432 13860 10434
rect 13169 10376 13174 10432
rect 13230 10376 13860 10432
rect 13169 10374 13860 10376
rect 13169 10371 13235 10374
rect 13854 10372 13860 10374
rect 13924 10372 13930 10436
rect 13077 10298 13143 10301
rect 11240 10296 13143 10298
rect 11240 10240 13082 10296
rect 13138 10240 13143 10296
rect 11240 10238 13143 10240
rect 7484 10236 7490 10238
rect 10593 10235 10659 10238
rect 13077 10235 13143 10238
rect 4337 10160 6378 10162
rect 4337 10104 4342 10160
rect 4398 10104 6378 10160
rect 4337 10102 6378 10104
rect 4337 10099 4403 10102
rect 7046 10100 7052 10164
rect 7116 10162 7122 10164
rect 10409 10162 10475 10165
rect 7116 10160 10475 10162
rect 7116 10104 10414 10160
rect 10470 10104 10475 10160
rect 7116 10102 10475 10104
rect 7116 10100 7122 10102
rect 10409 10099 10475 10102
rect 10593 10162 10659 10165
rect 13721 10162 13787 10165
rect 10593 10160 13787 10162
rect 10593 10104 10598 10160
rect 10654 10104 13726 10160
rect 13782 10104 13787 10160
rect 10593 10102 13787 10104
rect 10593 10099 10659 10102
rect 13721 10099 13787 10102
rect 6310 10026 6316 10028
rect 3190 9966 6316 10026
rect 0 9890 480 9920
rect 1669 9890 1735 9893
rect 0 9888 1735 9890
rect 0 9832 1674 9888
rect 1730 9832 1735 9888
rect 0 9830 1735 9832
rect 0 9800 480 9830
rect 1669 9827 1735 9830
rect 1853 9890 1919 9893
rect 3190 9890 3250 9966
rect 6310 9964 6316 9966
rect 6380 9964 6386 10028
rect 6862 9964 6868 10028
rect 6932 10026 6938 10028
rect 14641 10026 14707 10029
rect 6932 10024 14707 10026
rect 6932 9968 14646 10024
rect 14702 9968 14707 10024
rect 6932 9966 14707 9968
rect 6932 9964 6938 9966
rect 14641 9963 14707 9966
rect 1853 9888 3250 9890
rect 1853 9832 1858 9888
rect 1914 9832 3250 9888
rect 1853 9830 3250 9832
rect 1853 9827 1919 9830
rect 4838 9828 4844 9892
rect 4908 9890 4914 9892
rect 5206 9890 5212 9892
rect 4908 9830 5212 9890
rect 4908 9828 4914 9830
rect 5206 9828 5212 9830
rect 5276 9828 5282 9892
rect 9990 9828 9996 9892
rect 10060 9890 10066 9892
rect 10542 9890 10548 9892
rect 10060 9830 10548 9890
rect 10060 9828 10066 9830
rect 10542 9828 10548 9830
rect 10612 9828 10618 9892
rect 11973 9890 12039 9893
rect 12750 9890 12756 9892
rect 11973 9888 12756 9890
rect 11973 9832 11978 9888
rect 12034 9832 12756 9888
rect 11973 9830 12756 9832
rect 11973 9827 12039 9830
rect 12750 9828 12756 9830
rect 12820 9828 12826 9892
rect 3409 9824 3729 9825
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 9759 3729 9760
rect 8340 9824 8660 9825
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 9759 8660 9760
rect 13270 9824 13590 9825
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 9759 13590 9760
rect 5165 9754 5231 9757
rect 7649 9754 7715 9757
rect 7833 9754 7899 9757
rect 5165 9752 7899 9754
rect 5165 9696 5170 9752
rect 5226 9696 7654 9752
rect 7710 9696 7838 9752
rect 7894 9696 7899 9752
rect 5165 9694 7899 9696
rect 5165 9691 5231 9694
rect 7649 9691 7715 9694
rect 7833 9691 7899 9694
rect 9070 9692 9076 9756
rect 9140 9754 9146 9756
rect 9765 9754 9831 9757
rect 10133 9756 10199 9757
rect 10133 9754 10180 9756
rect 9140 9752 9831 9754
rect 9140 9696 9770 9752
rect 9826 9696 9831 9752
rect 9140 9694 9831 9696
rect 10088 9752 10180 9754
rect 10088 9696 10138 9752
rect 10088 9694 10180 9696
rect 9140 9692 9146 9694
rect 9765 9691 9831 9694
rect 10133 9692 10180 9694
rect 10244 9692 10250 9756
rect 10317 9754 10383 9757
rect 11646 9754 11652 9756
rect 10317 9752 11652 9754
rect 10317 9696 10322 9752
rect 10378 9696 11652 9752
rect 10317 9694 11652 9696
rect 10133 9691 10199 9692
rect 10317 9691 10383 9694
rect 11646 9692 11652 9694
rect 11716 9692 11722 9756
rect 13905 9754 13971 9757
rect 14038 9754 14044 9756
rect 13905 9752 14044 9754
rect 13905 9696 13910 9752
rect 13966 9696 14044 9752
rect 13905 9694 14044 9696
rect 13905 9691 13971 9694
rect 14038 9692 14044 9694
rect 14108 9692 14114 9756
rect 2773 9618 2839 9621
rect 10409 9618 10475 9621
rect 2773 9616 10475 9618
rect 2773 9560 2778 9616
rect 2834 9560 10414 9616
rect 10470 9560 10475 9616
rect 2773 9558 10475 9560
rect 2773 9555 2839 9558
rect 10409 9555 10475 9558
rect 10542 9556 10548 9620
rect 10612 9618 10618 9620
rect 15009 9618 15075 9621
rect 10612 9616 15075 9618
rect 10612 9560 15014 9616
rect 15070 9560 15075 9616
rect 10612 9558 15075 9560
rect 10612 9556 10618 9558
rect 15009 9555 15075 9558
rect 1945 9482 2011 9485
rect 13629 9482 13695 9485
rect 1945 9480 13695 9482
rect 1945 9424 1950 9480
rect 2006 9424 13634 9480
rect 13690 9424 13695 9480
rect 1945 9422 13695 9424
rect 1945 9419 2011 9422
rect 13629 9419 13695 9422
rect 6678 9284 6684 9348
rect 6748 9346 6754 9348
rect 10542 9346 10548 9348
rect 6748 9286 10548 9346
rect 6748 9284 6754 9286
rect 10542 9284 10548 9286
rect 10612 9284 10618 9348
rect 11329 9346 11395 9349
rect 14273 9346 14339 9349
rect 11329 9344 14339 9346
rect 11329 9288 11334 9344
rect 11390 9288 14278 9344
rect 14334 9288 14339 9344
rect 11329 9286 14339 9288
rect 11329 9283 11395 9286
rect 14273 9283 14339 9286
rect 5874 9280 6194 9281
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6194 9280
rect 5874 9215 6194 9216
rect 10805 9280 11125 9281
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 9215 11125 9216
rect 3601 9210 3667 9213
rect 5073 9210 5139 9213
rect 3601 9208 5139 9210
rect 3601 9152 3606 9208
rect 3662 9152 5078 9208
rect 5134 9152 5139 9208
rect 3601 9150 5139 9152
rect 3601 9147 3667 9150
rect 5073 9147 5139 9150
rect 6310 9148 6316 9212
rect 6380 9210 6386 9212
rect 9213 9210 9279 9213
rect 6380 9208 9279 9210
rect 6380 9152 9218 9208
rect 9274 9152 9279 9208
rect 6380 9150 9279 9152
rect 6380 9148 6386 9150
rect 9213 9147 9279 9150
rect 9622 9148 9628 9212
rect 9692 9210 9698 9212
rect 10542 9210 10548 9212
rect 9692 9150 10548 9210
rect 9692 9148 9698 9150
rect 10542 9148 10548 9150
rect 10612 9148 10618 9212
rect 11646 9148 11652 9212
rect 11716 9210 11722 9212
rect 11973 9210 12039 9213
rect 12157 9212 12223 9213
rect 12433 9212 12499 9213
rect 12157 9210 12204 9212
rect 11716 9208 12039 9210
rect 11716 9152 11978 9208
rect 12034 9152 12039 9208
rect 11716 9150 12039 9152
rect 12112 9208 12204 9210
rect 12112 9152 12162 9208
rect 12112 9150 12204 9152
rect 11716 9148 11722 9150
rect 11973 9147 12039 9150
rect 12157 9148 12204 9150
rect 12268 9148 12274 9212
rect 12382 9148 12388 9212
rect 12452 9210 12499 9212
rect 12452 9208 12544 9210
rect 12494 9152 12544 9208
rect 12452 9150 12544 9152
rect 12985 9208 13051 9213
rect 12985 9152 12990 9208
rect 13046 9152 13051 9208
rect 12452 9148 12499 9150
rect 12157 9147 12223 9148
rect 12433 9147 12499 9148
rect 12985 9147 13051 9152
rect 1577 9074 1643 9077
rect 12525 9074 12591 9077
rect 1577 9072 12591 9074
rect 1577 9016 1582 9072
rect 1638 9016 12530 9072
rect 12586 9016 12591 9072
rect 1577 9014 12591 9016
rect 1577 9011 1643 9014
rect 12525 9011 12591 9014
rect 0 8938 480 8968
rect 2405 8938 2471 8941
rect 8753 8938 8819 8941
rect 0 8878 1410 8938
rect 0 8848 480 8878
rect 1350 8802 1410 8878
rect 2405 8936 8819 8938
rect 2405 8880 2410 8936
rect 2466 8880 8758 8936
rect 8814 8880 8819 8936
rect 2405 8878 8819 8880
rect 2405 8875 2471 8878
rect 8753 8875 8819 8878
rect 9213 8938 9279 8941
rect 10593 8938 10659 8941
rect 9213 8936 10659 8938
rect 9213 8880 9218 8936
rect 9274 8880 10598 8936
rect 10654 8880 10659 8936
rect 9213 8878 10659 8880
rect 9213 8875 9279 8878
rect 10593 8875 10659 8878
rect 11053 8938 11119 8941
rect 11462 8938 11468 8940
rect 11053 8936 11468 8938
rect 11053 8880 11058 8936
rect 11114 8880 11468 8936
rect 11053 8878 11468 8880
rect 11053 8875 11119 8878
rect 11462 8876 11468 8878
rect 11532 8876 11538 8940
rect 12988 8938 13048 9147
rect 11608 8878 13048 8938
rect 2865 8802 2931 8805
rect 1350 8800 2931 8802
rect 1350 8744 2870 8800
rect 2926 8744 2931 8800
rect 1350 8742 2931 8744
rect 2865 8739 2931 8742
rect 6177 8802 6243 8805
rect 7925 8802 7991 8805
rect 6177 8800 7991 8802
rect 6177 8744 6182 8800
rect 6238 8744 7930 8800
rect 7986 8744 7991 8800
rect 6177 8742 7991 8744
rect 6177 8739 6243 8742
rect 7925 8739 7991 8742
rect 8886 8740 8892 8804
rect 8956 8802 8962 8804
rect 11608 8802 11668 8878
rect 8956 8742 11668 8802
rect 11881 8802 11947 8805
rect 12198 8802 12204 8804
rect 11881 8800 12204 8802
rect 11881 8744 11886 8800
rect 11942 8744 12204 8800
rect 11881 8742 12204 8744
rect 8956 8740 8962 8742
rect 11881 8739 11947 8742
rect 12198 8740 12204 8742
rect 12268 8740 12274 8804
rect 13670 8740 13676 8804
rect 13740 8802 13746 8804
rect 14181 8802 14247 8805
rect 13740 8800 14247 8802
rect 13740 8744 14186 8800
rect 14242 8744 14247 8800
rect 13740 8742 14247 8744
rect 13740 8740 13746 8742
rect 14181 8739 14247 8742
rect 3409 8736 3729 8737
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 8671 3729 8672
rect 8340 8736 8660 8737
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 8671 8660 8672
rect 13270 8736 13590 8737
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 8671 13590 8672
rect 3918 8604 3924 8668
rect 3988 8666 3994 8668
rect 7465 8666 7531 8669
rect 7598 8666 7604 8668
rect 3988 8606 7344 8666
rect 3988 8604 3994 8606
rect 2313 8530 2379 8533
rect 6310 8530 6316 8532
rect 2313 8528 6316 8530
rect 2313 8472 2318 8528
rect 2374 8472 6316 8528
rect 2313 8470 6316 8472
rect 2313 8467 2379 8470
rect 6310 8468 6316 8470
rect 6380 8468 6386 8532
rect 6729 8530 6795 8533
rect 6913 8530 6979 8533
rect 6729 8528 6979 8530
rect 6729 8472 6734 8528
rect 6790 8472 6918 8528
rect 6974 8472 6979 8528
rect 6729 8470 6979 8472
rect 7284 8530 7344 8606
rect 7465 8664 7604 8666
rect 7465 8608 7470 8664
rect 7526 8608 7604 8664
rect 7465 8606 7604 8608
rect 7465 8603 7531 8606
rect 7598 8604 7604 8606
rect 7668 8604 7674 8668
rect 8109 8666 8175 8669
rect 13077 8666 13143 8669
rect 7744 8664 8175 8666
rect 7744 8608 8114 8664
rect 8170 8608 8175 8664
rect 7744 8606 8175 8608
rect 7744 8530 7804 8606
rect 8109 8603 8175 8606
rect 8756 8664 13143 8666
rect 8756 8608 13082 8664
rect 13138 8608 13143 8664
rect 8756 8606 13143 8608
rect 7284 8470 7804 8530
rect 8017 8530 8083 8533
rect 8756 8530 8816 8606
rect 13077 8603 13143 8606
rect 12801 8530 12867 8533
rect 8017 8528 8816 8530
rect 8017 8472 8022 8528
rect 8078 8472 8816 8528
rect 8017 8470 8816 8472
rect 8894 8528 12867 8530
rect 8894 8472 12806 8528
rect 12862 8472 12867 8528
rect 8894 8470 12867 8472
rect 6729 8467 6795 8470
rect 6913 8467 6979 8470
rect 8017 8467 8083 8470
rect 3325 8394 3391 8397
rect 8894 8394 8954 8470
rect 12801 8467 12867 8470
rect 11053 8394 11119 8397
rect 3325 8392 8954 8394
rect 3325 8336 3330 8392
rect 3386 8336 8954 8392
rect 3325 8334 8954 8336
rect 9078 8392 11119 8394
rect 9078 8336 11058 8392
rect 11114 8336 11119 8392
rect 9078 8334 11119 8336
rect 3325 8331 3391 8334
rect 2957 8258 3023 8261
rect 4654 8258 4660 8260
rect 2957 8256 4660 8258
rect 2957 8200 2962 8256
rect 3018 8200 4660 8256
rect 2957 8198 4660 8200
rect 2957 8195 3023 8198
rect 4654 8196 4660 8198
rect 4724 8196 4730 8260
rect 5390 8196 5396 8260
rect 5460 8258 5466 8260
rect 5533 8258 5599 8261
rect 5460 8256 5599 8258
rect 5460 8200 5538 8256
rect 5594 8200 5599 8256
rect 5460 8198 5599 8200
rect 5460 8196 5466 8198
rect 5533 8195 5599 8198
rect 7097 8258 7163 8261
rect 9078 8258 9138 8334
rect 11053 8331 11119 8334
rect 11329 8394 11395 8397
rect 13813 8394 13879 8397
rect 11329 8392 13879 8394
rect 11329 8336 11334 8392
rect 11390 8336 13818 8392
rect 13874 8336 13879 8392
rect 11329 8334 13879 8336
rect 11329 8331 11395 8334
rect 13813 8331 13879 8334
rect 9305 8260 9371 8261
rect 7097 8256 9138 8258
rect 7097 8200 7102 8256
rect 7158 8200 9138 8256
rect 7097 8198 9138 8200
rect 7097 8195 7163 8198
rect 9254 8196 9260 8260
rect 9324 8258 9371 8260
rect 9324 8256 9416 8258
rect 9366 8200 9416 8256
rect 9324 8198 9416 8200
rect 9324 8196 9371 8198
rect 9622 8196 9628 8260
rect 9692 8258 9698 8260
rect 9765 8258 9831 8261
rect 9692 8256 9831 8258
rect 9692 8200 9770 8256
rect 9826 8200 9831 8256
rect 9692 8198 9831 8200
rect 9692 8196 9698 8198
rect 9305 8195 9371 8196
rect 9765 8195 9831 8198
rect 11278 8196 11284 8260
rect 11348 8258 11354 8260
rect 11605 8258 11671 8261
rect 11348 8256 11671 8258
rect 11348 8200 11610 8256
rect 11666 8200 11671 8256
rect 11348 8198 11671 8200
rect 11348 8196 11354 8198
rect 11605 8195 11671 8198
rect 12157 8258 12223 8261
rect 14733 8258 14799 8261
rect 12157 8256 14799 8258
rect 12157 8200 12162 8256
rect 12218 8200 14738 8256
rect 14794 8200 14799 8256
rect 12157 8198 14799 8200
rect 12157 8195 12223 8198
rect 14733 8195 14799 8198
rect 5874 8192 6194 8193
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6194 8192
rect 5874 8127 6194 8128
rect 10805 8192 11125 8193
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 8127 11125 8128
rect 3969 8122 4035 8125
rect 1902 8120 4035 8122
rect 1902 8064 3974 8120
rect 4030 8064 4035 8120
rect 1902 8062 4035 8064
rect 0 7850 480 7880
rect 1902 7850 1962 8062
rect 3969 8059 4035 8062
rect 6269 8122 6335 8125
rect 10358 8122 10364 8124
rect 6269 8120 10364 8122
rect 6269 8064 6274 8120
rect 6330 8064 10364 8120
rect 6269 8062 10364 8064
rect 6269 8059 6335 8062
rect 10358 8060 10364 8062
rect 10428 8060 10434 8124
rect 11697 8122 11763 8125
rect 13997 8122 14063 8125
rect 11697 8120 14063 8122
rect 11697 8064 11702 8120
rect 11758 8064 14002 8120
rect 14058 8064 14063 8120
rect 11697 8062 14063 8064
rect 11697 8059 11763 8062
rect 13997 8059 14063 8062
rect 2037 7986 2103 7989
rect 13813 7986 13879 7989
rect 2037 7984 13879 7986
rect 2037 7928 2042 7984
rect 2098 7928 13818 7984
rect 13874 7928 13879 7984
rect 2037 7926 13879 7928
rect 2037 7923 2103 7926
rect 13813 7923 13879 7926
rect 14089 7984 14155 7989
rect 14089 7928 14094 7984
rect 14150 7928 14155 7984
rect 14089 7923 14155 7928
rect 0 7790 1962 7850
rect 2497 7850 2563 7853
rect 5441 7850 5507 7853
rect 11605 7850 11671 7853
rect 2497 7848 5320 7850
rect 2497 7792 2502 7848
rect 2558 7792 5320 7848
rect 2497 7790 5320 7792
rect 0 7760 480 7790
rect 2497 7787 2563 7790
rect 4838 7652 4844 7716
rect 4908 7714 4914 7716
rect 4981 7714 5047 7717
rect 4908 7712 5047 7714
rect 4908 7656 4986 7712
rect 5042 7656 5047 7712
rect 4908 7654 5047 7656
rect 5260 7714 5320 7790
rect 5441 7848 11671 7850
rect 5441 7792 5446 7848
rect 5502 7792 11610 7848
rect 11666 7792 11671 7848
rect 5441 7790 11671 7792
rect 5441 7787 5507 7790
rect 11605 7787 11671 7790
rect 11830 7788 11836 7852
rect 11900 7850 11906 7852
rect 11973 7850 12039 7853
rect 11900 7848 12039 7850
rect 11900 7792 11978 7848
rect 12034 7792 12039 7848
rect 11900 7790 12039 7792
rect 11900 7788 11906 7790
rect 11973 7787 12039 7790
rect 12341 7850 12407 7853
rect 12934 7850 12940 7852
rect 12341 7848 12940 7850
rect 12341 7792 12346 7848
rect 12402 7792 12940 7848
rect 12341 7790 12940 7792
rect 12341 7787 12407 7790
rect 12934 7788 12940 7790
rect 13004 7788 13010 7852
rect 14092 7850 14152 7923
rect 13080 7790 14152 7850
rect 6494 7714 6500 7716
rect 5260 7654 6500 7714
rect 4908 7652 4914 7654
rect 4981 7651 5047 7654
rect 6494 7652 6500 7654
rect 6564 7652 6570 7716
rect 7465 7714 7531 7717
rect 8017 7714 8083 7717
rect 7465 7712 8083 7714
rect 7465 7656 7470 7712
rect 7526 7656 8022 7712
rect 8078 7656 8083 7712
rect 7465 7654 8083 7656
rect 7465 7651 7531 7654
rect 8017 7651 8083 7654
rect 8201 7712 8267 7717
rect 8201 7656 8206 7712
rect 8262 7656 8267 7712
rect 8201 7651 8267 7656
rect 9029 7714 9095 7717
rect 13080 7714 13140 7790
rect 9029 7712 13140 7714
rect 9029 7656 9034 7712
rect 9090 7656 13140 7712
rect 9029 7654 13140 7656
rect 9029 7651 9095 7654
rect 3409 7648 3729 7649
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 7583 3729 7584
rect 4061 7578 4127 7581
rect 6269 7578 6335 7581
rect 8204 7578 8264 7651
rect 8340 7648 8660 7649
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 7583 8660 7584
rect 13270 7648 13590 7649
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 7583 13590 7584
rect 4061 7576 8264 7578
rect 4061 7520 4066 7576
rect 4122 7520 6274 7576
rect 6330 7520 8264 7576
rect 4061 7518 8264 7520
rect 8937 7578 9003 7581
rect 9070 7578 9076 7580
rect 8937 7576 9076 7578
rect 8937 7520 8942 7576
rect 8998 7520 9076 7576
rect 8937 7518 9076 7520
rect 4061 7515 4127 7518
rect 6269 7515 6335 7518
rect 8937 7515 9003 7518
rect 9070 7516 9076 7518
rect 9140 7516 9146 7580
rect 9438 7516 9444 7580
rect 9508 7578 9514 7580
rect 9508 7518 12404 7578
rect 9508 7516 9514 7518
rect 2773 7442 2839 7445
rect 11053 7442 11119 7445
rect 2773 7440 11119 7442
rect 2773 7384 2778 7440
rect 2834 7384 11058 7440
rect 11114 7384 11119 7440
rect 2773 7382 11119 7384
rect 12344 7442 12404 7518
rect 13261 7442 13327 7445
rect 12344 7440 13327 7442
rect 12344 7384 13266 7440
rect 13322 7384 13327 7440
rect 12344 7382 13327 7384
rect 2773 7379 2839 7382
rect 11053 7379 11119 7382
rect 13261 7379 13327 7382
rect 4521 7306 4587 7309
rect 10225 7306 10291 7309
rect 11605 7306 11671 7309
rect 13261 7306 13327 7309
rect 4521 7304 10291 7306
rect 4521 7248 4526 7304
rect 4582 7248 10230 7304
rect 10286 7248 10291 7304
rect 4521 7246 10291 7248
rect 4521 7243 4587 7246
rect 10225 7243 10291 7246
rect 10596 7246 11530 7306
rect 4337 7170 4403 7173
rect 5441 7170 5507 7173
rect 4337 7168 5507 7170
rect 4337 7112 4342 7168
rect 4398 7112 5446 7168
rect 5502 7112 5507 7168
rect 4337 7110 5507 7112
rect 4337 7107 4403 7110
rect 5441 7107 5507 7110
rect 6494 7108 6500 7172
rect 6564 7170 6570 7172
rect 7925 7170 7991 7173
rect 8385 7170 8451 7173
rect 6564 7168 8451 7170
rect 6564 7112 7930 7168
rect 7986 7112 8390 7168
rect 8446 7112 8451 7168
rect 6564 7110 8451 7112
rect 6564 7108 6570 7110
rect 7925 7107 7991 7110
rect 8385 7107 8451 7110
rect 8661 7170 8727 7173
rect 9581 7170 9647 7173
rect 10596 7170 10656 7246
rect 8661 7168 10656 7170
rect 8661 7112 8666 7168
rect 8722 7112 9586 7168
rect 9642 7112 10656 7168
rect 8661 7110 10656 7112
rect 8661 7107 8727 7110
rect 9581 7107 9647 7110
rect 5874 7104 6194 7105
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6194 7104
rect 5874 7039 6194 7040
rect 10805 7104 11125 7105
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 7039 11125 7040
rect 4286 6972 4292 7036
rect 4356 7034 4362 7036
rect 4429 7034 4495 7037
rect 5717 7034 5783 7037
rect 9581 7034 9647 7037
rect 9857 7036 9923 7037
rect 9806 7034 9812 7036
rect 4356 7032 5783 7034
rect 4356 6976 4434 7032
rect 4490 6976 5722 7032
rect 5778 6976 5783 7032
rect 4356 6974 5783 6976
rect 4356 6972 4362 6974
rect 4429 6971 4495 6974
rect 5717 6971 5783 6974
rect 6272 7032 9647 7034
rect 6272 6976 9586 7032
rect 9642 6976 9647 7032
rect 6272 6974 9647 6976
rect 9766 6974 9812 7034
rect 9876 7032 9923 7036
rect 9918 6976 9923 7032
rect 1393 6898 1459 6901
rect 4153 6898 4219 6901
rect 6272 6898 6332 6974
rect 9581 6971 9647 6974
rect 9806 6972 9812 6974
rect 9876 6972 9923 6976
rect 11470 7034 11530 7246
rect 11605 7304 13327 7306
rect 11605 7248 11610 7304
rect 11666 7248 13266 7304
rect 13322 7248 13327 7304
rect 11605 7246 13327 7248
rect 11605 7243 11671 7246
rect 13261 7243 13327 7246
rect 12157 7170 12223 7173
rect 13169 7170 13235 7173
rect 12157 7168 13235 7170
rect 12157 7112 12162 7168
rect 12218 7112 13174 7168
rect 13230 7112 13235 7168
rect 12157 7110 13235 7112
rect 12157 7107 12223 7110
rect 13169 7107 13235 7110
rect 13353 7034 13419 7037
rect 11470 7032 13419 7034
rect 11470 6976 13358 7032
rect 13414 6976 13419 7032
rect 11470 6974 13419 6976
rect 9857 6971 9923 6972
rect 13353 6971 13419 6974
rect 1393 6896 4219 6898
rect 1393 6840 1398 6896
rect 1454 6840 4158 6896
rect 4214 6840 4219 6896
rect 1393 6838 4219 6840
rect 1393 6835 1459 6838
rect 4153 6835 4219 6838
rect 4294 6838 6332 6898
rect 0 6762 480 6792
rect 4294 6762 4354 6838
rect 7230 6836 7236 6900
rect 7300 6898 7306 6900
rect 9070 6898 9076 6900
rect 7300 6838 9076 6898
rect 7300 6836 7306 6838
rect 9070 6836 9076 6838
rect 9140 6836 9146 6900
rect 9397 6898 9463 6901
rect 16757 6898 16823 6901
rect 9397 6896 16823 6898
rect 9397 6840 9402 6896
rect 9458 6840 16762 6896
rect 16818 6840 16823 6896
rect 9397 6838 16823 6840
rect 9397 6835 9463 6838
rect 16757 6835 16823 6838
rect 0 6702 4354 6762
rect 4429 6762 4495 6765
rect 8293 6762 8359 6765
rect 4429 6760 8359 6762
rect 4429 6704 4434 6760
rect 4490 6704 8298 6760
rect 8354 6704 8359 6760
rect 4429 6702 8359 6704
rect 0 6672 480 6702
rect 4429 6699 4495 6702
rect 8293 6699 8359 6702
rect 8477 6762 8543 6765
rect 10041 6762 10107 6765
rect 14457 6762 14523 6765
rect 8477 6760 10107 6762
rect 8477 6704 8482 6760
rect 8538 6704 10046 6760
rect 10102 6704 10107 6760
rect 8477 6702 10107 6704
rect 8477 6699 8543 6702
rect 10041 6699 10107 6702
rect 10182 6760 14523 6762
rect 10182 6704 14462 6760
rect 14518 6704 14523 6760
rect 10182 6702 14523 6704
rect 4153 6626 4219 6629
rect 9949 6626 10015 6629
rect 10182 6626 10242 6702
rect 14457 6699 14523 6702
rect 4153 6624 7482 6626
rect 4153 6568 4158 6624
rect 4214 6568 7482 6624
rect 4153 6566 7482 6568
rect 4153 6563 4219 6566
rect 3409 6560 3729 6561
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 1853 6490 1919 6493
rect 4153 6490 4219 6493
rect 5257 6490 5323 6493
rect 7189 6490 7255 6493
rect 1853 6488 2698 6490
rect 1853 6432 1858 6488
rect 1914 6432 2698 6488
rect 1853 6430 2698 6432
rect 1853 6427 1919 6430
rect 2638 6354 2698 6430
rect 4153 6488 5323 6490
rect 4153 6432 4158 6488
rect 4214 6432 5262 6488
rect 5318 6432 5323 6488
rect 4153 6430 5323 6432
rect 4153 6427 4219 6430
rect 5257 6427 5323 6430
rect 5398 6488 7255 6490
rect 5398 6432 7194 6488
rect 7250 6432 7255 6488
rect 5398 6430 7255 6432
rect 7422 6490 7482 6566
rect 9949 6624 10242 6626
rect 9949 6568 9954 6624
rect 10010 6568 10242 6624
rect 9949 6566 10242 6568
rect 9949 6563 10015 6566
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 8201 6490 8267 6493
rect 7422 6488 8267 6490
rect 7422 6432 8206 6488
rect 8262 6432 8267 6488
rect 7422 6430 8267 6432
rect 4705 6354 4771 6357
rect 2638 6352 4771 6354
rect 2638 6296 4710 6352
rect 4766 6296 4771 6352
rect 2638 6294 4771 6296
rect 4705 6291 4771 6294
rect 4981 6354 5047 6357
rect 5398 6354 5458 6430
rect 7189 6427 7255 6430
rect 8201 6427 8267 6430
rect 8937 6490 9003 6493
rect 9397 6490 9463 6493
rect 10593 6492 10659 6493
rect 8937 6488 9463 6490
rect 8937 6432 8942 6488
rect 8998 6432 9402 6488
rect 9458 6432 9463 6488
rect 8937 6430 9463 6432
rect 8937 6427 9003 6430
rect 9397 6427 9463 6430
rect 10542 6428 10548 6492
rect 10612 6490 10659 6492
rect 10612 6488 10704 6490
rect 10654 6432 10704 6488
rect 10612 6430 10704 6432
rect 10612 6428 10659 6430
rect 10593 6427 10659 6428
rect 4981 6352 5458 6354
rect 4981 6296 4986 6352
rect 5042 6296 5458 6352
rect 4981 6294 5458 6296
rect 6729 6354 6795 6357
rect 15009 6354 15075 6357
rect 6729 6352 15075 6354
rect 6729 6296 6734 6352
rect 6790 6296 15014 6352
rect 15070 6296 15075 6352
rect 6729 6294 15075 6296
rect 4981 6291 5047 6294
rect 6729 6291 6795 6294
rect 15009 6291 15075 6294
rect 4061 6218 4127 6221
rect 11830 6218 11836 6220
rect 4061 6216 11836 6218
rect 4061 6160 4066 6216
rect 4122 6160 11836 6216
rect 4061 6158 11836 6160
rect 4061 6155 4127 6158
rect 11830 6156 11836 6158
rect 11900 6156 11906 6220
rect 4153 6082 4219 6085
rect 5441 6082 5507 6085
rect 4153 6080 5507 6082
rect 4153 6024 4158 6080
rect 4214 6024 5446 6080
rect 5502 6024 5507 6080
rect 4153 6022 5507 6024
rect 4153 6019 4219 6022
rect 5441 6019 5507 6022
rect 6310 6020 6316 6084
rect 6380 6082 6386 6084
rect 7281 6082 7347 6085
rect 6380 6080 7347 6082
rect 6380 6024 7286 6080
rect 7342 6024 7347 6080
rect 6380 6022 7347 6024
rect 6380 6020 6386 6022
rect 7281 6019 7347 6022
rect 7833 6082 7899 6085
rect 8201 6082 8267 6085
rect 7833 6080 8267 6082
rect 7833 6024 7838 6080
rect 7894 6024 8206 6080
rect 8262 6024 8267 6080
rect 7833 6022 8267 6024
rect 7833 6019 7899 6022
rect 8201 6019 8267 6022
rect 8569 6082 8635 6085
rect 8937 6082 9003 6085
rect 8569 6080 9003 6082
rect 8569 6024 8574 6080
rect 8630 6024 8942 6080
rect 8998 6024 9003 6080
rect 8569 6022 9003 6024
rect 8569 6019 8635 6022
rect 8937 6019 9003 6022
rect 9070 6020 9076 6084
rect 9140 6082 9146 6084
rect 10174 6082 10180 6084
rect 9140 6022 10180 6082
rect 9140 6020 9146 6022
rect 10174 6020 10180 6022
rect 10244 6082 10250 6084
rect 10501 6082 10567 6085
rect 10244 6080 10567 6082
rect 10244 6024 10506 6080
rect 10562 6024 10567 6080
rect 10244 6022 10567 6024
rect 10244 6020 10250 6022
rect 10501 6019 10567 6022
rect 11237 6082 11303 6085
rect 11462 6082 11468 6084
rect 11237 6080 11468 6082
rect 11237 6024 11242 6080
rect 11298 6024 11468 6080
rect 11237 6022 11468 6024
rect 11237 6019 11303 6022
rect 11462 6020 11468 6022
rect 11532 6020 11538 6084
rect 12433 6082 12499 6085
rect 12801 6082 12867 6085
rect 12433 6080 12867 6082
rect 12433 6024 12438 6080
rect 12494 6024 12806 6080
rect 12862 6024 12867 6080
rect 12433 6022 12867 6024
rect 12433 6019 12499 6022
rect 12801 6019 12867 6022
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 5022 5946 5028 5948
rect 2638 5886 5028 5946
rect 2638 5813 2698 5886
rect 5022 5884 5028 5886
rect 5092 5884 5098 5948
rect 6494 5884 6500 5948
rect 6564 5946 6570 5948
rect 9806 5946 9812 5948
rect 6564 5886 9812 5946
rect 6564 5884 6570 5886
rect 9806 5884 9812 5886
rect 9876 5884 9882 5948
rect 10041 5946 10107 5949
rect 10225 5946 10291 5949
rect 10041 5944 10291 5946
rect 10041 5888 10046 5944
rect 10102 5888 10230 5944
rect 10286 5888 10291 5944
rect 10041 5886 10291 5888
rect 10041 5883 10107 5886
rect 10225 5883 10291 5886
rect 2589 5808 2698 5813
rect 2589 5752 2594 5808
rect 2650 5752 2698 5808
rect 2589 5750 2698 5752
rect 2773 5810 2839 5813
rect 9305 5810 9371 5813
rect 2773 5808 9371 5810
rect 2773 5752 2778 5808
rect 2834 5752 9310 5808
rect 9366 5752 9371 5808
rect 2773 5750 9371 5752
rect 2589 5747 2655 5750
rect 2773 5747 2839 5750
rect 9305 5747 9371 5750
rect 10041 5810 10107 5813
rect 12566 5810 12572 5812
rect 10041 5808 12572 5810
rect 10041 5752 10046 5808
rect 10102 5752 12572 5808
rect 10041 5750 12572 5752
rect 10041 5747 10107 5750
rect 12566 5748 12572 5750
rect 12636 5748 12642 5812
rect 0 5674 480 5704
rect 3877 5674 3943 5677
rect 0 5672 3943 5674
rect 0 5616 3882 5672
rect 3938 5616 3943 5672
rect 0 5614 3943 5616
rect 0 5584 480 5614
rect 3877 5611 3943 5614
rect 4705 5674 4771 5677
rect 10501 5674 10567 5677
rect 4705 5672 10567 5674
rect 4705 5616 4710 5672
rect 4766 5616 10506 5672
rect 10562 5616 10567 5672
rect 4705 5614 10567 5616
rect 4705 5611 4771 5614
rect 10501 5611 10567 5614
rect 11053 5674 11119 5677
rect 12341 5674 12407 5677
rect 11053 5672 12407 5674
rect 11053 5616 11058 5672
rect 11114 5616 12346 5672
rect 12402 5616 12407 5672
rect 11053 5614 12407 5616
rect 11053 5611 11119 5614
rect 12341 5611 12407 5614
rect 4061 5538 4127 5541
rect 7230 5538 7236 5540
rect 4061 5536 7236 5538
rect 4061 5480 4066 5536
rect 4122 5480 7236 5536
rect 4061 5478 7236 5480
rect 4061 5475 4127 5478
rect 7230 5476 7236 5478
rect 7300 5476 7306 5540
rect 9765 5538 9831 5541
rect 12382 5538 12388 5540
rect 9765 5536 12388 5538
rect 9765 5480 9770 5536
rect 9826 5480 12388 5536
rect 9765 5478 12388 5480
rect 9765 5475 9831 5478
rect 12382 5476 12388 5478
rect 12452 5538 12458 5540
rect 12709 5538 12775 5541
rect 12452 5536 12775 5538
rect 12452 5480 12714 5536
rect 12770 5480 12775 5536
rect 12452 5478 12775 5480
rect 12452 5476 12458 5478
rect 12709 5475 12775 5478
rect 3409 5472 3729 5473
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 4613 5402 4679 5405
rect 7281 5402 7347 5405
rect 8109 5402 8175 5405
rect 4613 5400 6010 5402
rect 4613 5344 4618 5400
rect 4674 5344 6010 5400
rect 4613 5342 6010 5344
rect 4613 5339 4679 5342
rect 1853 5266 1919 5269
rect 5809 5266 5875 5269
rect 1853 5264 5875 5266
rect 1853 5208 1858 5264
rect 1914 5208 5814 5264
rect 5870 5208 5875 5264
rect 1853 5206 5875 5208
rect 5950 5266 6010 5342
rect 7281 5400 8175 5402
rect 7281 5344 7286 5400
rect 7342 5344 8114 5400
rect 8170 5344 8175 5400
rect 7281 5342 8175 5344
rect 7281 5339 7347 5342
rect 8109 5339 8175 5342
rect 9305 5402 9371 5405
rect 9673 5402 9739 5405
rect 9305 5400 9739 5402
rect 9305 5344 9310 5400
rect 9366 5344 9678 5400
rect 9734 5344 9739 5400
rect 9305 5342 9739 5344
rect 9305 5339 9371 5342
rect 9673 5339 9739 5342
rect 9949 5402 10015 5405
rect 10869 5402 10935 5405
rect 9949 5400 10935 5402
rect 9949 5344 9954 5400
rect 10010 5344 10874 5400
rect 10930 5344 10935 5400
rect 9949 5342 10935 5344
rect 9949 5339 10015 5342
rect 10869 5339 10935 5342
rect 11145 5402 11211 5405
rect 11421 5402 11487 5405
rect 11145 5400 11487 5402
rect 11145 5344 11150 5400
rect 11206 5344 11426 5400
rect 11482 5344 11487 5400
rect 11145 5342 11487 5344
rect 11145 5339 11211 5342
rect 11421 5339 11487 5342
rect 12249 5402 12315 5405
rect 12566 5402 12572 5404
rect 12249 5400 12572 5402
rect 12249 5344 12254 5400
rect 12310 5344 12572 5400
rect 12249 5342 12572 5344
rect 12249 5339 12315 5342
rect 12566 5340 12572 5342
rect 12636 5340 12642 5404
rect 14089 5266 14155 5269
rect 5950 5264 14155 5266
rect 5950 5208 14094 5264
rect 14150 5208 14155 5264
rect 5950 5206 14155 5208
rect 1853 5203 1919 5206
rect 5809 5203 5875 5206
rect 14089 5203 14155 5206
rect 4061 5128 4127 5133
rect 4061 5072 4066 5128
rect 4122 5072 4127 5128
rect 4061 5067 4127 5072
rect 5349 5130 5415 5133
rect 7005 5130 7071 5133
rect 5349 5128 7071 5130
rect 5349 5072 5354 5128
rect 5410 5072 7010 5128
rect 7066 5072 7071 5128
rect 5349 5070 7071 5072
rect 5349 5067 5415 5070
rect 7005 5067 7071 5070
rect 7230 5068 7236 5132
rect 7300 5130 7306 5132
rect 9765 5130 9831 5133
rect 7300 5128 9831 5130
rect 7300 5072 9770 5128
rect 9826 5072 9831 5128
rect 7300 5070 9831 5072
rect 7300 5068 7306 5070
rect 9765 5067 9831 5070
rect 9998 5070 14474 5130
rect 2681 4858 2747 4861
rect 4064 4858 4124 5067
rect 6637 4994 6703 4997
rect 9998 4994 10058 5070
rect 6637 4992 10058 4994
rect 6637 4936 6642 4992
rect 6698 4936 10058 4992
rect 6637 4934 10058 4936
rect 11237 4994 11303 4997
rect 11462 4994 11468 4996
rect 11237 4992 11468 4994
rect 11237 4936 11242 4992
rect 11298 4936 11468 4992
rect 11237 4934 11468 4936
rect 6637 4931 6703 4934
rect 11237 4931 11303 4934
rect 11462 4932 11468 4934
rect 11532 4932 11538 4996
rect 13813 4994 13879 4997
rect 12942 4992 13879 4994
rect 12942 4936 13818 4992
rect 13874 4936 13879 4992
rect 12942 4934 13879 4936
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 2681 4856 4124 4858
rect 2681 4800 2686 4856
rect 2742 4800 4124 4856
rect 2681 4798 4124 4800
rect 4521 4858 4587 4861
rect 5717 4858 5783 4861
rect 4521 4856 5783 4858
rect 4521 4800 4526 4856
rect 4582 4800 5722 4856
rect 5778 4800 5783 4856
rect 4521 4798 5783 4800
rect 2681 4795 2747 4798
rect 4521 4795 4587 4798
rect 5717 4795 5783 4798
rect 7005 4858 7071 4861
rect 8886 4858 8892 4860
rect 7005 4856 8892 4858
rect 7005 4800 7010 4856
rect 7066 4800 8892 4856
rect 7005 4798 8892 4800
rect 7005 4795 7071 4798
rect 8886 4796 8892 4798
rect 8956 4796 8962 4860
rect 9673 4858 9739 4861
rect 10593 4858 10659 4861
rect 9673 4856 10659 4858
rect 9673 4800 9678 4856
rect 9734 4800 10598 4856
rect 10654 4800 10659 4856
rect 9673 4798 10659 4800
rect 9673 4795 9739 4798
rect 10593 4795 10659 4798
rect 11646 4796 11652 4860
rect 11716 4858 11722 4860
rect 11881 4858 11947 4861
rect 11716 4856 11947 4858
rect 11716 4800 11886 4856
rect 11942 4800 11947 4856
rect 11716 4798 11947 4800
rect 11716 4796 11722 4798
rect 11881 4795 11947 4798
rect 12525 4858 12591 4861
rect 12750 4858 12756 4860
rect 12525 4856 12756 4858
rect 12525 4800 12530 4856
rect 12586 4800 12756 4856
rect 12525 4798 12756 4800
rect 12525 4795 12591 4798
rect 12750 4796 12756 4798
rect 12820 4796 12826 4860
rect 0 4722 480 4752
rect 4981 4722 5047 4725
rect 0 4720 5047 4722
rect 0 4664 4986 4720
rect 5042 4664 5047 4720
rect 0 4662 5047 4664
rect 0 4632 480 4662
rect 4981 4659 5047 4662
rect 5809 4722 5875 4725
rect 12942 4722 13002 4934
rect 13813 4931 13879 4934
rect 5809 4720 13002 4722
rect 5809 4664 5814 4720
rect 5870 4664 13002 4720
rect 5809 4662 13002 4664
rect 5809 4659 5875 4662
rect 3877 4586 3943 4589
rect 7005 4586 7071 4589
rect 3877 4584 7071 4586
rect 3877 4528 3882 4584
rect 3938 4528 7010 4584
rect 7066 4528 7071 4584
rect 3877 4526 7071 4528
rect 3877 4523 3943 4526
rect 7005 4523 7071 4526
rect 7373 4586 7439 4589
rect 11421 4586 11487 4589
rect 11881 4588 11947 4589
rect 11830 4586 11836 4588
rect 7373 4584 11487 4586
rect 7373 4528 7378 4584
rect 7434 4528 11426 4584
rect 11482 4528 11487 4584
rect 7373 4526 11487 4528
rect 11790 4526 11836 4586
rect 11900 4584 11947 4588
rect 12382 4586 12388 4588
rect 11942 4528 11947 4584
rect 7373 4523 7439 4526
rect 11421 4523 11487 4526
rect 11830 4524 11836 4526
rect 11900 4524 11947 4528
rect 11881 4523 11947 4524
rect 12160 4526 12388 4586
rect 5809 4450 5875 4453
rect 6862 4450 6868 4452
rect 5809 4448 6868 4450
rect 5809 4392 5814 4448
rect 5870 4392 6868 4448
rect 5809 4390 6868 4392
rect 5809 4387 5875 4390
rect 6862 4388 6868 4390
rect 6932 4388 6938 4452
rect 7189 4450 7255 4453
rect 8109 4450 8175 4453
rect 7189 4448 8175 4450
rect 7189 4392 7194 4448
rect 7250 4392 8114 4448
rect 8170 4392 8175 4448
rect 7189 4390 8175 4392
rect 7189 4387 7255 4390
rect 8109 4387 8175 4390
rect 8937 4450 9003 4453
rect 12160 4450 12220 4526
rect 12382 4524 12388 4526
rect 12452 4586 12458 4588
rect 14181 4586 14247 4589
rect 12452 4584 14247 4586
rect 12452 4528 14186 4584
rect 14242 4528 14247 4584
rect 12452 4526 14247 4528
rect 14414 4586 14474 5070
rect 16520 4586 17000 4616
rect 14414 4526 17000 4586
rect 12452 4524 12458 4526
rect 14181 4523 14247 4526
rect 16520 4496 17000 4526
rect 8937 4448 12220 4450
rect 8937 4392 8942 4448
rect 8998 4392 12220 4448
rect 8937 4390 12220 4392
rect 8937 4387 9003 4390
rect 3409 4384 3729 4385
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 3877 4314 3943 4317
rect 8109 4314 8175 4317
rect 3877 4312 8175 4314
rect 3877 4256 3882 4312
rect 3938 4256 8114 4312
rect 8170 4256 8175 4312
rect 3877 4254 8175 4256
rect 3877 4251 3943 4254
rect 8109 4251 8175 4254
rect 8886 4252 8892 4316
rect 8956 4314 8962 4316
rect 9029 4314 9095 4317
rect 9262 4316 9322 4390
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 4319 13590 4320
rect 8956 4312 9095 4314
rect 8956 4256 9034 4312
rect 9090 4256 9095 4312
rect 8956 4254 9095 4256
rect 8956 4252 8962 4254
rect 9029 4251 9095 4254
rect 9254 4252 9260 4316
rect 9324 4252 9330 4316
rect 9622 4252 9628 4316
rect 9692 4314 9698 4316
rect 10133 4314 10199 4317
rect 9692 4312 10199 4314
rect 9692 4256 10138 4312
rect 10194 4256 10199 4312
rect 9692 4254 10199 4256
rect 9692 4252 9698 4254
rect 10133 4251 10199 4254
rect 11145 4314 11211 4317
rect 11145 4312 13186 4314
rect 11145 4256 11150 4312
rect 11206 4256 13186 4312
rect 11145 4254 13186 4256
rect 11145 4251 11211 4254
rect 6494 4178 6500 4180
rect 5950 4118 6500 4178
rect 3785 4042 3851 4045
rect 5950 4042 6010 4118
rect 6494 4116 6500 4118
rect 6564 4116 6570 4180
rect 6729 4178 6795 4181
rect 12433 4178 12499 4181
rect 6729 4176 12499 4178
rect 6729 4120 6734 4176
rect 6790 4120 12438 4176
rect 12494 4120 12499 4176
rect 6729 4118 12499 4120
rect 13126 4178 13186 4254
rect 14641 4178 14707 4181
rect 13126 4176 14707 4178
rect 13126 4120 14646 4176
rect 14702 4120 14707 4176
rect 13126 4118 14707 4120
rect 6729 4115 6795 4118
rect 12433 4115 12499 4118
rect 14641 4115 14707 4118
rect 14917 4178 14983 4181
rect 15377 4178 15443 4181
rect 14917 4176 15443 4178
rect 14917 4120 14922 4176
rect 14978 4120 15382 4176
rect 15438 4120 15443 4176
rect 14917 4118 15443 4120
rect 14917 4115 14983 4118
rect 15377 4115 15443 4118
rect 3785 4040 6010 4042
rect 3785 3984 3790 4040
rect 3846 3984 6010 4040
rect 3785 3982 6010 3984
rect 6545 4042 6611 4045
rect 12525 4042 12591 4045
rect 14457 4042 14523 4045
rect 6545 4040 11346 4042
rect 6545 3984 6550 4040
rect 6606 3984 11346 4040
rect 6545 3982 11346 3984
rect 3785 3979 3851 3982
rect 6545 3979 6611 3982
rect 2865 3906 2931 3909
rect 2998 3906 3004 3908
rect 2865 3904 3004 3906
rect 2865 3848 2870 3904
rect 2926 3848 3004 3904
rect 2865 3846 3004 3848
rect 2865 3843 2931 3846
rect 2998 3844 3004 3846
rect 3068 3844 3074 3908
rect 6913 3906 6979 3909
rect 10501 3906 10567 3909
rect 6913 3904 10567 3906
rect 6913 3848 6918 3904
rect 6974 3848 10506 3904
rect 10562 3848 10567 3904
rect 6913 3846 10567 3848
rect 6913 3843 6979 3846
rect 10501 3843 10567 3846
rect 5874 3840 6194 3841
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 2037 3770 2103 3773
rect 5625 3772 5691 3773
rect 5574 3770 5580 3772
rect 2037 3768 5580 3770
rect 5644 3770 5691 3772
rect 7189 3770 7255 3773
rect 10409 3770 10475 3773
rect 5644 3768 5736 3770
rect 2037 3712 2042 3768
rect 2098 3712 5580 3768
rect 5686 3712 5736 3768
rect 2037 3710 5580 3712
rect 2037 3707 2103 3710
rect 5574 3708 5580 3710
rect 5644 3710 5736 3712
rect 7189 3768 10475 3770
rect 7189 3712 7194 3768
rect 7250 3712 10414 3768
rect 10470 3712 10475 3768
rect 7189 3710 10475 3712
rect 5644 3708 5691 3710
rect 5625 3707 5691 3708
rect 7189 3707 7255 3710
rect 10409 3707 10475 3710
rect 0 3634 480 3664
rect 3918 3634 3924 3636
rect 0 3574 3924 3634
rect 0 3544 480 3574
rect 3918 3572 3924 3574
rect 3988 3572 3994 3636
rect 4521 3634 4587 3637
rect 11145 3634 11211 3637
rect 4521 3632 11211 3634
rect 4521 3576 4526 3632
rect 4582 3576 11150 3632
rect 11206 3576 11211 3632
rect 4521 3574 11211 3576
rect 11286 3634 11346 3982
rect 12525 4040 14523 4042
rect 12525 3984 12530 4040
rect 12586 3984 14462 4040
rect 14518 3984 14523 4040
rect 12525 3982 14523 3984
rect 12525 3979 12591 3982
rect 14457 3979 14523 3982
rect 11697 3906 11763 3909
rect 13670 3906 13676 3908
rect 11697 3904 13676 3906
rect 11697 3848 11702 3904
rect 11758 3848 13676 3904
rect 11697 3846 13676 3848
rect 11697 3843 11763 3846
rect 13670 3844 13676 3846
rect 13740 3844 13746 3908
rect 11881 3770 11947 3773
rect 13813 3770 13879 3773
rect 11881 3768 13879 3770
rect 11881 3712 11886 3768
rect 11942 3712 13818 3768
rect 13874 3712 13879 3768
rect 11881 3710 13879 3712
rect 11881 3707 11947 3710
rect 13813 3707 13879 3710
rect 13445 3634 13511 3637
rect 11286 3632 13511 3634
rect 11286 3576 13450 3632
rect 13506 3576 13511 3632
rect 11286 3574 13511 3576
rect 4521 3571 4587 3574
rect 11145 3571 11211 3574
rect 13445 3571 13511 3574
rect 565 3498 631 3501
rect 9949 3498 10015 3501
rect 12014 3498 12020 3500
rect 565 3496 10015 3498
rect 565 3440 570 3496
rect 626 3440 9954 3496
rect 10010 3440 10015 3496
rect 565 3438 10015 3440
rect 565 3435 631 3438
rect 9949 3435 10015 3438
rect 10182 3438 12020 3498
rect 4429 3362 4495 3365
rect 5206 3362 5212 3364
rect 4429 3360 5212 3362
rect 4429 3304 4434 3360
rect 4490 3304 5212 3360
rect 4429 3302 5212 3304
rect 4429 3299 4495 3302
rect 5206 3300 5212 3302
rect 5276 3362 5282 3364
rect 6913 3362 6979 3365
rect 7097 3364 7163 3365
rect 5276 3360 6979 3362
rect 5276 3304 6918 3360
rect 6974 3304 6979 3360
rect 5276 3302 6979 3304
rect 5276 3300 5282 3302
rect 6913 3299 6979 3302
rect 7046 3300 7052 3364
rect 7116 3362 7163 3364
rect 7373 3364 7439 3365
rect 7373 3362 7420 3364
rect 7116 3360 7208 3362
rect 7158 3304 7208 3360
rect 7116 3302 7208 3304
rect 7328 3360 7420 3362
rect 7328 3304 7378 3360
rect 7328 3302 7420 3304
rect 7116 3300 7163 3302
rect 7097 3299 7163 3300
rect 7373 3300 7420 3302
rect 7484 3300 7490 3364
rect 9213 3362 9279 3365
rect 10182 3362 10242 3438
rect 12014 3436 12020 3438
rect 12084 3436 12090 3500
rect 12341 3498 12407 3501
rect 13353 3498 13419 3501
rect 13813 3500 13879 3501
rect 13813 3498 13860 3500
rect 12341 3496 13419 3498
rect 12341 3440 12346 3496
rect 12402 3440 13358 3496
rect 13414 3440 13419 3496
rect 12341 3438 13419 3440
rect 13768 3496 13860 3498
rect 13768 3440 13818 3496
rect 13768 3438 13860 3440
rect 12341 3435 12407 3438
rect 13353 3435 13419 3438
rect 13813 3436 13860 3438
rect 13924 3436 13930 3500
rect 13813 3435 13879 3436
rect 9213 3360 10242 3362
rect 9213 3304 9218 3360
rect 9274 3304 10242 3360
rect 9213 3302 10242 3304
rect 7373 3299 7439 3300
rect 9213 3299 9279 3302
rect 10542 3300 10548 3364
rect 10612 3362 10618 3364
rect 11421 3362 11487 3365
rect 13077 3362 13143 3365
rect 10612 3360 13143 3362
rect 10612 3304 11426 3360
rect 11482 3304 13082 3360
rect 13138 3304 13143 3360
rect 10612 3302 13143 3304
rect 10612 3300 10618 3302
rect 11421 3299 11487 3302
rect 13077 3299 13143 3302
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 3231 13590 3232
rect 4797 3226 4863 3229
rect 5257 3226 5323 3229
rect 4797 3224 5323 3226
rect 4797 3168 4802 3224
rect 4858 3168 5262 3224
rect 5318 3168 5323 3224
rect 4797 3166 5323 3168
rect 4797 3163 4863 3166
rect 5257 3163 5323 3166
rect 5533 3226 5599 3229
rect 8201 3226 8267 3229
rect 5533 3224 8267 3226
rect 5533 3168 5538 3224
rect 5594 3168 8206 3224
rect 8262 3168 8267 3224
rect 5533 3166 8267 3168
rect 5533 3163 5599 3166
rect 8201 3163 8267 3166
rect 8886 3164 8892 3228
rect 8956 3226 8962 3228
rect 11789 3226 11855 3229
rect 8956 3224 11855 3226
rect 8956 3168 11794 3224
rect 11850 3168 11855 3224
rect 8956 3166 11855 3168
rect 8956 3164 8962 3166
rect 11789 3163 11855 3166
rect 12198 3164 12204 3228
rect 12268 3226 12274 3228
rect 12709 3226 12775 3229
rect 12268 3224 12775 3226
rect 12268 3168 12714 3224
rect 12770 3168 12775 3224
rect 12268 3166 12775 3168
rect 12268 3164 12274 3166
rect 12709 3163 12775 3166
rect 5165 3090 5231 3093
rect 13721 3090 13787 3093
rect 5165 3088 13787 3090
rect 5165 3032 5170 3088
rect 5226 3032 13726 3088
rect 13782 3032 13787 3088
rect 5165 3030 13787 3032
rect 5165 3027 5231 3030
rect 13721 3027 13787 3030
rect 1025 2954 1091 2957
rect 4521 2954 4587 2957
rect 1025 2952 4587 2954
rect 1025 2896 1030 2952
rect 1086 2896 4526 2952
rect 4582 2896 4587 2952
rect 1025 2894 4587 2896
rect 1025 2891 1091 2894
rect 4521 2891 4587 2894
rect 4797 2954 4863 2957
rect 7046 2954 7052 2956
rect 4797 2952 7052 2954
rect 4797 2896 4802 2952
rect 4858 2896 7052 2952
rect 4797 2894 7052 2896
rect 4797 2891 4863 2894
rect 7046 2892 7052 2894
rect 7116 2892 7122 2956
rect 15009 2954 15075 2957
rect 7192 2952 15075 2954
rect 7192 2896 15014 2952
rect 15070 2896 15075 2952
rect 7192 2894 15075 2896
rect 2773 2818 2839 2821
rect 4429 2818 4495 2821
rect 2773 2816 4495 2818
rect 2773 2760 2778 2816
rect 2834 2760 4434 2816
rect 4490 2760 4495 2816
rect 2773 2758 4495 2760
rect 2773 2755 2839 2758
rect 4429 2755 4495 2758
rect 6729 2818 6795 2821
rect 7192 2818 7252 2894
rect 15009 2891 15075 2894
rect 6729 2816 7252 2818
rect 6729 2760 6734 2816
rect 6790 2760 7252 2816
rect 6729 2758 7252 2760
rect 7833 2818 7899 2821
rect 10041 2820 10107 2821
rect 7966 2818 7972 2820
rect 7833 2816 7972 2818
rect 7833 2760 7838 2816
rect 7894 2760 7972 2816
rect 7833 2758 7972 2760
rect 6729 2755 6795 2758
rect 7833 2755 7899 2758
rect 7966 2756 7972 2758
rect 8036 2756 8042 2820
rect 9990 2818 9996 2820
rect 9914 2758 9996 2818
rect 10060 2818 10107 2820
rect 10225 2818 10291 2821
rect 10060 2816 10291 2818
rect 10102 2760 10230 2816
rect 10286 2760 10291 2816
rect 9990 2756 9996 2758
rect 10060 2758 10291 2760
rect 10060 2756 10107 2758
rect 10041 2755 10107 2756
rect 10225 2755 10291 2758
rect 11789 2818 11855 2821
rect 14549 2818 14615 2821
rect 11789 2816 14615 2818
rect 11789 2760 11794 2816
rect 11850 2760 14554 2816
rect 14610 2760 14615 2816
rect 11789 2758 14615 2760
rect 11789 2755 11855 2758
rect 14549 2755 14615 2758
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 2773 2682 2839 2685
rect 5625 2682 5691 2685
rect 2773 2680 5691 2682
rect 2773 2624 2778 2680
rect 2834 2624 5630 2680
rect 5686 2624 5691 2680
rect 2773 2622 5691 2624
rect 2773 2619 2839 2622
rect 5625 2619 5691 2622
rect 6310 2620 6316 2684
rect 6380 2682 6386 2684
rect 6545 2682 6611 2685
rect 6380 2680 6611 2682
rect 6380 2624 6550 2680
rect 6606 2624 6611 2680
rect 6380 2622 6611 2624
rect 6380 2620 6386 2622
rect 6545 2619 6611 2622
rect 7005 2682 7071 2685
rect 8201 2684 8267 2685
rect 7782 2682 7788 2684
rect 7005 2680 7788 2682
rect 7005 2624 7010 2680
rect 7066 2624 7788 2680
rect 7005 2622 7788 2624
rect 7005 2619 7071 2622
rect 7782 2620 7788 2622
rect 7852 2620 7858 2684
rect 8150 2620 8156 2684
rect 8220 2682 8267 2684
rect 8569 2682 8635 2685
rect 9949 2682 10015 2685
rect 8220 2680 8312 2682
rect 8262 2624 8312 2680
rect 8220 2622 8312 2624
rect 8569 2680 10015 2682
rect 8569 2624 8574 2680
rect 8630 2624 9954 2680
rect 10010 2624 10015 2680
rect 8569 2622 10015 2624
rect 8220 2620 8267 2622
rect 8201 2619 8267 2620
rect 8569 2619 8635 2622
rect 9949 2619 10015 2622
rect 10174 2620 10180 2684
rect 10244 2682 10250 2684
rect 10593 2682 10659 2685
rect 11329 2684 11395 2685
rect 10244 2680 10659 2682
rect 10244 2624 10598 2680
rect 10654 2624 10659 2680
rect 10244 2622 10659 2624
rect 10244 2620 10250 2622
rect 10593 2619 10659 2622
rect 11278 2620 11284 2684
rect 11348 2682 11395 2684
rect 11973 2682 12039 2685
rect 13077 2682 13143 2685
rect 11348 2680 11440 2682
rect 11390 2624 11440 2680
rect 11348 2622 11440 2624
rect 11973 2680 13143 2682
rect 11973 2624 11978 2680
rect 12034 2624 13082 2680
rect 13138 2624 13143 2680
rect 11973 2622 13143 2624
rect 11348 2620 11395 2622
rect 11329 2619 11395 2620
rect 11973 2619 12039 2622
rect 13077 2619 13143 2622
rect 0 2546 480 2576
rect 4061 2546 4127 2549
rect 0 2544 4127 2546
rect 0 2488 4066 2544
rect 4122 2488 4127 2544
rect 0 2486 4127 2488
rect 0 2456 480 2486
rect 4061 2483 4127 2486
rect 5257 2546 5323 2549
rect 6678 2546 6684 2548
rect 5257 2544 6684 2546
rect 5257 2488 5262 2544
rect 5318 2488 6684 2544
rect 5257 2486 6684 2488
rect 5257 2483 5323 2486
rect 6678 2484 6684 2486
rect 6748 2484 6754 2548
rect 7046 2484 7052 2548
rect 7116 2546 7122 2548
rect 8753 2546 8819 2549
rect 13118 2546 13124 2548
rect 7116 2486 8402 2546
rect 7116 2484 7122 2486
rect 4981 2410 5047 2413
rect 7598 2410 7604 2412
rect 4981 2408 7604 2410
rect 4981 2352 4986 2408
rect 5042 2352 7604 2408
rect 4981 2350 7604 2352
rect 4981 2347 5047 2350
rect 7598 2348 7604 2350
rect 7668 2410 7674 2412
rect 7925 2410 7991 2413
rect 7668 2408 7991 2410
rect 7668 2352 7930 2408
rect 7986 2352 7991 2408
rect 7668 2350 7991 2352
rect 8342 2410 8402 2486
rect 8753 2544 13124 2546
rect 8753 2488 8758 2544
rect 8814 2488 13124 2544
rect 8753 2486 13124 2488
rect 8753 2483 8819 2486
rect 13118 2484 13124 2486
rect 13188 2484 13194 2548
rect 11789 2410 11855 2413
rect 8342 2408 11855 2410
rect 8342 2352 11794 2408
rect 11850 2352 11855 2408
rect 8342 2350 11855 2352
rect 7668 2348 7674 2350
rect 7925 2347 7991 2350
rect 11789 2347 11855 2350
rect 12566 2348 12572 2412
rect 12636 2410 12642 2412
rect 13077 2410 13143 2413
rect 12636 2408 13143 2410
rect 12636 2352 13082 2408
rect 13138 2352 13143 2408
rect 12636 2350 13143 2352
rect 12636 2348 12642 2350
rect 13077 2347 13143 2350
rect 5390 2212 5396 2276
rect 5460 2274 5466 2276
rect 7557 2274 7623 2277
rect 5460 2272 7623 2274
rect 5460 2216 7562 2272
rect 7618 2216 7623 2272
rect 5460 2214 7623 2216
rect 5460 2212 5466 2214
rect 7557 2211 7623 2214
rect 9305 2274 9371 2277
rect 13077 2274 13143 2277
rect 9305 2272 13143 2274
rect 9305 2216 9310 2272
rect 9366 2216 13082 2272
rect 13138 2216 13143 2272
rect 9305 2214 13143 2216
rect 9305 2211 9371 2214
rect 13077 2211 13143 2214
rect 3409 2208 3729 2209
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
rect 10358 2076 10364 2140
rect 10428 2138 10434 2140
rect 11237 2138 11303 2141
rect 10428 2136 11303 2138
rect 10428 2080 11242 2136
rect 11298 2080 11303 2136
rect 10428 2078 11303 2080
rect 10428 2076 10434 2078
rect 11237 2075 11303 2078
rect 4429 2002 4495 2005
rect 9438 2002 9444 2004
rect 4429 2000 9444 2002
rect 4429 1944 4434 2000
rect 4490 1944 9444 2000
rect 4429 1942 9444 1944
rect 4429 1939 4495 1942
rect 9438 1940 9444 1942
rect 9508 1940 9514 2004
rect 12934 1940 12940 2004
rect 13004 2002 13010 2004
rect 13353 2002 13419 2005
rect 13004 2000 13419 2002
rect 13004 1944 13358 2000
rect 13414 1944 13419 2000
rect 13004 1942 13419 1944
rect 13004 1940 13010 1942
rect 13353 1939 13419 1942
rect 4245 1866 4311 1869
rect 8886 1866 8892 1868
rect 4245 1864 8892 1866
rect 4245 1808 4250 1864
rect 4306 1808 8892 1864
rect 4245 1806 8892 1808
rect 4245 1803 4311 1806
rect 8886 1804 8892 1806
rect 8956 1804 8962 1868
rect 5993 1594 6059 1597
rect 9029 1594 9095 1597
rect 5993 1592 9095 1594
rect 5993 1536 5998 1592
rect 6054 1536 9034 1592
rect 9090 1536 9095 1592
rect 5993 1534 9095 1536
rect 5993 1531 6059 1534
rect 9029 1531 9095 1534
rect 12382 1532 12388 1596
rect 12452 1594 12458 1596
rect 12525 1594 12591 1597
rect 12452 1592 12591 1594
rect 12452 1536 12530 1592
rect 12586 1536 12591 1592
rect 12452 1534 12591 1536
rect 12452 1532 12458 1534
rect 12525 1531 12591 1534
rect 0 1458 480 1488
rect 14038 1458 14044 1460
rect 0 1398 14044 1458
rect 0 1368 480 1398
rect 14038 1396 14044 1398
rect 14108 1396 14114 1460
rect 10777 1322 10843 1325
rect 11278 1322 11284 1324
rect 10777 1320 11284 1322
rect 10777 1264 10782 1320
rect 10838 1264 11284 1320
rect 10777 1262 11284 1264
rect 10777 1259 10843 1262
rect 11278 1260 11284 1262
rect 11348 1260 11354 1324
rect 0 506 480 536
rect 2773 506 2839 509
rect 0 504 2839 506
rect 0 448 2778 504
rect 2834 448 2839 504
rect 0 446 2839 448
rect 0 416 480 446
rect 2773 443 2839 446
<< via3 >>
rect 12388 16084 12452 16148
rect 5882 15804 5946 15808
rect 5882 15748 5886 15804
rect 5886 15748 5942 15804
rect 5942 15748 5946 15804
rect 5882 15744 5946 15748
rect 5962 15804 6026 15808
rect 5962 15748 5966 15804
rect 5966 15748 6022 15804
rect 6022 15748 6026 15804
rect 5962 15744 6026 15748
rect 6042 15804 6106 15808
rect 6042 15748 6046 15804
rect 6046 15748 6102 15804
rect 6102 15748 6106 15804
rect 6042 15744 6106 15748
rect 6122 15804 6186 15808
rect 6122 15748 6126 15804
rect 6126 15748 6182 15804
rect 6182 15748 6186 15804
rect 6122 15744 6186 15748
rect 10813 15804 10877 15808
rect 10813 15748 10817 15804
rect 10817 15748 10873 15804
rect 10873 15748 10877 15804
rect 10813 15744 10877 15748
rect 10893 15804 10957 15808
rect 10893 15748 10897 15804
rect 10897 15748 10953 15804
rect 10953 15748 10957 15804
rect 10893 15744 10957 15748
rect 10973 15804 11037 15808
rect 10973 15748 10977 15804
rect 10977 15748 11033 15804
rect 11033 15748 11037 15804
rect 10973 15744 11037 15748
rect 11053 15804 11117 15808
rect 11053 15748 11057 15804
rect 11057 15748 11113 15804
rect 11113 15748 11117 15804
rect 11053 15744 11117 15748
rect 6868 15676 6932 15740
rect 3417 15260 3481 15264
rect 3417 15204 3421 15260
rect 3421 15204 3477 15260
rect 3477 15204 3481 15260
rect 3417 15200 3481 15204
rect 3497 15260 3561 15264
rect 3497 15204 3501 15260
rect 3501 15204 3557 15260
rect 3557 15204 3561 15260
rect 3497 15200 3561 15204
rect 3577 15260 3641 15264
rect 3577 15204 3581 15260
rect 3581 15204 3637 15260
rect 3637 15204 3641 15260
rect 3577 15200 3641 15204
rect 3657 15260 3721 15264
rect 3657 15204 3661 15260
rect 3661 15204 3717 15260
rect 3717 15204 3721 15260
rect 3657 15200 3721 15204
rect 8348 15260 8412 15264
rect 8348 15204 8352 15260
rect 8352 15204 8408 15260
rect 8408 15204 8412 15260
rect 8348 15200 8412 15204
rect 8428 15260 8492 15264
rect 8428 15204 8432 15260
rect 8432 15204 8488 15260
rect 8488 15204 8492 15260
rect 8428 15200 8492 15204
rect 8508 15260 8572 15264
rect 8508 15204 8512 15260
rect 8512 15204 8568 15260
rect 8568 15204 8572 15260
rect 8508 15200 8572 15204
rect 8588 15260 8652 15264
rect 8588 15204 8592 15260
rect 8592 15204 8648 15260
rect 8648 15204 8652 15260
rect 8588 15200 8652 15204
rect 13278 15260 13342 15264
rect 13278 15204 13282 15260
rect 13282 15204 13338 15260
rect 13338 15204 13342 15260
rect 13278 15200 13342 15204
rect 13358 15260 13422 15264
rect 13358 15204 13362 15260
rect 13362 15204 13418 15260
rect 13418 15204 13422 15260
rect 13358 15200 13422 15204
rect 13438 15260 13502 15264
rect 13438 15204 13442 15260
rect 13442 15204 13498 15260
rect 13498 15204 13502 15260
rect 13438 15200 13502 15204
rect 13518 15260 13582 15264
rect 13518 15204 13522 15260
rect 13522 15204 13578 15260
rect 13578 15204 13582 15260
rect 13518 15200 13582 15204
rect 6868 15132 6932 15196
rect 12204 14996 12268 15060
rect 5212 14724 5276 14788
rect 9628 14724 9692 14788
rect 9996 14724 10060 14788
rect 11652 14724 11716 14788
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 6122 14716 6186 14720
rect 6122 14660 6126 14716
rect 6126 14660 6182 14716
rect 6182 14660 6186 14716
rect 6122 14656 6186 14660
rect 10813 14716 10877 14720
rect 10813 14660 10817 14716
rect 10817 14660 10873 14716
rect 10873 14660 10877 14716
rect 10813 14656 10877 14660
rect 10893 14716 10957 14720
rect 10893 14660 10897 14716
rect 10897 14660 10953 14716
rect 10953 14660 10957 14716
rect 10893 14656 10957 14660
rect 10973 14716 11037 14720
rect 10973 14660 10977 14716
rect 10977 14660 11033 14716
rect 11033 14660 11037 14716
rect 10973 14656 11037 14660
rect 11053 14716 11117 14720
rect 11053 14660 11057 14716
rect 11057 14660 11113 14716
rect 11113 14660 11117 14716
rect 11053 14656 11117 14660
rect 5580 14588 5644 14652
rect 6316 14588 6380 14652
rect 7604 14316 7668 14380
rect 5396 14180 5460 14244
rect 13124 14316 13188 14380
rect 3417 14172 3481 14176
rect 3417 14116 3421 14172
rect 3421 14116 3477 14172
rect 3477 14116 3481 14172
rect 3417 14112 3481 14116
rect 3497 14172 3561 14176
rect 3497 14116 3501 14172
rect 3501 14116 3557 14172
rect 3557 14116 3561 14172
rect 3497 14112 3561 14116
rect 3577 14172 3641 14176
rect 3577 14116 3581 14172
rect 3581 14116 3637 14172
rect 3637 14116 3641 14172
rect 3577 14112 3641 14116
rect 3657 14172 3721 14176
rect 3657 14116 3661 14172
rect 3661 14116 3717 14172
rect 3717 14116 3721 14172
rect 3657 14112 3721 14116
rect 8348 14172 8412 14176
rect 8348 14116 8352 14172
rect 8352 14116 8408 14172
rect 8408 14116 8412 14172
rect 8348 14112 8412 14116
rect 8428 14172 8492 14176
rect 8428 14116 8432 14172
rect 8432 14116 8488 14172
rect 8488 14116 8492 14172
rect 8428 14112 8492 14116
rect 8508 14172 8572 14176
rect 8508 14116 8512 14172
rect 8512 14116 8568 14172
rect 8568 14116 8572 14172
rect 8508 14112 8572 14116
rect 8588 14172 8652 14176
rect 8588 14116 8592 14172
rect 8592 14116 8648 14172
rect 8648 14116 8652 14172
rect 8588 14112 8652 14116
rect 13278 14172 13342 14176
rect 13278 14116 13282 14172
rect 13282 14116 13338 14172
rect 13338 14116 13342 14172
rect 13278 14112 13342 14116
rect 13358 14172 13422 14176
rect 13358 14116 13362 14172
rect 13362 14116 13418 14172
rect 13418 14116 13422 14172
rect 13358 14112 13422 14116
rect 13438 14172 13502 14176
rect 13438 14116 13442 14172
rect 13442 14116 13498 14172
rect 13498 14116 13502 14172
rect 13438 14112 13502 14116
rect 13518 14172 13582 14176
rect 13518 14116 13522 14172
rect 13522 14116 13578 14172
rect 13578 14116 13582 14172
rect 13518 14112 13582 14116
rect 9628 14044 9692 14108
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 6122 13628 6186 13632
rect 6122 13572 6126 13628
rect 6126 13572 6182 13628
rect 6182 13572 6186 13628
rect 6122 13568 6186 13572
rect 8156 13772 8220 13836
rect 6684 13636 6748 13700
rect 12572 13636 12636 13700
rect 10813 13628 10877 13632
rect 10813 13572 10817 13628
rect 10817 13572 10873 13628
rect 10873 13572 10877 13628
rect 10813 13568 10877 13572
rect 10893 13628 10957 13632
rect 10893 13572 10897 13628
rect 10897 13572 10953 13628
rect 10953 13572 10957 13628
rect 10893 13568 10957 13572
rect 10973 13628 11037 13632
rect 10973 13572 10977 13628
rect 10977 13572 11033 13628
rect 11033 13572 11037 13628
rect 10973 13568 11037 13572
rect 11053 13628 11117 13632
rect 11053 13572 11057 13628
rect 11057 13572 11113 13628
rect 11113 13572 11117 13628
rect 11053 13568 11117 13572
rect 9812 13560 9876 13564
rect 9812 13504 9862 13560
rect 9862 13504 9876 13560
rect 9812 13500 9876 13504
rect 10548 13560 10612 13564
rect 10548 13504 10562 13560
rect 10562 13504 10612 13560
rect 10548 13500 10612 13504
rect 11836 13500 11900 13564
rect 12020 13500 12084 13564
rect 3417 13084 3481 13088
rect 3417 13028 3421 13084
rect 3421 13028 3477 13084
rect 3477 13028 3481 13084
rect 3417 13024 3481 13028
rect 3497 13084 3561 13088
rect 3497 13028 3501 13084
rect 3501 13028 3557 13084
rect 3557 13028 3561 13084
rect 3497 13024 3561 13028
rect 3577 13084 3641 13088
rect 3577 13028 3581 13084
rect 3581 13028 3637 13084
rect 3637 13028 3641 13084
rect 3577 13024 3641 13028
rect 3657 13084 3721 13088
rect 3657 13028 3661 13084
rect 3661 13028 3717 13084
rect 3717 13028 3721 13084
rect 3657 13024 3721 13028
rect 5580 13092 5644 13156
rect 8348 13084 8412 13088
rect 8348 13028 8352 13084
rect 8352 13028 8408 13084
rect 8408 13028 8412 13084
rect 8348 13024 8412 13028
rect 8428 13084 8492 13088
rect 8428 13028 8432 13084
rect 8432 13028 8488 13084
rect 8488 13028 8492 13084
rect 8428 13024 8492 13028
rect 8508 13084 8572 13088
rect 8508 13028 8512 13084
rect 8512 13028 8568 13084
rect 8568 13028 8572 13084
rect 8508 13024 8572 13028
rect 8588 13084 8652 13088
rect 8588 13028 8592 13084
rect 8592 13028 8648 13084
rect 8648 13028 8652 13084
rect 8588 13024 8652 13028
rect 13278 13084 13342 13088
rect 13278 13028 13282 13084
rect 13282 13028 13338 13084
rect 13338 13028 13342 13084
rect 13278 13024 13342 13028
rect 13358 13084 13422 13088
rect 13358 13028 13362 13084
rect 13362 13028 13418 13084
rect 13418 13028 13422 13084
rect 13358 13024 13422 13028
rect 13438 13084 13502 13088
rect 13438 13028 13442 13084
rect 13442 13028 13498 13084
rect 13498 13028 13502 13084
rect 13438 13024 13502 13028
rect 13518 13084 13582 13088
rect 13518 13028 13522 13084
rect 13522 13028 13578 13084
rect 13578 13028 13582 13084
rect 13518 13024 13582 13028
rect 6500 12880 6564 12884
rect 6500 12824 6550 12880
rect 6550 12824 6564 12880
rect 6500 12820 6564 12824
rect 7420 12956 7484 13020
rect 9260 12956 9324 13020
rect 10180 12956 10244 13020
rect 11284 12820 11348 12884
rect 9444 12548 9508 12612
rect 10364 12548 10428 12612
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 6122 12540 6186 12544
rect 6122 12484 6126 12540
rect 6126 12484 6182 12540
rect 6182 12484 6186 12540
rect 6122 12480 6186 12484
rect 10813 12540 10877 12544
rect 10813 12484 10817 12540
rect 10817 12484 10873 12540
rect 10873 12484 10877 12540
rect 10813 12480 10877 12484
rect 10893 12540 10957 12544
rect 10893 12484 10897 12540
rect 10897 12484 10953 12540
rect 10953 12484 10957 12540
rect 10893 12480 10957 12484
rect 10973 12540 11037 12544
rect 10973 12484 10977 12540
rect 10977 12484 11033 12540
rect 11033 12484 11037 12540
rect 10973 12480 11037 12484
rect 11053 12540 11117 12544
rect 11053 12484 11057 12540
rect 11057 12484 11113 12540
rect 11113 12484 11117 12540
rect 11053 12480 11117 12484
rect 4844 12412 4908 12476
rect 4292 12276 4356 12340
rect 3004 12140 3068 12204
rect 3417 11996 3481 12000
rect 3417 11940 3421 11996
rect 3421 11940 3477 11996
rect 3477 11940 3481 11996
rect 3417 11936 3481 11940
rect 3497 11996 3561 12000
rect 3497 11940 3501 11996
rect 3501 11940 3557 11996
rect 3557 11940 3561 11996
rect 3497 11936 3561 11940
rect 3577 11996 3641 12000
rect 3577 11940 3581 11996
rect 3581 11940 3637 11996
rect 3637 11940 3641 11996
rect 3577 11936 3641 11940
rect 3657 11996 3721 12000
rect 3657 11940 3661 11996
rect 3661 11940 3717 11996
rect 3717 11940 3721 11996
rect 3657 11936 3721 11940
rect 7420 12004 7484 12068
rect 8348 11996 8412 12000
rect 8348 11940 8352 11996
rect 8352 11940 8408 11996
rect 8408 11940 8412 11996
rect 8348 11936 8412 11940
rect 8428 11996 8492 12000
rect 8428 11940 8432 11996
rect 8432 11940 8488 11996
rect 8488 11940 8492 11996
rect 8428 11936 8492 11940
rect 8508 11996 8572 12000
rect 8508 11940 8512 11996
rect 8512 11940 8568 11996
rect 8568 11940 8572 11996
rect 8508 11936 8572 11940
rect 8588 11996 8652 12000
rect 8588 11940 8592 11996
rect 8592 11940 8648 11996
rect 8648 11940 8652 11996
rect 8588 11936 8652 11940
rect 13278 11996 13342 12000
rect 13278 11940 13282 11996
rect 13282 11940 13338 11996
rect 13338 11940 13342 11996
rect 13278 11936 13342 11940
rect 13358 11996 13422 12000
rect 13358 11940 13362 11996
rect 13362 11940 13418 11996
rect 13418 11940 13422 11996
rect 13358 11936 13422 11940
rect 13438 11996 13502 12000
rect 13438 11940 13442 11996
rect 13442 11940 13498 11996
rect 13498 11940 13502 11996
rect 13438 11936 13502 11940
rect 13518 11996 13582 12000
rect 13518 11940 13522 11996
rect 13522 11940 13578 11996
rect 13578 11940 13582 11996
rect 13518 11936 13582 11940
rect 9076 11868 9140 11932
rect 6316 11460 6380 11524
rect 7972 11460 8036 11524
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 6122 11452 6186 11456
rect 6122 11396 6126 11452
rect 6126 11396 6182 11452
rect 6182 11396 6186 11452
rect 6122 11392 6186 11396
rect 10813 11452 10877 11456
rect 10813 11396 10817 11452
rect 10817 11396 10873 11452
rect 10873 11396 10877 11452
rect 10813 11392 10877 11396
rect 10893 11452 10957 11456
rect 10893 11396 10897 11452
rect 10897 11396 10953 11452
rect 10953 11396 10957 11452
rect 10893 11392 10957 11396
rect 10973 11452 11037 11456
rect 10973 11396 10977 11452
rect 10977 11396 11033 11452
rect 11033 11396 11037 11452
rect 10973 11392 11037 11396
rect 11053 11452 11117 11456
rect 11053 11396 11057 11452
rect 11057 11396 11113 11452
rect 11113 11396 11117 11452
rect 11053 11392 11117 11396
rect 6316 11324 6380 11388
rect 8754 11188 8818 11252
rect 3417 10908 3481 10912
rect 3417 10852 3421 10908
rect 3421 10852 3477 10908
rect 3477 10852 3481 10908
rect 3417 10848 3481 10852
rect 3497 10908 3561 10912
rect 3497 10852 3501 10908
rect 3501 10852 3557 10908
rect 3557 10852 3561 10908
rect 3497 10848 3561 10852
rect 3577 10908 3641 10912
rect 3577 10852 3581 10908
rect 3581 10852 3637 10908
rect 3637 10852 3641 10908
rect 3577 10848 3641 10852
rect 3657 10908 3721 10912
rect 3657 10852 3661 10908
rect 3661 10852 3717 10908
rect 3717 10852 3721 10908
rect 3657 10848 3721 10852
rect 11836 11248 11900 11252
rect 11836 11192 11886 11248
rect 11886 11192 11900 11248
rect 11836 11188 11900 11192
rect 9444 10916 9508 10980
rect 9812 10976 9876 10980
rect 9812 10920 9826 10976
rect 9826 10920 9876 10976
rect 9812 10916 9876 10920
rect 8348 10908 8412 10912
rect 8348 10852 8352 10908
rect 8352 10852 8408 10908
rect 8408 10852 8412 10908
rect 8348 10848 8412 10852
rect 8428 10908 8492 10912
rect 8428 10852 8432 10908
rect 8432 10852 8488 10908
rect 8488 10852 8492 10908
rect 8428 10848 8492 10852
rect 8508 10908 8572 10912
rect 8508 10852 8512 10908
rect 8512 10852 8568 10908
rect 8568 10852 8572 10908
rect 8508 10848 8572 10852
rect 8588 10908 8652 10912
rect 8588 10852 8592 10908
rect 8592 10852 8648 10908
rect 8648 10852 8652 10908
rect 8588 10848 8652 10852
rect 7604 10780 7668 10844
rect 9260 10840 9324 10844
rect 9260 10784 9310 10840
rect 9310 10784 9324 10840
rect 9260 10780 9324 10784
rect 9996 10780 10060 10844
rect 13278 10908 13342 10912
rect 13278 10852 13282 10908
rect 13282 10852 13338 10908
rect 13338 10852 13342 10908
rect 13278 10848 13342 10852
rect 13358 10908 13422 10912
rect 13358 10852 13362 10908
rect 13362 10852 13418 10908
rect 13418 10852 13422 10908
rect 13358 10848 13422 10852
rect 13438 10908 13502 10912
rect 13438 10852 13442 10908
rect 13442 10852 13498 10908
rect 13498 10852 13502 10908
rect 13438 10848 13502 10852
rect 13518 10908 13582 10912
rect 13518 10852 13522 10908
rect 13522 10852 13578 10908
rect 13578 10852 13582 10908
rect 13518 10848 13582 10852
rect 12388 10780 12452 10844
rect 10364 10568 10428 10572
rect 10364 10512 10414 10568
rect 10414 10512 10428 10568
rect 10364 10508 10428 10512
rect 6500 10432 6564 10436
rect 6500 10376 6514 10432
rect 6514 10376 6564 10432
rect 6500 10372 6564 10376
rect 6684 10372 6748 10436
rect 7788 10372 7852 10436
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 6122 10364 6186 10368
rect 6122 10308 6126 10364
rect 6126 10308 6182 10364
rect 6182 10308 6186 10364
rect 6122 10304 6186 10308
rect 10813 10364 10877 10368
rect 10813 10308 10817 10364
rect 10817 10308 10873 10364
rect 10873 10308 10877 10364
rect 10813 10304 10877 10308
rect 10893 10364 10957 10368
rect 10893 10308 10897 10364
rect 10897 10308 10953 10364
rect 10953 10308 10957 10364
rect 10893 10304 10957 10308
rect 10973 10364 11037 10368
rect 10973 10308 10977 10364
rect 10977 10308 11033 10364
rect 11033 10308 11037 10364
rect 10973 10304 11037 10308
rect 11053 10364 11117 10368
rect 11053 10308 11057 10364
rect 11057 10308 11113 10364
rect 11113 10308 11117 10364
rect 11053 10304 11117 10308
rect 5212 10236 5276 10300
rect 7236 10236 7300 10300
rect 7420 10236 7484 10300
rect 11836 10372 11900 10436
rect 13860 10372 13924 10436
rect 7052 10100 7116 10164
rect 6316 9964 6380 10028
rect 6868 9964 6932 10028
rect 4844 9828 4908 9892
rect 5212 9828 5276 9892
rect 9996 9828 10060 9892
rect 10548 9828 10612 9892
rect 12756 9828 12820 9892
rect 3417 9820 3481 9824
rect 3417 9764 3421 9820
rect 3421 9764 3477 9820
rect 3477 9764 3481 9820
rect 3417 9760 3481 9764
rect 3497 9820 3561 9824
rect 3497 9764 3501 9820
rect 3501 9764 3557 9820
rect 3557 9764 3561 9820
rect 3497 9760 3561 9764
rect 3577 9820 3641 9824
rect 3577 9764 3581 9820
rect 3581 9764 3637 9820
rect 3637 9764 3641 9820
rect 3577 9760 3641 9764
rect 3657 9820 3721 9824
rect 3657 9764 3661 9820
rect 3661 9764 3717 9820
rect 3717 9764 3721 9820
rect 3657 9760 3721 9764
rect 8348 9820 8412 9824
rect 8348 9764 8352 9820
rect 8352 9764 8408 9820
rect 8408 9764 8412 9820
rect 8348 9760 8412 9764
rect 8428 9820 8492 9824
rect 8428 9764 8432 9820
rect 8432 9764 8488 9820
rect 8488 9764 8492 9820
rect 8428 9760 8492 9764
rect 8508 9820 8572 9824
rect 8508 9764 8512 9820
rect 8512 9764 8568 9820
rect 8568 9764 8572 9820
rect 8508 9760 8572 9764
rect 8588 9820 8652 9824
rect 8588 9764 8592 9820
rect 8592 9764 8648 9820
rect 8648 9764 8652 9820
rect 8588 9760 8652 9764
rect 13278 9820 13342 9824
rect 13278 9764 13282 9820
rect 13282 9764 13338 9820
rect 13338 9764 13342 9820
rect 13278 9760 13342 9764
rect 13358 9820 13422 9824
rect 13358 9764 13362 9820
rect 13362 9764 13418 9820
rect 13418 9764 13422 9820
rect 13358 9760 13422 9764
rect 13438 9820 13502 9824
rect 13438 9764 13442 9820
rect 13442 9764 13498 9820
rect 13498 9764 13502 9820
rect 13438 9760 13502 9764
rect 13518 9820 13582 9824
rect 13518 9764 13522 9820
rect 13522 9764 13578 9820
rect 13578 9764 13582 9820
rect 13518 9760 13582 9764
rect 9076 9692 9140 9756
rect 10180 9752 10244 9756
rect 10180 9696 10194 9752
rect 10194 9696 10244 9752
rect 10180 9692 10244 9696
rect 11652 9692 11716 9756
rect 14044 9692 14108 9756
rect 10548 9556 10612 9620
rect 6684 9284 6748 9348
rect 10548 9284 10612 9348
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 6122 9276 6186 9280
rect 6122 9220 6126 9276
rect 6126 9220 6182 9276
rect 6182 9220 6186 9276
rect 6122 9216 6186 9220
rect 10813 9276 10877 9280
rect 10813 9220 10817 9276
rect 10817 9220 10873 9276
rect 10873 9220 10877 9276
rect 10813 9216 10877 9220
rect 10893 9276 10957 9280
rect 10893 9220 10897 9276
rect 10897 9220 10953 9276
rect 10953 9220 10957 9276
rect 10893 9216 10957 9220
rect 10973 9276 11037 9280
rect 10973 9220 10977 9276
rect 10977 9220 11033 9276
rect 11033 9220 11037 9276
rect 10973 9216 11037 9220
rect 11053 9276 11117 9280
rect 11053 9220 11057 9276
rect 11057 9220 11113 9276
rect 11113 9220 11117 9276
rect 11053 9216 11117 9220
rect 6316 9148 6380 9212
rect 9628 9148 9692 9212
rect 10548 9148 10612 9212
rect 11652 9148 11716 9212
rect 12204 9208 12268 9212
rect 12204 9152 12218 9208
rect 12218 9152 12268 9208
rect 12204 9148 12268 9152
rect 12388 9208 12452 9212
rect 12388 9152 12438 9208
rect 12438 9152 12452 9208
rect 12388 9148 12452 9152
rect 11468 8876 11532 8940
rect 8892 8740 8956 8804
rect 12204 8740 12268 8804
rect 13676 8740 13740 8804
rect 3417 8732 3481 8736
rect 3417 8676 3421 8732
rect 3421 8676 3477 8732
rect 3477 8676 3481 8732
rect 3417 8672 3481 8676
rect 3497 8732 3561 8736
rect 3497 8676 3501 8732
rect 3501 8676 3557 8732
rect 3557 8676 3561 8732
rect 3497 8672 3561 8676
rect 3577 8732 3641 8736
rect 3577 8676 3581 8732
rect 3581 8676 3637 8732
rect 3637 8676 3641 8732
rect 3577 8672 3641 8676
rect 3657 8732 3721 8736
rect 3657 8676 3661 8732
rect 3661 8676 3717 8732
rect 3717 8676 3721 8732
rect 3657 8672 3721 8676
rect 8348 8732 8412 8736
rect 8348 8676 8352 8732
rect 8352 8676 8408 8732
rect 8408 8676 8412 8732
rect 8348 8672 8412 8676
rect 8428 8732 8492 8736
rect 8428 8676 8432 8732
rect 8432 8676 8488 8732
rect 8488 8676 8492 8732
rect 8428 8672 8492 8676
rect 8508 8732 8572 8736
rect 8508 8676 8512 8732
rect 8512 8676 8568 8732
rect 8568 8676 8572 8732
rect 8508 8672 8572 8676
rect 8588 8732 8652 8736
rect 8588 8676 8592 8732
rect 8592 8676 8648 8732
rect 8648 8676 8652 8732
rect 8588 8672 8652 8676
rect 13278 8732 13342 8736
rect 13278 8676 13282 8732
rect 13282 8676 13338 8732
rect 13338 8676 13342 8732
rect 13278 8672 13342 8676
rect 13358 8732 13422 8736
rect 13358 8676 13362 8732
rect 13362 8676 13418 8732
rect 13418 8676 13422 8732
rect 13358 8672 13422 8676
rect 13438 8732 13502 8736
rect 13438 8676 13442 8732
rect 13442 8676 13498 8732
rect 13498 8676 13502 8732
rect 13438 8672 13502 8676
rect 13518 8732 13582 8736
rect 13518 8676 13522 8732
rect 13522 8676 13578 8732
rect 13578 8676 13582 8732
rect 13518 8672 13582 8676
rect 3924 8604 3988 8668
rect 6316 8468 6380 8532
rect 7604 8604 7668 8668
rect 4660 8196 4724 8260
rect 5396 8196 5460 8260
rect 9260 8256 9324 8260
rect 9260 8200 9310 8256
rect 9310 8200 9324 8256
rect 9260 8196 9324 8200
rect 9628 8196 9692 8260
rect 11284 8196 11348 8260
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 6122 8188 6186 8192
rect 6122 8132 6126 8188
rect 6126 8132 6182 8188
rect 6182 8132 6186 8188
rect 6122 8128 6186 8132
rect 10813 8188 10877 8192
rect 10813 8132 10817 8188
rect 10817 8132 10873 8188
rect 10873 8132 10877 8188
rect 10813 8128 10877 8132
rect 10893 8188 10957 8192
rect 10893 8132 10897 8188
rect 10897 8132 10953 8188
rect 10953 8132 10957 8188
rect 10893 8128 10957 8132
rect 10973 8188 11037 8192
rect 10973 8132 10977 8188
rect 10977 8132 11033 8188
rect 11033 8132 11037 8188
rect 10973 8128 11037 8132
rect 11053 8188 11117 8192
rect 11053 8132 11057 8188
rect 11057 8132 11113 8188
rect 11113 8132 11117 8188
rect 11053 8128 11117 8132
rect 10364 8060 10428 8124
rect 4844 7652 4908 7716
rect 11836 7788 11900 7852
rect 12940 7788 13004 7852
rect 6500 7652 6564 7716
rect 3417 7644 3481 7648
rect 3417 7588 3421 7644
rect 3421 7588 3477 7644
rect 3477 7588 3481 7644
rect 3417 7584 3481 7588
rect 3497 7644 3561 7648
rect 3497 7588 3501 7644
rect 3501 7588 3557 7644
rect 3557 7588 3561 7644
rect 3497 7584 3561 7588
rect 3577 7644 3641 7648
rect 3577 7588 3581 7644
rect 3581 7588 3637 7644
rect 3637 7588 3641 7644
rect 3577 7584 3641 7588
rect 3657 7644 3721 7648
rect 3657 7588 3661 7644
rect 3661 7588 3717 7644
rect 3717 7588 3721 7644
rect 3657 7584 3721 7588
rect 8348 7644 8412 7648
rect 8348 7588 8352 7644
rect 8352 7588 8408 7644
rect 8408 7588 8412 7644
rect 8348 7584 8412 7588
rect 8428 7644 8492 7648
rect 8428 7588 8432 7644
rect 8432 7588 8488 7644
rect 8488 7588 8492 7644
rect 8428 7584 8492 7588
rect 8508 7644 8572 7648
rect 8508 7588 8512 7644
rect 8512 7588 8568 7644
rect 8568 7588 8572 7644
rect 8508 7584 8572 7588
rect 8588 7644 8652 7648
rect 8588 7588 8592 7644
rect 8592 7588 8648 7644
rect 8648 7588 8652 7644
rect 8588 7584 8652 7588
rect 13278 7644 13342 7648
rect 13278 7588 13282 7644
rect 13282 7588 13338 7644
rect 13338 7588 13342 7644
rect 13278 7584 13342 7588
rect 13358 7644 13422 7648
rect 13358 7588 13362 7644
rect 13362 7588 13418 7644
rect 13418 7588 13422 7644
rect 13358 7584 13422 7588
rect 13438 7644 13502 7648
rect 13438 7588 13442 7644
rect 13442 7588 13498 7644
rect 13498 7588 13502 7644
rect 13438 7584 13502 7588
rect 13518 7644 13582 7648
rect 13518 7588 13522 7644
rect 13522 7588 13578 7644
rect 13578 7588 13582 7644
rect 13518 7584 13582 7588
rect 9076 7516 9140 7580
rect 9444 7516 9508 7580
rect 6500 7108 6564 7172
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 6122 7100 6186 7104
rect 6122 7044 6126 7100
rect 6126 7044 6182 7100
rect 6182 7044 6186 7100
rect 6122 7040 6186 7044
rect 10813 7100 10877 7104
rect 10813 7044 10817 7100
rect 10817 7044 10873 7100
rect 10873 7044 10877 7100
rect 10813 7040 10877 7044
rect 10893 7100 10957 7104
rect 10893 7044 10897 7100
rect 10897 7044 10953 7100
rect 10953 7044 10957 7100
rect 10893 7040 10957 7044
rect 10973 7100 11037 7104
rect 10973 7044 10977 7100
rect 10977 7044 11033 7100
rect 11033 7044 11037 7100
rect 10973 7040 11037 7044
rect 11053 7100 11117 7104
rect 11053 7044 11057 7100
rect 11057 7044 11113 7100
rect 11113 7044 11117 7100
rect 11053 7040 11117 7044
rect 4292 6972 4356 7036
rect 9812 7032 9876 7036
rect 9812 6976 9862 7032
rect 9862 6976 9876 7032
rect 9812 6972 9876 6976
rect 7236 6836 7300 6900
rect 9076 6836 9140 6900
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 10548 6488 10612 6492
rect 10548 6432 10598 6488
rect 10598 6432 10612 6488
rect 10548 6428 10612 6432
rect 11836 6156 11900 6220
rect 6316 6020 6380 6084
rect 9076 6020 9140 6084
rect 10180 6020 10244 6084
rect 11468 6020 11532 6084
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 5028 5884 5092 5948
rect 6500 5884 6564 5948
rect 9812 5884 9876 5948
rect 12572 5748 12636 5812
rect 7236 5476 7300 5540
rect 12388 5476 12452 5540
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 12572 5340 12636 5404
rect 7236 5068 7300 5132
rect 11468 4932 11532 4996
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 8892 4796 8956 4860
rect 11652 4796 11716 4860
rect 12756 4796 12820 4860
rect 11836 4584 11900 4588
rect 11836 4528 11886 4584
rect 11886 4528 11900 4584
rect 11836 4524 11900 4528
rect 6868 4388 6932 4452
rect 12388 4524 12452 4588
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 8892 4252 8956 4316
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 9260 4252 9324 4316
rect 9628 4252 9692 4316
rect 6500 4116 6564 4180
rect 3004 3844 3068 3908
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 5580 3768 5644 3772
rect 5580 3712 5630 3768
rect 5630 3712 5644 3768
rect 5580 3708 5644 3712
rect 3924 3572 3988 3636
rect 13676 3844 13740 3908
rect 5212 3300 5276 3364
rect 7052 3360 7116 3364
rect 7052 3304 7102 3360
rect 7102 3304 7116 3360
rect 7052 3300 7116 3304
rect 7420 3360 7484 3364
rect 7420 3304 7434 3360
rect 7434 3304 7484 3360
rect 7420 3300 7484 3304
rect 12020 3436 12084 3500
rect 13860 3496 13924 3500
rect 13860 3440 13874 3496
rect 13874 3440 13924 3496
rect 13860 3436 13924 3440
rect 10548 3300 10612 3364
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 8892 3164 8956 3228
rect 12204 3164 12268 3228
rect 7052 2892 7116 2956
rect 7972 2756 8036 2820
rect 9996 2816 10060 2820
rect 9996 2760 10046 2816
rect 10046 2760 10060 2816
rect 9996 2756 10060 2760
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 6316 2620 6380 2684
rect 7788 2620 7852 2684
rect 8156 2680 8220 2684
rect 8156 2624 8206 2680
rect 8206 2624 8220 2680
rect 8156 2620 8220 2624
rect 10180 2620 10244 2684
rect 11284 2680 11348 2684
rect 11284 2624 11334 2680
rect 11334 2624 11348 2680
rect 11284 2620 11348 2624
rect 6684 2484 6748 2548
rect 7052 2484 7116 2548
rect 7604 2348 7668 2412
rect 13124 2484 13188 2548
rect 12572 2348 12636 2412
rect 5396 2212 5460 2276
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
rect 10364 2076 10428 2140
rect 9444 1940 9508 2004
rect 12940 1940 13004 2004
rect 8892 1804 8956 1868
rect 12388 1532 12452 1596
rect 14044 1396 14108 1460
rect 11284 1260 11348 1324
<< metal4 >>
rect 12387 16148 12453 16149
rect 12387 16084 12388 16148
rect 12452 16084 12453 16148
rect 12387 16083 12453 16084
rect 3409 15264 3729 15824
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 14176 3729 15200
rect 5874 15808 6195 15824
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6195 15808
rect 5211 14788 5277 14789
rect 5211 14724 5212 14788
rect 5276 14724 5277 14788
rect 5211 14723 5277 14724
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 13088 3729 14112
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3003 12204 3069 12205
rect 3003 12140 3004 12204
rect 3068 12140 3069 12204
rect 3003 12139 3069 12140
rect 3006 3909 3066 12139
rect 3409 12000 3729 13024
rect 4843 12476 4909 12477
rect 4843 12412 4844 12476
rect 4908 12412 4909 12476
rect 4843 12411 4909 12412
rect 4291 12340 4357 12341
rect 4291 12276 4292 12340
rect 4356 12276 4357 12340
rect 4291 12275 4357 12276
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 10912 3729 11936
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 9824 3729 10848
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 8736 3729 9760
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 7648 3729 8672
rect 3923 8668 3989 8669
rect 3923 8604 3924 8668
rect 3988 8604 3989 8668
rect 3923 8603 3989 8604
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 6560 3729 7584
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 5472 3729 6496
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3003 3908 3069 3909
rect 3003 3844 3004 3908
rect 3068 3844 3069 3908
rect 3003 3843 3069 3844
rect 3409 3296 3729 4320
rect 3926 3637 3986 8603
rect 4294 7037 4354 12275
rect 4846 9893 4906 12411
rect 5214 10301 5274 14723
rect 5874 14720 6195 15744
rect 6867 15740 6933 15741
rect 6867 15676 6868 15740
rect 6932 15676 6933 15740
rect 6867 15675 6933 15676
rect 6870 15197 6930 15675
rect 8340 15264 8660 15824
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 6867 15196 6933 15197
rect 6867 15132 6868 15196
rect 6932 15132 6933 15196
rect 6867 15131 6933 15132
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6195 14720
rect 5579 14652 5645 14653
rect 5579 14588 5580 14652
rect 5644 14588 5645 14652
rect 5579 14587 5645 14588
rect 5395 14244 5461 14245
rect 5395 14180 5396 14244
rect 5460 14180 5461 14244
rect 5395 14179 5461 14180
rect 5211 10300 5277 10301
rect 5211 10236 5212 10300
rect 5276 10236 5277 10300
rect 5211 10235 5277 10236
rect 5398 10026 5458 14179
rect 5582 13157 5642 14587
rect 5874 13632 6195 14656
rect 6315 14652 6381 14653
rect 6315 14588 6316 14652
rect 6380 14588 6381 14652
rect 6315 14587 6381 14588
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6195 13632
rect 5579 13156 5645 13157
rect 5579 13092 5580 13156
rect 5644 13092 5645 13156
rect 5579 13091 5645 13092
rect 5030 9966 5458 10026
rect 4843 9892 4909 9893
rect 4843 9828 4844 9892
rect 4908 9828 4909 9892
rect 4843 9827 4909 9828
rect 4662 8261 4722 9062
rect 4659 8260 4725 8261
rect 4659 8196 4660 8260
rect 4724 8196 4725 8260
rect 4659 8195 4725 8196
rect 4843 7716 4909 7717
rect 4843 7652 4844 7716
rect 4908 7652 4909 7716
rect 4843 7651 4909 7652
rect 4291 7036 4357 7037
rect 4291 6972 4292 7036
rect 4356 6972 4357 7036
rect 4291 6971 4357 6972
rect 4846 4538 4906 7651
rect 5030 5949 5090 9966
rect 5211 9892 5277 9893
rect 5211 9828 5212 9892
rect 5276 9828 5277 9892
rect 5211 9827 5277 9828
rect 5027 5948 5093 5949
rect 5027 5884 5028 5948
rect 5092 5884 5093 5948
rect 5027 5883 5093 5884
rect 3923 3636 3989 3637
rect 3923 3572 3924 3636
rect 3988 3572 3989 3636
rect 3923 3571 3989 3572
rect 5214 3365 5274 9827
rect 5395 8260 5461 8261
rect 5395 8196 5396 8260
rect 5460 8196 5461 8260
rect 5395 8195 5461 8196
rect 5211 3364 5277 3365
rect 5211 3300 5212 3364
rect 5276 3300 5277 3364
rect 5211 3299 5277 3300
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 2208 3729 3232
rect 5398 2277 5458 8195
rect 5582 3773 5642 13091
rect 5874 12544 6195 13568
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6195 12544
rect 5874 11456 6195 12480
rect 6318 11525 6378 14587
rect 6683 13700 6749 13701
rect 6683 13636 6684 13700
rect 6748 13636 6749 13700
rect 6683 13635 6749 13636
rect 6499 12884 6565 12885
rect 6499 12820 6500 12884
rect 6564 12820 6565 12884
rect 6499 12819 6565 12820
rect 6315 11524 6381 11525
rect 6315 11460 6316 11524
rect 6380 11460 6381 11524
rect 6315 11459 6381 11460
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6195 11456
rect 5874 10368 6195 11392
rect 6315 11388 6381 11389
rect 6315 11324 6316 11388
rect 6380 11324 6381 11388
rect 6315 11323 6381 11324
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6195 10368
rect 5874 9280 6195 10304
rect 6318 10029 6378 11323
rect 6502 10437 6562 12819
rect 6686 10437 6746 13635
rect 6870 12882 6930 15131
rect 7603 14380 7669 14381
rect 7603 14316 7604 14380
rect 7668 14316 7669 14380
rect 7603 14315 7669 14316
rect 7419 13020 7485 13021
rect 7419 12956 7420 13020
rect 7484 12956 7485 13020
rect 7419 12955 7485 12956
rect 6870 12822 7298 12882
rect 6499 10436 6565 10437
rect 6499 10372 6500 10436
rect 6564 10372 6565 10436
rect 6499 10371 6565 10372
rect 6683 10436 6749 10437
rect 6683 10372 6684 10436
rect 6748 10372 6749 10436
rect 6683 10371 6749 10372
rect 7238 10301 7298 12822
rect 7422 12069 7482 12955
rect 7419 12068 7485 12069
rect 7419 12004 7420 12068
rect 7484 12004 7485 12068
rect 7419 12003 7485 12004
rect 7606 10845 7666 14315
rect 8340 14176 8660 15200
rect 10805 15808 11125 15824
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 9627 14788 9693 14789
rect 9627 14724 9628 14788
rect 9692 14724 9693 14788
rect 9627 14723 9693 14724
rect 9995 14788 10061 14789
rect 9995 14724 9996 14788
rect 10060 14724 10061 14788
rect 9995 14723 10061 14724
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8155 13836 8221 13837
rect 8155 13772 8156 13836
rect 8220 13772 8221 13836
rect 8155 13771 8221 13772
rect 7971 11524 8037 11525
rect 7971 11460 7972 11524
rect 8036 11460 8037 11524
rect 7971 11459 8037 11460
rect 7603 10844 7669 10845
rect 7603 10780 7604 10844
rect 7668 10780 7669 10844
rect 7603 10779 7669 10780
rect 7787 10436 7853 10437
rect 7787 10372 7788 10436
rect 7852 10372 7853 10436
rect 7787 10371 7853 10372
rect 7235 10300 7301 10301
rect 7235 10236 7236 10300
rect 7300 10236 7301 10300
rect 7235 10235 7301 10236
rect 7419 10300 7485 10301
rect 7419 10236 7420 10300
rect 7484 10236 7485 10300
rect 7419 10235 7485 10236
rect 7051 10164 7117 10165
rect 7051 10100 7052 10164
rect 7116 10100 7117 10164
rect 7051 10099 7117 10100
rect 6315 10028 6381 10029
rect 6315 9964 6316 10028
rect 6380 9964 6381 10028
rect 6315 9963 6381 9964
rect 6867 10028 6933 10029
rect 6867 9964 6868 10028
rect 6932 9964 6933 10028
rect 6867 9963 6933 9964
rect 6683 9348 6749 9349
rect 6683 9284 6684 9348
rect 6748 9284 6749 9348
rect 6683 9283 6749 9284
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6195 9280
rect 5874 8192 6195 9216
rect 6315 9212 6381 9213
rect 6315 9148 6316 9212
rect 6380 9148 6381 9212
rect 6315 9147 6381 9148
rect 6318 8533 6378 9147
rect 6315 8532 6381 8533
rect 6315 8468 6316 8532
rect 6380 8468 6381 8532
rect 6315 8467 6381 8468
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6195 8192
rect 5874 7104 6195 8128
rect 6499 7716 6565 7717
rect 6499 7652 6500 7716
rect 6564 7652 6565 7716
rect 6499 7651 6565 7652
rect 6502 7173 6562 7651
rect 6499 7172 6565 7173
rect 6499 7108 6500 7172
rect 6564 7108 6565 7172
rect 6499 7107 6565 7108
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6195 7104
rect 5874 6016 6195 7040
rect 6315 6084 6381 6085
rect 6315 6020 6316 6084
rect 6380 6020 6381 6084
rect 6315 6019 6381 6020
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5874 3840 6195 4864
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5579 3772 5645 3773
rect 5579 3708 5580 3772
rect 5644 3708 5645 3772
rect 5579 3707 5645 3708
rect 5874 2752 6195 3776
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 5395 2276 5461 2277
rect 5395 2212 5396 2276
rect 5460 2212 5461 2276
rect 5395 2211 5461 2212
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 5874 2128 6195 2688
rect 6318 2685 6378 6019
rect 6499 5948 6565 5949
rect 6499 5884 6500 5948
rect 6564 5884 6565 5948
rect 6499 5883 6565 5884
rect 6502 4181 6562 5883
rect 6499 4180 6565 4181
rect 6499 4116 6500 4180
rect 6564 4116 6565 4180
rect 6499 4115 6565 4116
rect 6315 2684 6381 2685
rect 6315 2620 6316 2684
rect 6380 2620 6381 2684
rect 6315 2619 6381 2620
rect 6686 2549 6746 9283
rect 6870 4453 6930 9963
rect 6867 4452 6933 4453
rect 6867 4388 6868 4452
rect 6932 4388 6933 4452
rect 6867 4387 6933 4388
rect 7054 3365 7114 10099
rect 7238 6901 7298 10235
rect 7235 6900 7301 6901
rect 7235 6836 7236 6900
rect 7300 6836 7301 6900
rect 7235 6835 7301 6836
rect 7235 5540 7301 5541
rect 7235 5476 7236 5540
rect 7300 5476 7301 5540
rect 7235 5475 7301 5476
rect 7238 5133 7298 5475
rect 7235 5132 7301 5133
rect 7235 5068 7236 5132
rect 7300 5068 7301 5132
rect 7235 5067 7301 5068
rect 7422 3365 7482 10235
rect 7603 8668 7669 8669
rect 7603 8604 7604 8668
rect 7668 8604 7669 8668
rect 7603 8603 7669 8604
rect 7051 3364 7117 3365
rect 7051 3300 7052 3364
rect 7116 3300 7117 3364
rect 7051 3299 7117 3300
rect 7419 3364 7485 3365
rect 7419 3300 7420 3364
rect 7484 3300 7485 3364
rect 7419 3299 7485 3300
rect 7051 2956 7117 2957
rect 7051 2892 7052 2956
rect 7116 2892 7117 2956
rect 7051 2891 7117 2892
rect 7054 2549 7114 2891
rect 6683 2548 6749 2549
rect 6683 2484 6684 2548
rect 6748 2484 6749 2548
rect 6683 2483 6749 2484
rect 7051 2548 7117 2549
rect 7051 2484 7052 2548
rect 7116 2484 7117 2548
rect 7051 2483 7117 2484
rect 7606 2413 7666 8603
rect 7790 2685 7850 10371
rect 7974 2821 8034 11459
rect 7971 2820 8037 2821
rect 7971 2756 7972 2820
rect 8036 2756 8037 2820
rect 7971 2755 8037 2756
rect 8158 2685 8218 13771
rect 8340 13088 8660 14112
rect 9630 14109 9690 14723
rect 9627 14108 9693 14109
rect 9627 14044 9628 14108
rect 9692 14044 9693 14108
rect 9627 14043 9693 14044
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 12000 8660 13024
rect 9259 13020 9325 13021
rect 9259 12956 9260 13020
rect 9324 12956 9325 13020
rect 9259 12955 9325 12956
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 10912 8660 11936
rect 9075 11932 9141 11933
rect 9075 11868 9076 11932
rect 9140 11868 9141 11932
rect 9075 11867 9141 11868
rect 8753 11252 8819 11253
rect 8753 11188 8754 11252
rect 8818 11250 8819 11252
rect 9078 11250 9138 11867
rect 8818 11190 9138 11250
rect 8818 11188 8819 11190
rect 8753 11187 8819 11188
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 9824 8660 10848
rect 9262 10845 9322 12955
rect 9443 12612 9509 12613
rect 9443 12548 9444 12612
rect 9508 12548 9509 12612
rect 9443 12547 9509 12548
rect 9446 10981 9506 12547
rect 9443 10980 9509 10981
rect 9443 10916 9444 10980
rect 9508 10916 9509 10980
rect 9443 10915 9509 10916
rect 9259 10844 9325 10845
rect 9259 10780 9260 10844
rect 9324 10780 9325 10844
rect 9259 10779 9325 10780
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 8736 8660 9760
rect 9075 9756 9141 9757
rect 9075 9692 9076 9756
rect 9140 9692 9141 9756
rect 9075 9691 9141 9692
rect 8891 8804 8957 8805
rect 8891 8740 8892 8804
rect 8956 8740 8957 8804
rect 8891 8739 8957 8740
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 7648 8660 8672
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 6560 8660 7584
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 5472 8660 6496
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8894 4861 8954 8739
rect 9078 7581 9138 9691
rect 9630 9298 9690 14043
rect 9811 13564 9877 13565
rect 9811 13500 9812 13564
rect 9876 13500 9877 13564
rect 9811 13499 9877 13500
rect 9814 10981 9874 13499
rect 9811 10980 9877 10981
rect 9811 10916 9812 10980
rect 9876 10916 9877 10980
rect 9811 10915 9877 10916
rect 9998 10845 10058 14723
rect 10805 14720 11125 15744
rect 12203 15060 12269 15061
rect 12203 14996 12204 15060
rect 12268 14996 12269 15060
rect 12203 14995 12269 14996
rect 11651 14788 11717 14789
rect 11651 14724 11652 14788
rect 11716 14724 11717 14788
rect 11651 14723 11717 14724
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 13632 11125 14656
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10547 13564 10613 13565
rect 10547 13500 10548 13564
rect 10612 13500 10613 13564
rect 10547 13499 10613 13500
rect 10179 13020 10245 13021
rect 10179 12956 10180 13020
rect 10244 12956 10245 13020
rect 10179 12955 10245 12956
rect 9995 10844 10061 10845
rect 9995 10780 9996 10844
rect 10060 10780 10061 10844
rect 9995 10779 10061 10780
rect 9995 9892 10061 9893
rect 9995 9828 9996 9892
rect 10060 9828 10061 9892
rect 9995 9827 10061 9828
rect 9259 8260 9325 8261
rect 9259 8196 9260 8260
rect 9324 8196 9325 8260
rect 9259 8195 9325 8196
rect 9627 8260 9693 8261
rect 9627 8196 9628 8260
rect 9692 8196 9693 8260
rect 9627 8195 9693 8196
rect 9075 7580 9141 7581
rect 9075 7516 9076 7580
rect 9140 7516 9141 7580
rect 9075 7515 9141 7516
rect 9075 6900 9141 6901
rect 9075 6836 9076 6900
rect 9140 6836 9141 6900
rect 9075 6835 9141 6836
rect 9078 6085 9138 6835
rect 9075 6084 9141 6085
rect 9075 6020 9076 6084
rect 9140 6020 9141 6084
rect 9075 6019 9141 6020
rect 8891 4860 8957 4861
rect 8891 4796 8892 4860
rect 8956 4796 8957 4860
rect 8891 4795 8957 4796
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 3296 8660 4320
rect 9262 4317 9322 8195
rect 9443 7580 9509 7581
rect 9443 7516 9444 7580
rect 9508 7516 9509 7580
rect 9443 7515 9509 7516
rect 9259 4316 9325 4317
rect 8891 4252 8892 4302
rect 8956 4252 8957 4302
rect 8891 4251 8957 4252
rect 9259 4252 9260 4316
rect 9324 4252 9325 4316
rect 9259 4251 9325 4252
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 7787 2684 7853 2685
rect 7787 2620 7788 2684
rect 7852 2620 7853 2684
rect 7787 2619 7853 2620
rect 8155 2684 8221 2685
rect 8155 2620 8156 2684
rect 8220 2620 8221 2684
rect 8155 2619 8221 2620
rect 7603 2412 7669 2413
rect 7603 2348 7604 2412
rect 7668 2348 7669 2412
rect 7603 2347 7669 2348
rect 8340 2208 8660 3232
rect 8891 3228 8957 3229
rect 8891 3164 8892 3228
rect 8956 3164 8957 3228
rect 8891 3163 8957 3164
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 8894 1869 8954 3163
rect 9446 2005 9506 7515
rect 9630 4317 9690 8195
rect 9811 7036 9877 7037
rect 9811 6972 9812 7036
rect 9876 6972 9877 7036
rect 9811 6971 9877 6972
rect 9814 5949 9874 6971
rect 9811 5948 9877 5949
rect 9811 5884 9812 5948
rect 9876 5884 9877 5948
rect 9811 5883 9877 5884
rect 9627 4316 9693 4317
rect 9627 4252 9628 4316
rect 9692 4252 9693 4316
rect 9627 4251 9693 4252
rect 9998 2821 10058 9827
rect 10182 9757 10242 12955
rect 10363 12612 10429 12613
rect 10363 12548 10364 12612
rect 10428 12548 10429 12612
rect 10363 12547 10429 12548
rect 10366 10573 10426 12547
rect 10363 10572 10429 10573
rect 10363 10508 10364 10572
rect 10428 10508 10429 10572
rect 10363 10507 10429 10508
rect 10179 9756 10245 9757
rect 10179 9692 10180 9756
rect 10244 9692 10245 9756
rect 10179 9691 10245 9692
rect 10366 8125 10426 10507
rect 10550 9893 10610 13499
rect 10805 12544 11125 13568
rect 11283 12884 11349 12885
rect 11283 12820 11284 12884
rect 11348 12820 11349 12884
rect 11283 12819 11349 12820
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 11456 11125 12480
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 10368 11125 11392
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10547 9892 10613 9893
rect 10547 9828 10548 9892
rect 10612 9828 10613 9892
rect 10547 9827 10613 9828
rect 10547 9620 10613 9621
rect 10547 9556 10548 9620
rect 10612 9556 10613 9620
rect 10547 9555 10613 9556
rect 10550 9349 10610 9555
rect 10547 9348 10613 9349
rect 10547 9284 10548 9348
rect 10612 9284 10613 9348
rect 10547 9283 10613 9284
rect 10805 9280 11125 10304
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10547 9212 10613 9213
rect 10547 9148 10548 9212
rect 10612 9148 10613 9212
rect 10547 9147 10613 9148
rect 10363 8124 10429 8125
rect 10363 8060 10364 8124
rect 10428 8060 10429 8124
rect 10363 8059 10429 8060
rect 10179 6084 10245 6085
rect 10179 6020 10180 6084
rect 10244 6020 10245 6084
rect 10179 6019 10245 6020
rect 9995 2820 10061 2821
rect 9995 2756 9996 2820
rect 10060 2756 10061 2820
rect 9995 2755 10061 2756
rect 10182 2685 10242 6019
rect 10179 2684 10245 2685
rect 10179 2620 10180 2684
rect 10244 2620 10245 2684
rect 10179 2619 10245 2620
rect 10366 2141 10426 8059
rect 10550 6493 10610 9147
rect 10805 8192 11125 9216
rect 11286 8261 11346 12819
rect 11654 9757 11714 14723
rect 11835 13564 11901 13565
rect 11835 13500 11836 13564
rect 11900 13500 11901 13564
rect 11835 13499 11901 13500
rect 12019 13564 12085 13565
rect 12019 13500 12020 13564
rect 12084 13500 12085 13564
rect 12019 13499 12085 13500
rect 11838 11253 11898 13499
rect 11835 11252 11901 11253
rect 11835 11188 11836 11252
rect 11900 11188 11901 11252
rect 11835 11187 11901 11188
rect 11835 10436 11901 10437
rect 11835 10372 11836 10436
rect 11900 10372 11901 10436
rect 11835 10371 11901 10372
rect 11651 9756 11717 9757
rect 11651 9692 11652 9756
rect 11716 9692 11717 9756
rect 11651 9691 11717 9692
rect 11651 9212 11717 9213
rect 11651 9148 11652 9212
rect 11716 9148 11717 9212
rect 11651 9147 11717 9148
rect 11467 8940 11533 8941
rect 11467 8876 11468 8940
rect 11532 8876 11533 8940
rect 11467 8875 11533 8876
rect 11283 8260 11349 8261
rect 11283 8196 11284 8260
rect 11348 8196 11349 8260
rect 11283 8195 11349 8196
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 7104 11125 8128
rect 11470 7850 11530 8875
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10547 6492 10613 6493
rect 10547 6428 10548 6492
rect 10612 6428 10613 6492
rect 10547 6427 10613 6428
rect 10550 3365 10610 6427
rect 10805 6016 11125 7040
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 3840 11125 4864
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10547 3364 10613 3365
rect 10547 3300 10548 3364
rect 10612 3300 10613 3364
rect 10547 3299 10613 3300
rect 10805 2752 11125 3776
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10363 2140 10429 2141
rect 10363 2076 10364 2140
rect 10428 2076 10429 2140
rect 10805 2128 11125 2688
rect 11286 7790 11530 7850
rect 11286 2685 11346 7790
rect 11467 6084 11533 6085
rect 11467 6020 11468 6084
rect 11532 6020 11533 6084
rect 11467 6019 11533 6020
rect 11470 4997 11530 6019
rect 11467 4996 11533 4997
rect 11467 4932 11468 4996
rect 11532 4932 11533 4996
rect 11467 4931 11533 4932
rect 11654 4861 11714 9147
rect 11838 7853 11898 10371
rect 11835 7852 11901 7853
rect 11835 7788 11836 7852
rect 11900 7788 11901 7852
rect 11835 7787 11901 7788
rect 11835 6220 11901 6221
rect 11835 6156 11836 6220
rect 11900 6156 11901 6220
rect 11835 6155 11901 6156
rect 11651 4860 11717 4861
rect 11651 4858 11652 4860
rect 11470 4798 11652 4858
rect 11283 2684 11349 2685
rect 11283 2620 11284 2684
rect 11348 2620 11349 2684
rect 11283 2619 11349 2620
rect 11470 2546 11530 4798
rect 11651 4796 11652 4798
rect 11716 4796 11717 4860
rect 11651 4795 11717 4796
rect 11838 4589 11898 6155
rect 11835 4588 11901 4589
rect 11835 4524 11836 4588
rect 11900 4524 11901 4588
rect 11835 4523 11901 4524
rect 12022 3501 12082 13499
rect 12206 9213 12266 14995
rect 12390 10845 12450 16083
rect 13270 15264 13590 15824
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13123 14380 13189 14381
rect 13123 14316 13124 14380
rect 13188 14316 13189 14380
rect 13123 14315 13189 14316
rect 12571 13700 12637 13701
rect 12571 13636 12572 13700
rect 12636 13636 12637 13700
rect 12571 13635 12637 13636
rect 12387 10844 12453 10845
rect 12387 10780 12388 10844
rect 12452 10780 12453 10844
rect 12387 10779 12453 10780
rect 12203 9212 12269 9213
rect 12203 9148 12204 9212
rect 12268 9148 12269 9212
rect 12203 9147 12269 9148
rect 12387 9212 12453 9213
rect 12387 9148 12388 9212
rect 12452 9148 12453 9212
rect 12387 9147 12453 9148
rect 12203 8804 12269 8805
rect 12203 8740 12204 8804
rect 12268 8740 12269 8804
rect 12203 8739 12269 8740
rect 12019 3500 12085 3501
rect 12019 3436 12020 3500
rect 12084 3436 12085 3500
rect 12019 3435 12085 3436
rect 12206 3229 12266 8739
rect 12390 5541 12450 9147
rect 12574 5813 12634 13635
rect 12755 9892 12821 9893
rect 12755 9828 12756 9892
rect 12820 9828 12821 9892
rect 12755 9827 12821 9828
rect 12571 5812 12637 5813
rect 12571 5748 12572 5812
rect 12636 5748 12637 5812
rect 12571 5747 12637 5748
rect 12387 5540 12453 5541
rect 12387 5476 12388 5540
rect 12452 5476 12453 5540
rect 12387 5475 12453 5476
rect 12571 5404 12637 5405
rect 12571 5340 12572 5404
rect 12636 5340 12637 5404
rect 12571 5339 12637 5340
rect 12387 4588 12453 4589
rect 12387 4524 12388 4588
rect 12452 4524 12453 4588
rect 12387 4523 12453 4524
rect 12203 3228 12269 3229
rect 12203 3164 12204 3228
rect 12268 3164 12269 3228
rect 12203 3163 12269 3164
rect 11286 2486 11530 2546
rect 10363 2075 10429 2076
rect 9443 2004 9509 2005
rect 9443 1940 9444 2004
rect 9508 1940 9509 2004
rect 9443 1939 9509 1940
rect 8891 1868 8957 1869
rect 8891 1804 8892 1868
rect 8956 1804 8957 1868
rect 8891 1803 8957 1804
rect 11286 1325 11346 2486
rect 12390 1597 12450 4523
rect 12574 2413 12634 5339
rect 12758 4861 12818 9827
rect 12939 7852 13005 7853
rect 12939 7788 12940 7852
rect 13004 7788 13005 7852
rect 12939 7787 13005 7788
rect 12755 4860 12821 4861
rect 12755 4796 12756 4860
rect 12820 4796 12821 4860
rect 12755 4795 12821 4796
rect 12571 2412 12637 2413
rect 12571 2348 12572 2412
rect 12636 2348 12637 2412
rect 12571 2347 12637 2348
rect 12942 2005 13002 7787
rect 13126 2549 13186 14315
rect 13270 14176 13590 15200
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 13088 13590 14112
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 12000 13590 13024
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 10912 13590 11936
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 9824 13590 10848
rect 13859 10436 13925 10437
rect 13859 10372 13860 10436
rect 13924 10372 13925 10436
rect 13859 10371 13925 10372
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 8736 13590 9760
rect 13675 8804 13741 8805
rect 13675 8740 13676 8804
rect 13740 8740 13741 8804
rect 13675 8739 13741 8740
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 7648 13590 8672
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 6560 13590 7584
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 5472 13590 6496
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 3296 13590 4320
rect 13678 3909 13738 8739
rect 13675 3908 13741 3909
rect 13675 3844 13676 3908
rect 13740 3844 13741 3908
rect 13675 3843 13741 3844
rect 13862 3501 13922 10371
rect 14043 9756 14109 9757
rect 14043 9692 14044 9756
rect 14108 9692 14109 9756
rect 14043 9691 14109 9692
rect 13859 3500 13925 3501
rect 13859 3436 13860 3500
rect 13924 3436 13925 3500
rect 13859 3435 13925 3436
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13123 2548 13189 2549
rect 13123 2484 13124 2548
rect 13188 2484 13189 2548
rect 13123 2483 13189 2484
rect 13270 2208 13590 3232
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2128 13590 2144
rect 12939 2004 13005 2005
rect 12939 1940 12940 2004
rect 13004 1940 13005 2004
rect 12939 1939 13005 1940
rect 12387 1596 12453 1597
rect 12387 1532 12388 1596
rect 12452 1532 12453 1596
rect 12387 1531 12453 1532
rect 14046 1461 14106 9691
rect 14043 1460 14109 1461
rect 14043 1396 14044 1460
rect 14108 1396 14109 1460
rect 14043 1395 14109 1396
rect 11283 1324 11349 1325
rect 11283 1260 11284 1324
rect 11348 1260 11349 1324
rect 11283 1259 11349 1260
<< via4 >>
rect 4574 9062 4810 9298
rect 4758 4302 4994 4538
rect 9542 9212 9778 9298
rect 9542 9148 9628 9212
rect 9628 9148 9692 9212
rect 9692 9148 9778 9212
rect 9542 9062 9778 9148
rect 8806 4316 9042 4538
rect 8806 4302 8892 4316
rect 8892 4302 8956 4316
rect 8956 4302 9042 4316
<< metal5 >>
rect 4532 9298 9820 9340
rect 4532 9062 4574 9298
rect 4810 9062 9542 9298
rect 9778 9062 9820 9298
rect 4532 9020 9820 9062
rect 4716 4538 9084 4580
rect 4716 4302 4758 4538
rect 4994 4302 8806 4538
rect 9042 4302 9084 4538
rect 4716 4260 9084 4302
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2116 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2852 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _51_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4324 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1605641404
transform 1 0 6348 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5520 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5796 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1605641404
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7728 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1605641404
transform 1 0 8280 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 9844 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 9476 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90
timestamp 1605641404
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_87
timestamp 1605641404
transform 1 0 9108 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_94
timestamp 1605641404
transform 1 0 9752 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_104
timestamp 1605641404
transform 1 0 10672 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11040 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1605641404
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11776 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1605641404
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1605641404
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1605641404
transform 1 0 13616 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14444 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_134
timestamp 1605641404
transform 1 0 13432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1605641404
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1605641404
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1605641404
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1605641404
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_154
timestamp 1605641404
transform 1 0 15272 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 2852 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 4876 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1605641404
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 5428 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1605641404
transform 1 0 6900 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7728 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1605641404
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1605641404
transform 1 0 10488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10856 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12052 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1605641404
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12880 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13708 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1605641404
transform 1 0 14536 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1605641404
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2852 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 4876 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_3_35 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4324 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1605641404
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1605641404
transform 1 0 8280 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1605641404
transform 1 0 9844 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1605641404
transform 1 0 9476 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_87
timestamp 1605641404
transform 1 0 9108 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_94
timestamp 1605641404
transform 1 0 9752 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_104
timestamp 1605641404
transform 1 0 10672 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 11040 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1605641404
transform 1 0 11868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1605641404
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 13616 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1605641404
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1605641404
transform 1 0 14444 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1605641404
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_153
timestamp 1605641404
transform 1 0 15180 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2852 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1605641404
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5888 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_48
timestamp 1605641404
transform 1 0 5520 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1605641404
transform 1 0 7360 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7728 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1605641404
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1605641404
transform 1 0 10488 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1605641404
transform 1 0 10856 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_115
timestamp 1605641404
transform 1 0 11684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1605641404
transform 1 0 14444 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13248 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp 1605641404
transform 1 0 12880 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1605641404
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1605641404
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1564 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2392 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_20
timestamp 1605641404
transform 1 0 2944 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4876 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 3036 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1605641404
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _29_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1605641404
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7820 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1605641404
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1605641404
transform 1 0 10120 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1605641404
transform 1 0 9292 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1605641404
transform 1 0 10488 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_101
timestamp 1605641404
transform 1 0 10396 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1605641404
transform 1 0 11684 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_111
timestamp 1605641404
transform 1 0 11316 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1605641404
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13616 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1605641404
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1605641404
transform 1 0 14444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1605641404
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_153
timestamp 1605641404
transform 1 0 15180 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1605641404
transform 1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2116 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1564 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 2760 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_14
timestamp 1605641404
transform 1 0 2392 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4876 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4416 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 3036 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1605641404
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1605641404
transform 1 0 4508 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6256 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_52
timestamp 1605641404
transform 1 0 5888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1605641404
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8004 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1605641404
transform 1 0 8372 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6900 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 8096 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_72
timestamp 1605641404
transform 1 0 7728 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_72
timestamp 1605641404
transform 1 0 7728 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1605641404
transform 1 0 9476 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1605641404
transform 1 0 9844 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1605641404
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_94
timestamp 1605641404
transform 1 0 9752 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1605641404
transform 1 0 10120 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1605641404
transform 1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 11500 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1605641404
transform 1 0 11132 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_122
timestamp 1605641404
transform 1 0 12328 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_111
timestamp 1605641404
transform 1 0 11316 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1605641404
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12696 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13892 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13616 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1605641404
transform 1 0 13524 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1605641404
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1605641404
transform 1 0 14444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1605641404
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_148
timestamp 1605641404
transform 1 0 14720 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1605641404
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1605641404
transform 1 0 15180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2116 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1605641404
transform 1 0 1748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1605641404
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1605641404
transform 1 0 4876 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5244 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_61
timestamp 1605641404
transform 1 0 6716 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7084 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 8556 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1605641404
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1605641404
transform 1 0 11500 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1605641404
transform 1 0 11132 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_122
timestamp 1605641404
transform 1 0 12328 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 13892 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12696 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1605641404
transform 1 0 13524 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1605641404
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1605641404
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2208 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 3036 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4876 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_37
timestamp 1605641404
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1605641404
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8648 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_78
timestamp 1605641404
transform 1 0 8280 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1605641404
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1605641404
transform 1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_111
timestamp 1605641404
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1605641404
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1605641404
transform 1 0 13616 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1605641404
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_145
timestamp 1605641404
transform 1 0 14444 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1605641404
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1605641404
transform 1 0 15180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1564 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1605641404
transform 1 0 3588 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1605641404
transform 1 0 3220 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1605641404
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1605641404
transform 1 0 4876 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 5612 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 5244 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_48
timestamp 1605641404
transform 1 0 5520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 7452 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1605641404
transform 1 0 7084 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1605641404
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1605641404
transform 1 0 8924 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1605641404
transform 1 0 11500 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_109
timestamp 1605641404
transform 1 0 11132 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_122
timestamp 1605641404
transform 1 0 12328 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1605641404
transform 1 0 13892 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12696 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1605641404
transform 1 0 13524 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp 1605641404
transform 1 0 14720 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1605641404
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1840 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2668 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1605641404
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4876 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1605641404
transform 1 0 4048 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 3496 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1605641404
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8648 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_78
timestamp 1605641404
transform 1 0 8280 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1605641404
transform 1 0 10488 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_98
timestamp 1605641404
transform 1 0 10120 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1605641404
transform 1 0 11684 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_111
timestamp 1605641404
transform 1 0 11316 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1605641404
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1605641404
transform 1 0 13616 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp 1605641404
transform 1 0 13248 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_145
timestamp 1605641404
transform 1 0 14444 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1605641404
transform 1 0 14812 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1605641404
transform 1 0 15180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2760 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1932 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1605641404
transform 1 0 4324 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1605641404
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_32
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5796 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_12_44
timestamp 1605641404
transform 1 0 5152 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_50
timestamp 1605641404
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7636 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1605641404
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1605641404
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1605641404
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12052 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1605641404
transform 1 0 10856 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_115
timestamp 1605641404
transform 1 0 11684 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14168 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13248 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_128
timestamp 1605641404
transform 1 0 12880 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_138
timestamp 1605641404
transform 1 0 13800 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_148
timestamp 1605641404
transform 1 0 14720 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1605641404
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2760 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 1564 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2300 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 1472 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_14
timestamp 1605641404
transform 1 0 2392 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 3772 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4508 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 3128 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1605641404
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_36
timestamp 1605641404
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5704 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 5244 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_46
timestamp 1605641404
transform 1 0 5336 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7544 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1605641404
transform 1 0 8648 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1605641404
transform 1 0 8280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_66
timestamp 1605641404
transform 1 0 7176 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1605641404
transform 1 0 9844 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 1605641404
transform 1 0 9476 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_104
timestamp 1605641404
transform 1 0 10672 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_86
timestamp 1605641404
transform 1 0 9016 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1605641404
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12052 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1605641404
transform 1 0 11040 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10856 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_117
timestamp 1605641404
transform 1 0 11868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1605641404
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_115
timestamp 1605641404
transform 1 0 11684 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1605641404
transform 1 0 14444 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13616 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1605641404
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1605641404
transform 1 0 14444 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_128
timestamp 1605641404
transform 1 0 12880 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1605641404
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1605641404
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1605641404
transform 1 0 15180 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1605641404
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2208 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 4876 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 3036 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_37
timestamp 1605641404
transform 1 0 4508 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1605641404
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1605641404
transform 1 0 8648 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp 1605641404
transform 1 0 8280 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1605641404
transform 1 0 9844 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_91
timestamp 1605641404
transform 1 0 9476 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_104
timestamp 1605641404
transform 1 0 10672 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1605641404
transform 1 0 11040 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_117
timestamp 1605641404
transform 1 0 11868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1605641404
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13616 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1605641404
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_142
timestamp 1605641404
transform 1 0 14168 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14536 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1605641404
transform 1 0 15088 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_156
timestamp 1605641404
transform 1 0 15456 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2760 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1564 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_14
timestamp 1605641404
transform 1 0 2392 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4324 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1605641404
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_32
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5520 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_44
timestamp 1605641404
transform 1 0 5152 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7360 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_64
timestamp 1605641404
transform 1 0 6992 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 9200 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_84
timestamp 1605641404
transform 1 0 8832 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1605641404
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_102
timestamp 1605641404
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10856 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12052 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_115
timestamp 1605641404
transform 1 0 11684 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1605641404
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13248 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_128
timestamp 1605641404
transform 1 0 12880 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1605641404
transform 1 0 14076 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1605641404
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1605641404
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1605641404
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_17
timestamp 1605641404
transform 1 0 2668 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 3036 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4876 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_37
timestamp 1605641404
transform 1 0 4508 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1605641404
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1605641404
transform 1 0 8648 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_78
timestamp 1605641404
transform 1 0 8280 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1605641404
transform 1 0 10580 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1605641404
transform 1 0 9384 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_86
timestamp 1605641404
transform 1 0 9016 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_99
timestamp 1605641404
transform 1 0 10212 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1605641404
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 11868 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_106
timestamp 1605641404
transform 1 0 10856 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1605641404
transform 1 0 11500 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1605641404
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1605641404
transform 1 0 14352 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1605641404
transform 1 0 13616 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1605641404
transform 1 0 13248 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_140
timestamp 1605641404
transform 1 0 13984 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_148
timestamp 1605641404
transform 1 0 14720 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_156
timestamp 1605641404
transform 1 0 15456 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2760 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1564 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1605641404
transform 1 0 2392 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4692 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1605641404
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_35
timestamp 1605641404
transform 1 0 4324 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6532 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_55
timestamp 1605641404
transform 1 0 6164 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1605641404
transform 1 0 8372 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_75
timestamp 1605641404
transform 1 0 8004 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1605641404
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12052 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1605641404
transform 1 0 11500 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1605641404
transform 1 0 11132 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_116
timestamp 1605641404
transform 1 0 11776 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14168 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13248 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_128
timestamp 1605641404
transform 1 0 12880 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_138
timestamp 1605641404
transform 1 0 13800 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1605641404
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1605641404
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2116 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1605641404
transform 1 0 1932 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_18
timestamp 1605641404
transform 1 0 2760 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_7
timestamp 1605641404
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1605641404
transform 1 0 4324 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1605641404
transform 1 0 4324 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1605641404
transform 1 0 3128 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_31
timestamp 1605641404
transform 1 0 3956 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1605641404
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_38
timestamp 1605641404
transform 1 0 4600 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4968 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6808 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1605641404
transform 1 0 5520 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_44
timestamp 1605641404
transform 1 0 5152 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1605641404
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1605641404
transform 1 0 6440 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7728 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1605641404
transform 1 0 8372 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1605641404
transform 1 0 8004 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_68
timestamp 1605641404
transform 1 0 7360 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_81
timestamp 1605641404
transform 1 0 8556 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_71
timestamp 1605641404
transform 1 0 7636 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_78
timestamp 1605641404
transform 1 0 8280 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1605641404
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1605641404
transform 1 0 8924 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1605641404
transform 1 0 10028 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_101
timestamp 1605641404
transform 1 0 10396 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_94
timestamp 1605641404
transform 1 0 9752 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1605641404
transform 1 0 9752 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1605641404
transform 1 0 10120 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10396 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1605641404
transform 1 0 12236 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_114
timestamp 1605641404
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_117
timestamp 1605641404
transform 1 0 11868 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_124
timestamp 1605641404
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13616 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1605641404
transform 1 0 13892 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12696 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1605641404
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1605641404
transform 1 0 14444 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1605641404
transform 1 0 13524 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1605641404
transform 1 0 14812 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1605641404
transform 1 0 15180 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1605641404
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1605641404
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1605641404
transform 1 0 2300 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1605641404
transform 1 0 1564 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_9
timestamp 1605641404
transform 1 0 1932 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_17
timestamp 1605641404
transform 1 0 2668 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1605641404
transform 1 0 3496 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1605641404
transform 1 0 4140 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 3220 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_29
timestamp 1605641404
transform 1 0 3772 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1605641404
transform 1 0 5336 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_42
timestamp 1605641404
transform 1 0 4968 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_55
timestamp 1605641404
transform 1 0 6164 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8464 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1605641404
transform 1 0 7268 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_66
timestamp 1605641404
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_76
timestamp 1605641404
transform 1 0 8096 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10304 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1605641404
transform 1 0 9936 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1605641404
transform 1 0 11500 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_109
timestamp 1605641404
transform 1 0 11132 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_116
timestamp 1605641404
transform 1 0 11776 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13616 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1605641404
transform 1 0 13248 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_145
timestamp 1605641404
transform 1 0 14444 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1605641404
transform 1 0 14812 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1605641404
transform 1 0 15180 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1605641404
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2484 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_11
timestamp 1605641404
transform 1 0 2116 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4324 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1605641404
transform 1 0 3496 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_21
timestamp 1605641404
transform 1 0 3036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_25
timestamp 1605641404
transform 1 0 3404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1605641404
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_32
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6164 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_51
timestamp 1605641404
transform 1 0 5796 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7360 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 8556 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_64
timestamp 1605641404
transform 1 0 6992 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_77
timestamp 1605641404
transform 1 0 8188 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 1605641404
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1605641404
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12052 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_109
timestamp 1605641404
transform 1 0 11132 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_117
timestamp 1605641404
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1605641404
transform 1 0 14168 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13248 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_128
timestamp 1605641404
transform 1 0 12880 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_138
timestamp 1605641404
transform 1 0 13800 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_146
timestamp 1605641404
transform 1 0 14536 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1605641404
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1605641404
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1605641404
transform 1 0 1472 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1605641404
transform 1 0 2760 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1605641404
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_8
timestamp 1605641404
transform 1 0 1840 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_16
timestamp 1605641404
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1605641404
transform 1 0 3588 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4784 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_22
timestamp 1605641404
transform 1 0 3128 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_26
timestamp 1605641404
transform 1 0 3496 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_36
timestamp 1605641404
transform 1 0 4416 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1605641404
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1605641404
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_49
timestamp 1605641404
transform 1 0 5612 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1605641404
transform 1 0 6348 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1605641404
transform 1 0 7820 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1605641404
transform 1 0 8556 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_23_66
timestamp 1605641404
transform 1 0 7176 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_72
timestamp 1605641404
transform 1 0 7728 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_77
timestamp 1605641404
transform 1 0 8188 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1605641404
transform 1 0 9752 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_90
timestamp 1605641404
transform 1 0 9384 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_98
timestamp 1605641404
transform 1 0 10120 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1605641404
transform 1 0 11040 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_106
timestamp 1605641404
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1605641404
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1605641404
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1605641404
transform 1 0 13616 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1605641404
transform 1 0 14352 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_132
timestamp 1605641404
transform 1 0 13248 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 1605641404
transform 1 0 13984 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_148
timestamp 1605641404
transform 1 0 14720 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_156
timestamp 1605641404
transform 1 0 15456 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1605641404
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 2116 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_7
timestamp 1605641404
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1605641404
transform 1 0 4324 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1605641404
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_32
timestamp 1605641404
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1605641404
transform 1 0 5520 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 6808 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_44
timestamp 1605641404
transform 1 0 5152 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_52
timestamp 1605641404
transform 1 0 5888 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_60
timestamp 1605641404
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1605641404
transform 1 0 6900 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8096 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_72
timestamp 1605641404
transform 1 0 7728 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1605641404
transform 1 0 9752 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 9660 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1605641404
transform 1 0 8924 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_98
timestamp 1605641404
transform 1 0 10120 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12604 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1605641404
transform 1 0 10948 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 12512 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_106
timestamp 1605641404
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_116
timestamp 1605641404
transform 1 0 11776 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1605641404
transform 1 0 14260 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1605641404
transform 1 0 13524 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1605641404
transform 1 0 13156 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_139
timestamp 1605641404
transform 1 0 13892 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 15364 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_147
timestamp 1605641404
transform 1 0 14628 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_156
timestamp 1605641404
transform 1 0 15456 0 -1 15776
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 416 480 536 6 ccff_head
port 0 nsew default input
rlabel metal3 s 16520 13472 17000 13592 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 12898 0 12954 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 13818 0 13874 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 16302 0 16358 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 16762 0 16818 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 11242 0 11298 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 12070 0 12126 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 4434 0 4490 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 7010 0 7066 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 1030 0 1086 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 1858 0 1914 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 2686 0 2742 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 3146 0 3202 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 3606 0 3662 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 3974 0 4030 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 8666 17520 8722 18000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 12898 17520 12954 18000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 13358 17520 13414 18000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 13818 17520 13874 18000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 14186 17520 14242 18000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 14646 17520 14702 18000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 15014 17520 15070 18000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 15474 17520 15530 18000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 15934 17520 15990 18000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 16302 17520 16358 18000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 16762 17520 16818 18000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 9126 17520 9182 18000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 9494 17520 9550 18000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 9954 17520 10010 18000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 10414 17520 10470 18000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 10782 17520 10838 18000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 11242 17520 11298 18000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 11610 17520 11666 18000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 12070 17520 12126 18000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 12530 17520 12586 18000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 202 17520 258 18000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 4434 17520 4490 18000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 4802 17520 4858 18000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 5262 17520 5318 18000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 5722 17520 5778 18000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 6090 17520 6146 18000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 6550 17520 6606 18000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 7010 17520 7066 18000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 7378 17520 7434 18000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 7838 17520 7894 18000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 8206 17520 8262 18000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 570 17520 626 18000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 1030 17520 1086 18000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 1398 17520 1454 18000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 1858 17520 1914 18000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 2318 17520 2374 18000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 2686 17520 2742 18000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 3146 17520 3202 18000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 3606 17520 3662 18000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 3974 17520 4030 18000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 left_grid_pin_16_
port 82 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 left_grid_pin_17_
port 83 nsew default tristate
rlabel metal3 s 0 3544 480 3664 6 left_grid_pin_18_
port 84 nsew default tristate
rlabel metal3 s 0 4632 480 4752 6 left_grid_pin_19_
port 85 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 left_grid_pin_20_
port 86 nsew default tristate
rlabel metal3 s 0 6672 480 6792 6 left_grid_pin_21_
port 87 nsew default tristate
rlabel metal3 s 0 7760 480 7880 6 left_grid_pin_22_
port 88 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 left_grid_pin_23_
port 89 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 left_grid_pin_24_
port 90 nsew default tristate
rlabel metal3 s 0 10888 480 11008 6 left_grid_pin_25_
port 91 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 left_grid_pin_26_
port 92 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 left_grid_pin_27_
port 93 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 left_grid_pin_28_
port 94 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 left_grid_pin_29_
port 95 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 left_grid_pin_30_
port 96 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 left_grid_pin_31_
port 97 nsew default tristate
rlabel metal3 s 16520 4496 17000 4616 6 prog_clk
port 98 nsew default input
rlabel metal4 s 3409 2128 3729 15824 6 VPWR
port 99 nsew default input
rlabel metal4 s 5875 2128 6195 15824 6 VGND
port 100 nsew default input
<< properties >>
string FIXED_BBOX 0 0 17000 18000
<< end >>
