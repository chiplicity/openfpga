magic
tech sky130A
magscale 1 2
timestamp 1606928950
<< locali >>
rect 7573 7191 7607 7293
<< viali >>
rect 3985 15113 4019 15147
rect 4721 15113 4755 15147
rect 5549 15113 5583 15147
rect 7297 15113 7331 15147
rect 9505 15113 9539 15147
rect 3801 14909 3835 14943
rect 4537 14909 4571 14943
rect 5365 14909 5399 14943
rect 7113 14909 7147 14943
rect 9321 14909 9355 14943
rect 5733 13957 5767 13991
rect 4353 13821 4387 13855
rect 4609 13821 4643 13855
rect 4905 13481 4939 13515
rect 14841 13481 14875 13515
rect 2881 13345 2915 13379
rect 3249 13345 3283 13379
rect 5089 13345 5123 13379
rect 14657 13345 14691 13379
rect 3341 13141 3375 13175
rect 7389 12801 7423 12835
rect 7297 12733 7331 12767
rect 7205 12665 7239 12699
rect 6837 12597 6871 12631
rect 6101 12325 6135 12359
rect 8309 12257 8343 12291
rect 8401 12189 8435 12223
rect 8493 12189 8527 12223
rect 7389 12053 7423 12087
rect 7941 12053 7975 12087
rect 9229 11849 9263 11883
rect 7389 11713 7423 11747
rect 7205 11645 7239 11679
rect 7849 11645 7883 11679
rect 8094 11577 8128 11611
rect 6837 11509 6871 11543
rect 7297 11509 7331 11543
rect 6745 11305 6779 11339
rect 6653 11237 6687 11271
rect 7542 11237 7576 11271
rect 7297 11169 7331 11203
rect 10057 11169 10091 11203
rect 6929 11101 6963 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 6285 11033 6319 11067
rect 8677 10965 8711 10999
rect 9689 10965 9723 10999
rect 7389 10693 7423 10727
rect 9045 10693 9079 10727
rect 4077 10625 4111 10659
rect 5089 10625 5123 10659
rect 7665 10625 7699 10659
rect 9781 10625 9815 10659
rect 9873 10625 9907 10659
rect 10885 10625 10919 10659
rect 3224 10557 3258 10591
rect 7573 10557 7607 10591
rect 10793 10557 10827 10591
rect 4169 10489 4203 10523
rect 7932 10489 7966 10523
rect 9689 10489 9723 10523
rect 3295 10421 3329 10455
rect 9321 10421 9355 10455
rect 10333 10421 10367 10455
rect 10701 10421 10735 10455
rect 6653 10217 6687 10251
rect 9689 10217 9723 10251
rect 1593 10149 1627 10183
rect 2513 10149 2547 10183
rect 7564 10149 7598 10183
rect 6745 10081 6779 10115
rect 7297 10081 7331 10115
rect 1501 10013 1535 10047
rect 6929 10013 6963 10047
rect 6285 9877 6319 9911
rect 8677 9877 8711 9911
rect 7757 9537 7791 9571
rect 7849 9537 7883 9571
rect 8769 9537 8803 9571
rect 8861 9537 8895 9571
rect 7665 9401 7699 9435
rect 7297 9333 7331 9367
rect 8309 9333 8343 9367
rect 8677 9333 8711 9367
rect 12541 8993 12575 9027
rect 12725 8925 12759 8959
rect 7205 8041 7239 8075
rect 7021 7905 7055 7939
rect 5089 7497 5123 7531
rect 6377 7497 6411 7531
rect 7389 7497 7423 7531
rect 9689 7497 9723 7531
rect 10425 7497 10459 7531
rect 10977 7497 11011 7531
rect 11805 7497 11839 7531
rect 12633 7497 12667 7531
rect 7941 7429 7975 7463
rect 3249 7293 3283 7327
rect 4905 7293 4939 7327
rect 5641 7293 5675 7327
rect 6193 7293 6227 7327
rect 7205 7293 7239 7327
rect 7573 7293 7607 7327
rect 7757 7293 7791 7327
rect 8309 7293 8343 7327
rect 8953 7293 8987 7327
rect 9505 7293 9539 7327
rect 10241 7293 10275 7327
rect 10793 7293 10827 7327
rect 11621 7293 11655 7327
rect 12449 7293 12483 7327
rect 3525 7225 3559 7259
rect 5825 7157 5859 7191
rect 7573 7157 7607 7191
rect 8493 7157 8527 7191
rect 9137 7157 9171 7191
rect 4813 6817 4847 6851
rect 5641 6817 5675 6851
rect 6285 6817 6319 6851
rect 6837 6817 6871 6851
rect 7389 6817 7423 6851
rect 7941 6817 7975 6851
rect 8493 6817 8527 6851
rect 9045 6817 9079 6851
rect 9965 6817 9999 6851
rect 10701 6817 10735 6851
rect 11437 6817 11471 6851
rect 11989 6817 12023 6851
rect 12541 6817 12575 6851
rect 6469 6681 6503 6715
rect 7021 6681 7055 6715
rect 10149 6681 10183 6715
rect 12173 6681 12207 6715
rect 4997 6613 5031 6647
rect 5825 6613 5859 6647
rect 7573 6613 7607 6647
rect 8125 6613 8159 6647
rect 8677 6613 8711 6647
rect 9229 6613 9263 6647
rect 10885 6613 10919 6647
rect 11621 6613 11655 6647
rect 12725 6613 12759 6647
rect 7941 6341 7975 6375
rect 9597 6341 9631 6375
rect 3709 6205 3743 6239
rect 4353 6205 4387 6239
rect 5181 6205 5215 6239
rect 7757 6205 7791 6239
rect 9413 6205 9447 6239
rect 10241 6205 10275 6239
rect 11529 6205 11563 6239
rect 3893 6069 3927 6103
rect 4537 6069 4571 6103
rect 5365 6069 5399 6103
rect 10425 6069 10459 6103
rect 11713 6069 11747 6103
rect 7573 5729 7607 5763
rect 9689 5729 9723 5763
rect 9873 5593 9907 5627
rect 7757 5525 7791 5559
<< metal1 >>
rect 1104 17434 15824 17456
rect 1104 17382 3447 17434
rect 3499 17382 3511 17434
rect 3563 17382 3575 17434
rect 3627 17382 3639 17434
rect 3691 17382 8378 17434
rect 8430 17382 8442 17434
rect 8494 17382 8506 17434
rect 8558 17382 8570 17434
rect 8622 17382 13308 17434
rect 13360 17382 13372 17434
rect 13424 17382 13436 17434
rect 13488 17382 13500 17434
rect 13552 17382 15824 17434
rect 1104 17360 15824 17382
rect 9766 17008 9772 17060
rect 9824 17048 9830 17060
rect 10962 17048 10968 17060
rect 9824 17020 10968 17048
rect 9824 17008 9830 17020
rect 10962 17008 10968 17020
rect 11020 17008 11026 17060
rect 1104 16890 15824 16912
rect 1104 16838 5912 16890
rect 5964 16838 5976 16890
rect 6028 16838 6040 16890
rect 6092 16838 6104 16890
rect 6156 16838 10843 16890
rect 10895 16838 10907 16890
rect 10959 16838 10971 16890
rect 11023 16838 11035 16890
rect 11087 16838 15824 16890
rect 1104 16816 15824 16838
rect 4798 16396 4804 16448
rect 4856 16436 4862 16448
rect 9306 16436 9312 16448
rect 4856 16408 9312 16436
rect 4856 16396 4862 16408
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 1104 16346 15824 16368
rect 1104 16294 3447 16346
rect 3499 16294 3511 16346
rect 3563 16294 3575 16346
rect 3627 16294 3639 16346
rect 3691 16294 8378 16346
rect 8430 16294 8442 16346
rect 8494 16294 8506 16346
rect 8558 16294 8570 16346
rect 8622 16294 13308 16346
rect 13360 16294 13372 16346
rect 13424 16294 13436 16346
rect 13488 16294 13500 16346
rect 13552 16294 15824 16346
rect 1104 16272 15824 16294
rect 3050 16192 3056 16244
rect 3108 16232 3114 16244
rect 6454 16232 6460 16244
rect 3108 16204 6460 16232
rect 3108 16192 3114 16204
rect 6454 16192 6460 16204
rect 6512 16192 6518 16244
rect 9122 16192 9128 16244
rect 9180 16232 9186 16244
rect 11330 16232 11336 16244
rect 9180 16204 11336 16232
rect 9180 16192 9186 16204
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 5534 16124 5540 16176
rect 5592 16164 5598 16176
rect 8202 16164 8208 16176
rect 5592 16136 8208 16164
rect 5592 16124 5598 16136
rect 8202 16124 8208 16136
rect 8260 16124 8266 16176
rect 6362 16056 6368 16108
rect 6420 16096 6426 16108
rect 8110 16096 8116 16108
rect 6420 16068 8116 16096
rect 6420 16056 6426 16068
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 3878 15988 3884 16040
rect 3936 16028 3942 16040
rect 5626 16028 5632 16040
rect 3936 16000 5632 16028
rect 3936 15988 3942 16000
rect 5626 15988 5632 16000
rect 5684 15988 5690 16040
rect 6822 15988 6828 16040
rect 6880 16028 6886 16040
rect 7834 16028 7840 16040
rect 6880 16000 7840 16028
rect 6880 15988 6886 16000
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 8662 15988 8668 16040
rect 8720 16028 8726 16040
rect 9582 16028 9588 16040
rect 8720 16000 9588 16028
rect 8720 15988 8726 16000
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 14550 15988 14556 16040
rect 14608 16028 14614 16040
rect 16298 16028 16304 16040
rect 14608 16000 16304 16028
rect 14608 15988 14614 16000
rect 16298 15988 16304 16000
rect 16356 15988 16362 16040
rect 3326 15920 3332 15972
rect 3384 15960 3390 15972
rect 6362 15960 6368 15972
rect 3384 15932 6368 15960
rect 3384 15920 3390 15932
rect 6362 15920 6368 15932
rect 6420 15920 6426 15972
rect 7926 15920 7932 15972
rect 7984 15960 7990 15972
rect 12618 15960 12624 15972
rect 7984 15932 12624 15960
rect 7984 15920 7990 15932
rect 12618 15920 12624 15932
rect 12676 15920 12682 15972
rect 4706 15852 4712 15904
rect 4764 15892 4770 15904
rect 6822 15892 6828 15904
rect 4764 15864 6828 15892
rect 4764 15852 4770 15864
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 8018 15852 8024 15904
rect 8076 15892 8082 15904
rect 12158 15892 12164 15904
rect 8076 15864 12164 15892
rect 8076 15852 8082 15864
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 1104 15802 15824 15824
rect 1104 15750 5912 15802
rect 5964 15750 5976 15802
rect 6028 15750 6040 15802
rect 6092 15750 6104 15802
rect 6156 15750 10843 15802
rect 10895 15750 10907 15802
rect 10959 15750 10971 15802
rect 11023 15750 11035 15802
rect 11087 15750 15824 15802
rect 1104 15728 15824 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 4706 15688 4712 15700
rect 1452 15660 4712 15688
rect 1452 15648 1458 15660
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 6270 15648 6276 15700
rect 6328 15688 6334 15700
rect 10042 15688 10048 15700
rect 6328 15660 10048 15688
rect 6328 15648 6334 15660
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 9398 15580 9404 15632
rect 9456 15620 9462 15632
rect 14274 15620 14280 15632
rect 9456 15592 14280 15620
rect 9456 15580 9462 15592
rect 14274 15580 14280 15592
rect 14332 15580 14338 15632
rect 1026 15444 1032 15496
rect 1084 15484 1090 15496
rect 5074 15484 5080 15496
rect 1084 15456 5080 15484
rect 1084 15444 1090 15456
rect 5074 15444 5080 15456
rect 5132 15444 5138 15496
rect 9306 15444 9312 15496
rect 9364 15484 9370 15496
rect 13170 15484 13176 15496
rect 9364 15456 13176 15484
rect 9364 15444 9370 15456
rect 13170 15444 13176 15456
rect 13228 15444 13234 15496
rect 14366 15444 14372 15496
rect 14424 15484 14430 15496
rect 15930 15484 15936 15496
rect 14424 15456 15936 15484
rect 14424 15444 14430 15456
rect 15930 15444 15936 15456
rect 15988 15444 15994 15496
rect 2222 15376 2228 15428
rect 2280 15416 2286 15428
rect 5534 15416 5540 15428
rect 2280 15388 5540 15416
rect 2280 15376 2286 15388
rect 5534 15376 5540 15388
rect 5592 15376 5598 15428
rect 7006 15376 7012 15428
rect 7064 15416 7070 15428
rect 9674 15416 9680 15428
rect 7064 15388 9680 15416
rect 7064 15376 7070 15388
rect 9674 15376 9680 15388
rect 9732 15376 9738 15428
rect 198 15308 204 15360
rect 256 15348 262 15360
rect 2866 15348 2872 15360
rect 256 15320 2872 15348
rect 256 15308 262 15320
rect 2866 15308 2872 15320
rect 2924 15308 2930 15360
rect 7190 15308 7196 15360
rect 7248 15348 7254 15360
rect 9490 15348 9496 15360
rect 7248 15320 9496 15348
rect 7248 15308 7254 15320
rect 9490 15308 9496 15320
rect 9548 15308 9554 15360
rect 1104 15258 15824 15280
rect 1104 15206 3447 15258
rect 3499 15206 3511 15258
rect 3563 15206 3575 15258
rect 3627 15206 3639 15258
rect 3691 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 13308 15258
rect 13360 15206 13372 15258
rect 13424 15206 13436 15258
rect 13488 15206 13500 15258
rect 13552 15206 15824 15258
rect 1104 15184 15824 15206
rect 566 15104 572 15156
rect 624 15144 630 15156
rect 3973 15147 4031 15153
rect 3973 15144 3985 15147
rect 624 15116 3985 15144
rect 624 15104 630 15116
rect 3973 15113 3985 15116
rect 4019 15113 4031 15147
rect 4706 15144 4712 15156
rect 4667 15116 4712 15144
rect 3973 15107 4031 15113
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 5534 15144 5540 15156
rect 5495 15116 5540 15144
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 6822 15104 6828 15156
rect 6880 15144 6886 15156
rect 7285 15147 7343 15153
rect 7285 15144 7297 15147
rect 6880 15116 7297 15144
rect 6880 15104 6886 15116
rect 7285 15113 7297 15116
rect 7331 15113 7343 15147
rect 9490 15144 9496 15156
rect 9451 15116 9496 15144
rect 7285 15107 7343 15113
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 6730 15008 6736 15020
rect 4540 14980 6736 15008
rect 4540 14949 4568 14980
rect 6730 14968 6736 14980
rect 6788 14968 6794 15020
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14909 4583 14943
rect 4525 14903 4583 14909
rect 5353 14943 5411 14949
rect 5353 14909 5365 14943
rect 5399 14940 5411 14943
rect 7101 14943 7159 14949
rect 5399 14912 7052 14940
rect 5399 14909 5411 14912
rect 5353 14903 5411 14909
rect 3804 14872 3832 14903
rect 6546 14872 6552 14884
rect 3804 14844 6552 14872
rect 6546 14832 6552 14844
rect 6604 14832 6610 14884
rect 7024 14872 7052 14912
rect 7101 14909 7113 14943
rect 7147 14940 7159 14943
rect 8938 14940 8944 14952
rect 7147 14912 8944 14940
rect 7147 14909 7159 14912
rect 7101 14903 7159 14909
rect 8938 14900 8944 14912
rect 8996 14900 9002 14952
rect 9309 14943 9367 14949
rect 9309 14909 9321 14943
rect 9355 14940 9367 14943
rect 9858 14940 9864 14952
rect 9355 14912 9864 14940
rect 9355 14909 9367 14912
rect 9309 14903 9367 14909
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 8018 14872 8024 14884
rect 7024 14844 8024 14872
rect 8018 14832 8024 14844
rect 8076 14832 8082 14884
rect 1104 14714 15824 14736
rect 1104 14662 5912 14714
rect 5964 14662 5976 14714
rect 6028 14662 6040 14714
rect 6092 14662 6104 14714
rect 6156 14662 10843 14714
rect 10895 14662 10907 14714
rect 10959 14662 10971 14714
rect 11023 14662 11035 14714
rect 11087 14662 15824 14714
rect 1104 14640 15824 14662
rect 1104 14170 15824 14192
rect 1104 14118 3447 14170
rect 3499 14118 3511 14170
rect 3563 14118 3575 14170
rect 3627 14118 3639 14170
rect 3691 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 13308 14170
rect 13360 14118 13372 14170
rect 13424 14118 13436 14170
rect 13488 14118 13500 14170
rect 13552 14118 15824 14170
rect 1104 14096 15824 14118
rect 5721 13991 5779 13997
rect 5721 13957 5733 13991
rect 5767 13988 5779 13991
rect 7374 13988 7380 14000
rect 5767 13960 7380 13988
rect 5767 13957 5779 13960
rect 5721 13951 5779 13957
rect 7374 13948 7380 13960
rect 7432 13948 7438 14000
rect 3786 13880 3792 13932
rect 3844 13920 3850 13932
rect 3844 13892 4476 13920
rect 3844 13880 3850 13892
rect 4338 13852 4344 13864
rect 4299 13824 4344 13852
rect 4338 13812 4344 13824
rect 4396 13812 4402 13864
rect 4448 13852 4476 13892
rect 4597 13855 4655 13861
rect 4597 13852 4609 13855
rect 4448 13824 4609 13852
rect 4597 13821 4609 13824
rect 4643 13821 4655 13855
rect 4597 13815 4655 13821
rect 1104 13626 15824 13648
rect 1104 13574 5912 13626
rect 5964 13574 5976 13626
rect 6028 13574 6040 13626
rect 6092 13574 6104 13626
rect 6156 13574 10843 13626
rect 10895 13574 10907 13626
rect 10959 13574 10971 13626
rect 11023 13574 11035 13626
rect 11087 13574 15824 13626
rect 1104 13552 15824 13574
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 4893 13515 4951 13521
rect 4893 13512 4905 13515
rect 4396 13484 4905 13512
rect 4396 13472 4402 13484
rect 4893 13481 4905 13484
rect 4939 13481 4951 13515
rect 4893 13475 4951 13481
rect 13722 13472 13728 13524
rect 13780 13512 13786 13524
rect 14829 13515 14887 13521
rect 14829 13512 14841 13515
rect 13780 13484 14841 13512
rect 13780 13472 13786 13484
rect 14829 13481 14841 13484
rect 14875 13481 14887 13515
rect 14829 13475 14887 13481
rect 2866 13376 2872 13388
rect 2827 13348 2872 13376
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 3237 13379 3295 13385
rect 3237 13345 3249 13379
rect 3283 13345 3295 13379
rect 3237 13339 3295 13345
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13376 5135 13379
rect 7190 13376 7196 13388
rect 5123 13348 7196 13376
rect 5123 13345 5135 13348
rect 5077 13339 5135 13345
rect 3252 13308 3280 13339
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 14645 13379 14703 13385
rect 14645 13376 14657 13379
rect 13832 13348 14657 13376
rect 9214 13308 9220 13320
rect 3252 13280 9220 13308
rect 9214 13268 9220 13280
rect 9272 13268 9278 13320
rect 13832 13184 13860 13348
rect 14645 13345 14657 13348
rect 14691 13345 14703 13379
rect 14645 13339 14703 13345
rect 3326 13172 3332 13184
rect 3287 13144 3332 13172
rect 3326 13132 3332 13144
rect 3384 13132 3390 13184
rect 13814 13132 13820 13184
rect 13872 13132 13878 13184
rect 1104 13082 15824 13104
rect 1104 13030 3447 13082
rect 3499 13030 3511 13082
rect 3563 13030 3575 13082
rect 3627 13030 3639 13082
rect 3691 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 13308 13082
rect 13360 13030 13372 13082
rect 13424 13030 13436 13082
rect 13488 13030 13500 13082
rect 13552 13030 15824 13082
rect 1104 13008 15824 13030
rect 7374 12832 7380 12844
rect 7335 12804 7380 12832
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 6730 12724 6736 12776
rect 6788 12764 6794 12776
rect 6914 12764 6920 12776
rect 6788 12736 6920 12764
rect 6788 12724 6794 12736
rect 6914 12724 6920 12736
rect 6972 12764 6978 12776
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 6972 12736 7297 12764
rect 6972 12724 6978 12736
rect 7285 12733 7297 12736
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 7006 12656 7012 12708
rect 7064 12696 7070 12708
rect 7193 12699 7251 12705
rect 7193 12696 7205 12699
rect 7064 12668 7205 12696
rect 7064 12656 7070 12668
rect 7193 12665 7205 12668
rect 7239 12665 7251 12699
rect 7193 12659 7251 12665
rect 6270 12588 6276 12640
rect 6328 12628 6334 12640
rect 6825 12631 6883 12637
rect 6825 12628 6837 12631
rect 6328 12600 6837 12628
rect 6328 12588 6334 12600
rect 6825 12597 6837 12600
rect 6871 12597 6883 12631
rect 6825 12591 6883 12597
rect 9214 12588 9220 12640
rect 9272 12628 9278 12640
rect 13722 12628 13728 12640
rect 9272 12600 13728 12628
rect 9272 12588 9278 12600
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 1104 12538 15824 12560
rect 1104 12486 5912 12538
rect 5964 12486 5976 12538
rect 6028 12486 6040 12538
rect 6092 12486 6104 12538
rect 6156 12486 10843 12538
rect 10895 12486 10907 12538
rect 10959 12486 10971 12538
rect 11023 12486 11035 12538
rect 11087 12486 15824 12538
rect 1104 12464 15824 12486
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 8846 12424 8852 12436
rect 6696 12396 8852 12424
rect 6696 12384 6702 12396
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 6089 12359 6147 12365
rect 6089 12325 6101 12359
rect 6135 12356 6147 12359
rect 11146 12356 11152 12368
rect 6135 12328 11152 12356
rect 6135 12325 6147 12328
rect 6089 12319 6147 12325
rect 11146 12316 11152 12328
rect 11204 12316 11210 12368
rect 8297 12291 8355 12297
rect 8297 12257 8309 12291
rect 8343 12288 8355 12291
rect 9858 12288 9864 12300
rect 8343 12260 9864 12288
rect 8343 12257 8355 12260
rect 8297 12251 8355 12257
rect 9858 12248 9864 12260
rect 9916 12288 9922 12300
rect 10502 12288 10508 12300
rect 9916 12260 10508 12288
rect 9916 12248 9922 12260
rect 10502 12248 10508 12260
rect 10560 12248 10566 12300
rect 8018 12180 8024 12232
rect 8076 12220 8082 12232
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 8076 12192 8401 12220
rect 8076 12180 8082 12192
rect 8389 12189 8401 12192
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 7282 12112 7288 12164
rect 7340 12152 7346 12164
rect 8496 12152 8524 12183
rect 7340 12124 8524 12152
rect 7340 12112 7346 12124
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 7377 12087 7435 12093
rect 7377 12084 7389 12087
rect 7248 12056 7389 12084
rect 7248 12044 7254 12056
rect 7377 12053 7389 12056
rect 7423 12053 7435 12087
rect 7377 12047 7435 12053
rect 7929 12087 7987 12093
rect 7929 12053 7941 12087
rect 7975 12084 7987 12087
rect 8754 12084 8760 12096
rect 7975 12056 8760 12084
rect 7975 12053 7987 12056
rect 7929 12047 7987 12053
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 1104 11994 15824 12016
rect 1104 11942 3447 11994
rect 3499 11942 3511 11994
rect 3563 11942 3575 11994
rect 3627 11942 3639 11994
rect 3691 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 13308 11994
rect 13360 11942 13372 11994
rect 13424 11942 13436 11994
rect 13488 11942 13500 11994
rect 13552 11942 15824 11994
rect 1104 11920 15824 11942
rect 8018 11840 8024 11892
rect 8076 11880 8082 11892
rect 9214 11880 9220 11892
rect 8076 11852 8892 11880
rect 9175 11852 9220 11880
rect 8076 11840 8082 11852
rect 7282 11772 7288 11824
rect 7340 11812 7346 11824
rect 8864 11812 8892 11852
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 10226 11812 10232 11824
rect 7340 11784 7420 11812
rect 8864 11784 10232 11812
rect 7340 11772 7346 11784
rect 7392 11753 7420 11784
rect 10226 11772 10232 11784
rect 10284 11772 10290 11824
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 6638 11636 6644 11688
rect 6696 11676 6702 11688
rect 7193 11679 7251 11685
rect 7193 11676 7205 11679
rect 6696 11648 7205 11676
rect 6696 11636 6702 11648
rect 7193 11645 7205 11648
rect 7239 11645 7251 11679
rect 7193 11639 7251 11645
rect 7282 11636 7288 11688
rect 7340 11676 7346 11688
rect 7837 11679 7895 11685
rect 7837 11676 7849 11679
rect 7340 11648 7849 11676
rect 7340 11636 7346 11648
rect 7837 11645 7849 11648
rect 7883 11645 7895 11679
rect 7837 11639 7895 11645
rect 6546 11568 6552 11620
rect 6604 11608 6610 11620
rect 6604 11580 7788 11608
rect 6604 11568 6610 11580
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 7300 11549 7328 11580
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6788 11512 6837 11540
rect 6788 11500 6794 11512
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 7285 11543 7343 11549
rect 7285 11509 7297 11543
rect 7331 11509 7343 11543
rect 7285 11503 7343 11509
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 7650 11540 7656 11552
rect 7524 11512 7656 11540
rect 7524 11500 7530 11512
rect 7650 11500 7656 11512
rect 7708 11500 7714 11552
rect 7760 11540 7788 11580
rect 8018 11568 8024 11620
rect 8076 11617 8082 11620
rect 8076 11611 8140 11617
rect 8076 11577 8094 11611
rect 8128 11577 8140 11611
rect 8076 11571 8140 11577
rect 8076 11568 8082 11571
rect 8938 11540 8944 11552
rect 7760 11512 8944 11540
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 1104 11450 15824 11472
rect 1104 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 6104 11450
rect 6156 11398 10843 11450
rect 10895 11398 10907 11450
rect 10959 11398 10971 11450
rect 11023 11398 11035 11450
rect 11087 11398 15824 11450
rect 1104 11376 15824 11398
rect 6730 11336 6736 11348
rect 6691 11308 6736 11336
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 12986 11336 12992 11348
rect 9876 11308 12992 11336
rect 6270 11228 6276 11280
rect 6328 11268 6334 11280
rect 6641 11271 6699 11277
rect 6641 11268 6653 11271
rect 6328 11240 6653 11268
rect 6328 11228 6334 11240
rect 6641 11237 6653 11240
rect 6687 11237 6699 11271
rect 6641 11231 6699 11237
rect 7374 11228 7380 11280
rect 7432 11268 7438 11280
rect 7530 11271 7588 11277
rect 7530 11268 7542 11271
rect 7432 11240 7542 11268
rect 7432 11228 7438 11240
rect 7530 11237 7542 11240
rect 7576 11237 7588 11271
rect 7530 11231 7588 11237
rect 7282 11200 7288 11212
rect 7243 11172 7288 11200
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 6963 11104 7328 11132
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 6273 11067 6331 11073
rect 6273 11033 6285 11067
rect 6319 11064 6331 11067
rect 7098 11064 7104 11076
rect 6319 11036 7104 11064
rect 6319 11033 6331 11036
rect 6273 11027 6331 11033
rect 7098 11024 7104 11036
rect 7156 11024 7162 11076
rect 7300 10996 7328 11104
rect 9030 11092 9036 11144
rect 9088 11132 9094 11144
rect 9876 11132 9904 11308
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 10042 11200 10048 11212
rect 9955 11172 10048 11200
rect 10042 11160 10048 11172
rect 10100 11200 10106 11212
rect 10318 11200 10324 11212
rect 10100 11172 10324 11200
rect 10100 11160 10106 11172
rect 10318 11160 10324 11172
rect 10376 11160 10382 11212
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 9088 11104 10149 11132
rect 9088 11092 9094 11104
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 10244 11064 10272 11095
rect 10870 11064 10876 11076
rect 8680 11036 10876 11064
rect 8680 11008 8708 11036
rect 10870 11024 10876 11036
rect 10928 11024 10934 11076
rect 8662 10996 8668 11008
rect 7300 10968 8668 10996
rect 8662 10956 8668 10968
rect 8720 10956 8726 11008
rect 9674 10996 9680 11008
rect 9635 10968 9680 10996
rect 9674 10956 9680 10968
rect 9732 10956 9738 11008
rect 1104 10906 15824 10928
rect 1104 10854 3447 10906
rect 3499 10854 3511 10906
rect 3563 10854 3575 10906
rect 3627 10854 3639 10906
rect 3691 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 13308 10906
rect 13360 10854 13372 10906
rect 13424 10854 13436 10906
rect 13488 10854 13500 10906
rect 13552 10854 15824 10906
rect 1104 10832 15824 10854
rect 13630 10792 13636 10804
rect 5092 10764 13636 10792
rect 4062 10656 4068 10668
rect 4023 10628 4068 10656
rect 4062 10616 4068 10628
rect 4120 10616 4126 10668
rect 5092 10665 5120 10764
rect 13630 10752 13636 10764
rect 13688 10792 13694 10804
rect 13814 10792 13820 10804
rect 13688 10764 13820 10792
rect 13688 10752 13694 10764
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 7282 10684 7288 10736
rect 7340 10724 7346 10736
rect 7377 10727 7435 10733
rect 7377 10724 7389 10727
rect 7340 10696 7389 10724
rect 7340 10684 7346 10696
rect 7377 10693 7389 10696
rect 7423 10724 7435 10727
rect 9033 10727 9091 10733
rect 7423 10696 7696 10724
rect 7423 10693 7435 10696
rect 7377 10687 7435 10693
rect 7668 10665 7696 10696
rect 9033 10693 9045 10727
rect 9079 10724 9091 10727
rect 9079 10696 9904 10724
rect 9079 10693 9091 10696
rect 9033 10687 9091 10693
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10625 5135 10659
rect 5077 10619 5135 10625
rect 7653 10659 7711 10665
rect 7653 10625 7665 10659
rect 7699 10625 7711 10659
rect 7653 10619 7711 10625
rect 1578 10548 1584 10600
rect 1636 10588 1642 10600
rect 3212 10591 3270 10597
rect 3212 10588 3224 10591
rect 1636 10560 3224 10588
rect 1636 10548 1642 10560
rect 3212 10557 3224 10560
rect 3258 10588 3270 10591
rect 3326 10588 3332 10600
rect 3258 10560 3332 10588
rect 3258 10557 3270 10560
rect 3212 10551 3270 10557
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 7190 10548 7196 10600
rect 7248 10588 7254 10600
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 7248 10560 7573 10588
rect 7248 10548 7254 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 9048 10588 9076 10687
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 9876 10665 9904 10696
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9732 10628 9781 10656
rect 9732 10616 9738 10628
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 9769 10619 9827 10625
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10625 9919 10659
rect 10870 10656 10876 10668
rect 10831 10628 10876 10656
rect 9861 10619 9919 10625
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 7800 10560 9076 10588
rect 7800 10548 7806 10560
rect 10594 10548 10600 10600
rect 10652 10588 10658 10600
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10652 10560 10793 10588
rect 10652 10548 10658 10560
rect 10781 10557 10793 10560
rect 10827 10588 10839 10591
rect 15470 10588 15476 10600
rect 10827 10560 15476 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 15470 10548 15476 10560
rect 15528 10548 15534 10600
rect 4157 10523 4215 10529
rect 4157 10489 4169 10523
rect 4203 10489 4215 10523
rect 4157 10483 4215 10489
rect 7920 10523 7978 10529
rect 7920 10489 7932 10523
rect 7966 10520 7978 10523
rect 8662 10520 8668 10532
rect 7966 10492 8668 10520
rect 7966 10489 7978 10492
rect 7920 10483 7978 10489
rect 3283 10455 3341 10461
rect 3283 10421 3295 10455
rect 3329 10452 3341 10455
rect 4172 10452 4200 10483
rect 8662 10480 8668 10492
rect 8720 10480 8726 10532
rect 9677 10523 9735 10529
rect 9677 10489 9689 10523
rect 9723 10520 9735 10523
rect 9723 10492 10364 10520
rect 9723 10489 9735 10492
rect 9677 10483 9735 10489
rect 3329 10424 4200 10452
rect 3329 10421 3341 10424
rect 3283 10415 3341 10421
rect 6730 10412 6736 10464
rect 6788 10452 6794 10464
rect 9122 10452 9128 10464
rect 6788 10424 9128 10452
rect 6788 10412 6794 10424
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9306 10452 9312 10464
rect 9267 10424 9312 10452
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 10336 10461 10364 10492
rect 10321 10455 10379 10461
rect 10321 10421 10333 10455
rect 10367 10421 10379 10455
rect 10686 10452 10692 10464
rect 10647 10424 10692 10452
rect 10321 10415 10379 10421
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 1104 10362 15824 10384
rect 1104 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 6104 10362
rect 6156 10310 10843 10362
rect 10895 10310 10907 10362
rect 10959 10310 10971 10362
rect 11023 10310 11035 10362
rect 11087 10310 15824 10362
rect 1104 10288 15824 10310
rect 6641 10251 6699 10257
rect 6641 10217 6653 10251
rect 6687 10248 6699 10251
rect 9306 10248 9312 10260
rect 6687 10220 9312 10248
rect 6687 10217 6699 10220
rect 6641 10211 6699 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 9677 10251 9735 10257
rect 9677 10217 9689 10251
rect 9723 10248 9735 10251
rect 10686 10248 10692 10260
rect 9723 10220 10692 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 1578 10180 1584 10192
rect 1539 10152 1584 10180
rect 1578 10140 1584 10152
rect 1636 10140 1642 10192
rect 2501 10183 2559 10189
rect 2501 10149 2513 10183
rect 2547 10180 2559 10183
rect 2774 10180 2780 10192
rect 2547 10152 2780 10180
rect 2547 10149 2559 10152
rect 2501 10143 2559 10149
rect 2774 10140 2780 10152
rect 2832 10140 2838 10192
rect 7552 10183 7610 10189
rect 7552 10149 7564 10183
rect 7598 10180 7610 10183
rect 7742 10180 7748 10192
rect 7598 10152 7748 10180
rect 7598 10149 7610 10152
rect 7552 10143 7610 10149
rect 7742 10140 7748 10152
rect 7800 10140 7806 10192
rect 6733 10115 6791 10121
rect 6733 10081 6745 10115
rect 6779 10112 6791 10115
rect 7190 10112 7196 10124
rect 6779 10084 7196 10112
rect 6779 10081 6791 10084
rect 6733 10075 6791 10081
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 7340 10084 7385 10112
rect 7340 10072 7346 10084
rect 1489 10047 1547 10053
rect 1489 10013 1501 10047
rect 1535 10013 1547 10047
rect 1489 10007 1547 10013
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10013 6975 10047
rect 6917 10007 6975 10013
rect 1504 9976 1532 10007
rect 2958 9976 2964 9988
rect 1504 9948 2964 9976
rect 2958 9936 2964 9948
rect 3016 9936 3022 9988
rect 6270 9908 6276 9920
rect 6231 9880 6276 9908
rect 6270 9868 6276 9880
rect 6328 9868 6334 9920
rect 6932 9908 6960 10007
rect 8018 9908 8024 9920
rect 6932 9880 8024 9908
rect 8018 9868 8024 9880
rect 8076 9908 8082 9920
rect 8665 9911 8723 9917
rect 8665 9908 8677 9911
rect 8076 9880 8677 9908
rect 8076 9868 8082 9880
rect 8665 9877 8677 9880
rect 8711 9877 8723 9911
rect 8665 9871 8723 9877
rect 1104 9818 15824 9840
rect 1104 9766 3447 9818
rect 3499 9766 3511 9818
rect 3563 9766 3575 9818
rect 3627 9766 3639 9818
rect 3691 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 13308 9818
rect 13360 9766 13372 9818
rect 13424 9766 13436 9818
rect 13488 9766 13500 9818
rect 13552 9766 15824 9818
rect 1104 9744 15824 9766
rect 6914 9596 6920 9648
rect 6972 9596 6978 9648
rect 7006 9596 7012 9648
rect 7064 9596 7070 9648
rect 7098 9596 7104 9648
rect 7156 9636 7162 9648
rect 7156 9608 7788 9636
rect 7156 9596 7162 9608
rect 6932 9512 6960 9596
rect 6914 9460 6920 9512
rect 6972 9460 6978 9512
rect 4338 9392 4344 9444
rect 4396 9432 4402 9444
rect 7024 9432 7052 9596
rect 7760 9577 7788 9608
rect 8662 9596 8668 9648
rect 8720 9636 8726 9648
rect 8720 9608 8892 9636
rect 8720 9596 8726 9608
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9537 7803 9571
rect 7745 9531 7803 9537
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 8754 9568 8760 9580
rect 7892 9540 7937 9568
rect 8715 9540 8760 9568
rect 7892 9528 7898 9540
rect 8754 9528 8760 9540
rect 8812 9528 8818 9580
rect 8864 9577 8892 9608
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 4396 9404 7052 9432
rect 7653 9435 7711 9441
rect 4396 9392 4402 9404
rect 7653 9401 7665 9435
rect 7699 9432 7711 9435
rect 7699 9404 8340 9432
rect 7699 9401 7711 9404
rect 7653 9395 7711 9401
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 8312 9373 8340 9404
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 7248 9336 7297 9364
rect 7248 9324 7254 9336
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 7285 9327 7343 9333
rect 8297 9367 8355 9373
rect 8297 9333 8309 9367
rect 8343 9333 8355 9367
rect 8297 9327 8355 9333
rect 8665 9367 8723 9373
rect 8665 9333 8677 9367
rect 8711 9364 8723 9367
rect 8846 9364 8852 9376
rect 8711 9336 8852 9364
rect 8711 9333 8723 9336
rect 8665 9327 8723 9333
rect 8846 9324 8852 9336
rect 8904 9364 8910 9376
rect 9490 9364 9496 9376
rect 8904 9336 9496 9364
rect 8904 9324 8910 9336
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 1104 9274 15824 9296
rect 1104 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 6104 9274
rect 6156 9222 10843 9274
rect 10895 9222 10907 9274
rect 10959 9222 10971 9274
rect 11023 9222 11035 9274
rect 11087 9222 15824 9274
rect 1104 9200 15824 9222
rect 12526 9024 12532 9036
rect 12487 8996 12532 9024
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 12713 8959 12771 8965
rect 12713 8956 12725 8959
rect 11204 8928 12725 8956
rect 11204 8916 11210 8928
rect 12713 8925 12725 8928
rect 12759 8925 12771 8959
rect 12713 8919 12771 8925
rect 1104 8730 15824 8752
rect 1104 8678 3447 8730
rect 3499 8678 3511 8730
rect 3563 8678 3575 8730
rect 3627 8678 3639 8730
rect 3691 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 13308 8730
rect 13360 8678 13372 8730
rect 13424 8678 13436 8730
rect 13488 8678 13500 8730
rect 13552 8678 15824 8730
rect 1104 8656 15824 8678
rect 1104 8186 15824 8208
rect 1104 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 6104 8186
rect 6156 8134 10843 8186
rect 10895 8134 10907 8186
rect 10959 8134 10971 8186
rect 11023 8134 11035 8186
rect 11087 8134 15824 8186
rect 1104 8112 15824 8134
rect 6454 8032 6460 8084
rect 6512 8072 6518 8084
rect 7193 8075 7251 8081
rect 7193 8072 7205 8075
rect 6512 8044 7205 8072
rect 6512 8032 6518 8044
rect 7193 8041 7205 8044
rect 7239 8041 7251 8075
rect 7193 8035 7251 8041
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7936 7067 7939
rect 9306 7936 9312 7948
rect 7055 7908 9312 7936
rect 7055 7905 7067 7908
rect 7009 7899 7067 7905
rect 9306 7896 9312 7908
rect 9364 7896 9370 7948
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 11790 7868 11796 7880
rect 7524 7840 11796 7868
rect 7524 7828 7530 7840
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 2682 7760 2688 7812
rect 2740 7800 2746 7812
rect 6362 7800 6368 7812
rect 2740 7772 6368 7800
rect 2740 7760 2746 7772
rect 6362 7760 6368 7772
rect 6420 7760 6426 7812
rect 7650 7760 7656 7812
rect 7708 7800 7714 7812
rect 10962 7800 10968 7812
rect 7708 7772 10968 7800
rect 7708 7760 7714 7772
rect 10962 7760 10968 7772
rect 11020 7760 11026 7812
rect 5166 7692 5172 7744
rect 5224 7732 5230 7744
rect 9122 7732 9128 7744
rect 5224 7704 9128 7732
rect 5224 7692 5230 7704
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 12618 7732 12624 7744
rect 9640 7704 12624 7732
rect 9640 7692 9646 7704
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 1104 7642 15824 7664
rect 1104 7590 3447 7642
rect 3499 7590 3511 7642
rect 3563 7590 3575 7642
rect 3627 7590 3639 7642
rect 3691 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 13308 7642
rect 13360 7590 13372 7642
rect 13424 7590 13436 7642
rect 13488 7590 13500 7642
rect 13552 7590 15824 7642
rect 1104 7568 15824 7590
rect 5074 7528 5080 7540
rect 5035 7500 5080 7528
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 6362 7528 6368 7540
rect 6323 7500 6368 7528
rect 6362 7488 6368 7500
rect 6420 7488 6426 7540
rect 6454 7488 6460 7540
rect 6512 7528 6518 7540
rect 7377 7531 7435 7537
rect 7377 7528 7389 7531
rect 6512 7500 7389 7528
rect 6512 7488 6518 7500
rect 7377 7497 7389 7500
rect 7423 7497 7435 7531
rect 7377 7491 7435 7497
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 9677 7531 9735 7537
rect 9677 7528 9689 7531
rect 8260 7500 9689 7528
rect 8260 7488 8266 7500
rect 9677 7497 9689 7500
rect 9723 7497 9735 7531
rect 10413 7531 10471 7537
rect 10413 7528 10425 7531
rect 9677 7491 9735 7497
rect 9784 7500 10425 7528
rect 5626 7420 5632 7472
rect 5684 7460 5690 7472
rect 7929 7463 7987 7469
rect 7929 7460 7941 7463
rect 5684 7432 7941 7460
rect 5684 7420 5690 7432
rect 7929 7429 7941 7432
rect 7975 7429 7987 7463
rect 7929 7423 7987 7429
rect 8110 7420 8116 7472
rect 8168 7460 8174 7472
rect 9784 7460 9812 7500
rect 10413 7497 10425 7500
rect 10459 7497 10471 7531
rect 10962 7528 10968 7540
rect 10923 7500 10968 7528
rect 10413 7491 10471 7497
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11790 7528 11796 7540
rect 11751 7500 11796 7528
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 12618 7528 12624 7540
rect 12579 7500 12624 7528
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 13998 7460 14004 7472
rect 8168 7432 9812 7460
rect 10244 7432 14004 7460
rect 8168 7420 8174 7432
rect 6270 7392 6276 7404
rect 3252 7364 6276 7392
rect 3252 7333 3280 7364
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 10042 7392 10048 7404
rect 8312 7364 10048 7392
rect 3237 7327 3295 7333
rect 3237 7293 3249 7327
rect 3283 7293 3295 7327
rect 3237 7287 3295 7293
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7324 4951 7327
rect 5534 7324 5540 7336
rect 4939 7296 5540 7324
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 6181 7327 6239 7333
rect 6181 7293 6193 7327
rect 6227 7324 6239 7327
rect 7098 7324 7104 7336
rect 6227 7296 7104 7324
rect 6227 7293 6239 7296
rect 6181 7287 6239 7293
rect 3050 7216 3056 7268
rect 3108 7256 3114 7268
rect 3513 7259 3571 7265
rect 3513 7256 3525 7259
rect 3108 7228 3525 7256
rect 3108 7216 3114 7228
rect 3513 7225 3525 7228
rect 3559 7225 3571 7259
rect 5644 7256 5672 7287
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 8312 7333 8340 7364
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 7193 7327 7251 7333
rect 7193 7293 7205 7327
rect 7239 7324 7251 7327
rect 7561 7327 7619 7333
rect 7561 7324 7573 7327
rect 7239 7296 7573 7324
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 7561 7293 7573 7296
rect 7607 7293 7619 7327
rect 7561 7287 7619 7293
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 8297 7327 8355 7333
rect 8297 7293 8309 7327
rect 8343 7293 8355 7327
rect 8297 7287 8355 7293
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7293 8999 7327
rect 9490 7324 9496 7336
rect 9451 7296 9496 7324
rect 8941 7287 8999 7293
rect 7650 7256 7656 7268
rect 5644 7228 7656 7256
rect 3513 7219 3571 7225
rect 7650 7216 7656 7228
rect 7708 7216 7714 7268
rect 7760 7256 7788 7287
rect 8846 7256 8852 7268
rect 7760 7228 8852 7256
rect 8846 7216 8852 7228
rect 8904 7216 8910 7268
rect 8956 7256 8984 7287
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 10244 7333 10272 7432
rect 13998 7420 14004 7432
rect 14056 7420 14062 7472
rect 15010 7392 15016 7404
rect 10796 7364 15016 7392
rect 10796 7333 10824 7364
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 10229 7327 10287 7333
rect 10229 7293 10241 7327
rect 10275 7293 10287 7327
rect 10229 7287 10287 7293
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 11609 7327 11667 7333
rect 11609 7293 11621 7327
rect 11655 7293 11667 7327
rect 11609 7287 11667 7293
rect 12437 7327 12495 7333
rect 12437 7293 12449 7327
rect 12483 7324 12495 7327
rect 16850 7324 16856 7336
rect 12483 7296 16856 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 10686 7256 10692 7268
rect 8956 7228 10692 7256
rect 10686 7216 10692 7228
rect 10744 7216 10750 7268
rect 11624 7256 11652 7287
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 13722 7256 13728 7268
rect 11624 7228 13728 7256
rect 13722 7216 13728 7228
rect 13780 7216 13786 7268
rect 1854 7148 1860 7200
rect 1912 7188 1918 7200
rect 5813 7191 5871 7197
rect 5813 7188 5825 7191
rect 1912 7160 5825 7188
rect 1912 7148 1918 7160
rect 5813 7157 5825 7160
rect 5859 7157 5871 7191
rect 5813 7151 5871 7157
rect 7561 7191 7619 7197
rect 7561 7157 7573 7191
rect 7607 7188 7619 7191
rect 8294 7188 8300 7200
rect 7607 7160 8300 7188
rect 7607 7157 7619 7160
rect 7561 7151 7619 7157
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 8478 7188 8484 7200
rect 8439 7160 8484 7188
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 9122 7188 9128 7200
rect 9083 7160 9128 7188
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 1104 7098 15824 7120
rect 1104 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 6104 7098
rect 6156 7046 10843 7098
rect 10895 7046 10907 7098
rect 10959 7046 10971 7098
rect 11023 7046 11035 7098
rect 11087 7046 15824 7098
rect 1104 7024 15824 7046
rect 4430 6944 4436 6996
rect 4488 6984 4494 6996
rect 8478 6984 8484 6996
rect 4488 6956 8484 6984
rect 4488 6944 4494 6956
rect 8478 6944 8484 6956
rect 8536 6944 8542 6996
rect 9490 6944 9496 6996
rect 9548 6984 9554 6996
rect 13814 6984 13820 6996
rect 9548 6956 13820 6984
rect 9548 6944 9554 6956
rect 13814 6944 13820 6956
rect 13872 6944 13878 6996
rect 8202 6916 8208 6928
rect 6288 6888 8208 6916
rect 4798 6848 4804 6860
rect 4759 6820 4804 6848
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 5626 6848 5632 6860
rect 5587 6820 5632 6848
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 6288 6857 6316 6888
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 15102 6916 15108 6928
rect 8404 6888 9536 6916
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6817 6331 6851
rect 6273 6811 6331 6817
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 6825 6851 6883 6857
rect 6825 6848 6837 6851
rect 6788 6820 6837 6848
rect 6788 6808 6794 6820
rect 6825 6817 6837 6820
rect 6871 6817 6883 6851
rect 6825 6811 6883 6817
rect 7377 6851 7435 6857
rect 7377 6817 7389 6851
rect 7423 6817 7435 6851
rect 7926 6848 7932 6860
rect 7887 6820 7932 6848
rect 7377 6811 7435 6817
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 7392 6780 7420 6811
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 8404 6780 8432 6888
rect 8481 6851 8539 6857
rect 8481 6817 8493 6851
rect 8527 6817 8539 6851
rect 8481 6811 8539 6817
rect 9033 6851 9091 6857
rect 9033 6817 9045 6851
rect 9079 6848 9091 6851
rect 9398 6848 9404 6860
rect 9079 6820 9404 6848
rect 9079 6817 9091 6820
rect 9033 6811 9091 6817
rect 4948 6752 7052 6780
rect 7392 6752 8432 6780
rect 8496 6780 8524 6811
rect 9398 6808 9404 6820
rect 9456 6808 9462 6860
rect 9214 6780 9220 6792
rect 8496 6752 9220 6780
rect 4948 6740 4954 6752
rect 4614 6672 4620 6724
rect 4672 6712 4678 6724
rect 7024 6721 7052 6752
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9508 6780 9536 6888
rect 10704 6888 15108 6916
rect 9950 6848 9956 6860
rect 9911 6820 9956 6848
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 10704 6857 10732 6888
rect 15102 6876 15108 6888
rect 15160 6876 15166 6928
rect 10689 6851 10747 6857
rect 10689 6817 10701 6851
rect 10735 6817 10747 6851
rect 10689 6811 10747 6817
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6817 11483 6851
rect 11974 6848 11980 6860
rect 11935 6820 11980 6848
rect 11425 6811 11483 6817
rect 10410 6780 10416 6792
rect 9508 6752 10416 6780
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 11440 6780 11468 6811
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 12529 6851 12587 6857
rect 12529 6817 12541 6851
rect 12575 6848 12587 6851
rect 16758 6848 16764 6860
rect 12575 6820 16764 6848
rect 12575 6817 12587 6820
rect 12529 6811 12587 6817
rect 16758 6808 16764 6820
rect 16816 6808 16822 6860
rect 14550 6780 14556 6792
rect 11440 6752 14556 6780
rect 14550 6740 14556 6752
rect 14608 6740 14614 6792
rect 6457 6715 6515 6721
rect 6457 6712 6469 6715
rect 4672 6684 6469 6712
rect 4672 6672 4678 6684
rect 6457 6681 6469 6684
rect 6503 6681 6515 6715
rect 6457 6675 6515 6681
rect 7009 6715 7067 6721
rect 7009 6681 7021 6715
rect 7055 6681 7067 6715
rect 10134 6712 10140 6724
rect 7009 6675 7067 6681
rect 7116 6684 9260 6712
rect 10095 6684 10140 6712
rect 4982 6644 4988 6656
rect 4943 6616 4988 6644
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 5074 6604 5080 6656
rect 5132 6644 5138 6656
rect 5813 6647 5871 6653
rect 5813 6644 5825 6647
rect 5132 6616 5825 6644
rect 5132 6604 5138 6616
rect 5813 6613 5825 6616
rect 5859 6613 5871 6647
rect 5813 6607 5871 6613
rect 5902 6604 5908 6656
rect 5960 6644 5966 6656
rect 7116 6644 7144 6684
rect 7558 6644 7564 6656
rect 5960 6616 7144 6644
rect 7519 6616 7564 6644
rect 5960 6604 5966 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 8110 6644 8116 6656
rect 8071 6616 8116 6644
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 8662 6644 8668 6656
rect 8623 6616 8668 6644
rect 8662 6604 8668 6616
rect 8720 6604 8726 6656
rect 9232 6653 9260 6684
rect 10134 6672 10140 6684
rect 10192 6672 10198 6724
rect 12158 6712 12164 6724
rect 12119 6684 12164 6712
rect 12158 6672 12164 6684
rect 12216 6672 12222 6724
rect 9217 6647 9275 6653
rect 9217 6613 9229 6647
rect 9263 6613 9275 6647
rect 9217 6607 9275 6613
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 10873 6647 10931 6653
rect 10873 6644 10885 6647
rect 9732 6616 10885 6644
rect 9732 6604 9738 6616
rect 10873 6613 10885 6616
rect 10919 6613 10931 6647
rect 11606 6644 11612 6656
rect 11567 6616 11612 6644
rect 10873 6607 10931 6613
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 12710 6644 12716 6656
rect 12671 6616 12716 6644
rect 12710 6604 12716 6616
rect 12768 6604 12774 6656
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 4798 6400 4804 6452
rect 4856 6440 4862 6452
rect 8662 6440 8668 6452
rect 4856 6412 8668 6440
rect 4856 6400 4862 6412
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 9858 6440 9864 6452
rect 8772 6412 9864 6440
rect 7929 6375 7987 6381
rect 7929 6341 7941 6375
rect 7975 6341 7987 6375
rect 7929 6335 7987 6341
rect 7834 6304 7840 6316
rect 7576 6276 7840 6304
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6205 3755 6239
rect 4338 6236 4344 6248
rect 4299 6208 4344 6236
rect 3697 6199 3755 6205
rect 3712 6168 3740 6199
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 5169 6239 5227 6245
rect 5169 6205 5181 6239
rect 5215 6236 5227 6239
rect 7576 6236 7604 6276
rect 7834 6264 7840 6276
rect 7892 6264 7898 6316
rect 7944 6248 7972 6335
rect 8018 6332 8024 6384
rect 8076 6372 8082 6384
rect 8772 6372 8800 6412
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 14274 6440 14280 6452
rect 12032 6412 14280 6440
rect 12032 6400 12038 6412
rect 14274 6400 14280 6412
rect 14332 6400 14338 6452
rect 8076 6344 8800 6372
rect 8076 6332 8082 6344
rect 9490 6332 9496 6384
rect 9548 6372 9554 6384
rect 9585 6375 9643 6381
rect 9585 6372 9597 6375
rect 9548 6344 9597 6372
rect 9548 6332 9554 6344
rect 9585 6341 9597 6344
rect 9631 6341 9643 6375
rect 9585 6335 9643 6341
rect 9950 6332 9956 6384
rect 10008 6372 10014 6384
rect 14182 6372 14188 6384
rect 10008 6344 14188 6372
rect 10008 6332 10014 6344
rect 14182 6332 14188 6344
rect 14240 6332 14246 6384
rect 14642 6304 14648 6316
rect 10244 6276 14648 6304
rect 7742 6236 7748 6248
rect 5215 6208 7604 6236
rect 7703 6208 7748 6236
rect 5215 6205 5227 6208
rect 5169 6199 5227 6205
rect 7742 6196 7748 6208
rect 7800 6196 7806 6248
rect 7926 6196 7932 6248
rect 7984 6196 7990 6248
rect 9398 6236 9404 6248
rect 9359 6208 9404 6236
rect 9398 6196 9404 6208
rect 9456 6196 9462 6248
rect 10244 6245 10272 6276
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 10229 6239 10287 6245
rect 10229 6205 10241 6239
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 11517 6239 11575 6245
rect 11517 6205 11529 6239
rect 11563 6236 11575 6239
rect 14366 6236 14372 6248
rect 11563 6208 14372 6236
rect 11563 6205 11575 6208
rect 11517 6199 11575 6205
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 6546 6168 6552 6180
rect 3712 6140 6552 6168
rect 6546 6128 6552 6140
rect 6604 6128 6610 6180
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 7432 6140 11744 6168
rect 7432 6128 7438 6140
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 3881 6103 3939 6109
rect 3881 6100 3893 6103
rect 1452 6072 3893 6100
rect 1452 6060 1458 6072
rect 3881 6069 3893 6072
rect 3927 6069 3939 6103
rect 4522 6100 4528 6112
rect 4483 6072 4528 6100
rect 3881 6063 3939 6069
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 5350 6100 5356 6112
rect 5311 6072 5356 6100
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 9766 6100 9772 6112
rect 8260 6072 9772 6100
rect 8260 6060 8266 6072
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10410 6100 10416 6112
rect 10371 6072 10416 6100
rect 10410 6060 10416 6072
rect 10468 6060 10474 6112
rect 11716 6109 11744 6140
rect 11701 6103 11759 6109
rect 11701 6069 11713 6103
rect 11747 6069 11759 6103
rect 11701 6063 11759 6069
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 11882 5896 11888 5908
rect 8680 5868 11888 5896
rect 7742 5788 7748 5840
rect 7800 5828 7806 5840
rect 8680 5828 8708 5868
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 7800 5800 8708 5828
rect 7800 5788 7806 5800
rect 9398 5788 9404 5840
rect 9456 5828 9462 5840
rect 14090 5828 14096 5840
rect 9456 5800 14096 5828
rect 9456 5788 9462 5800
rect 14090 5788 14096 5800
rect 14148 5788 14154 5840
rect 7561 5763 7619 5769
rect 7561 5729 7573 5763
rect 7607 5760 7619 5763
rect 9030 5760 9036 5772
rect 7607 5732 9036 5760
rect 7607 5729 7619 5732
rect 7561 5723 7619 5729
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 10594 5760 10600 5772
rect 9723 5732 10600 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 10502 5692 10508 5704
rect 5684 5664 10508 5692
rect 5684 5652 5690 5664
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 7006 5584 7012 5636
rect 7064 5624 7070 5636
rect 9861 5627 9919 5633
rect 9861 5624 9873 5627
rect 7064 5596 9873 5624
rect 7064 5584 7070 5596
rect 9861 5593 9873 5596
rect 9907 5593 9919 5627
rect 9861 5587 9919 5593
rect 4430 5516 4436 5568
rect 4488 5556 4494 5568
rect 7745 5559 7803 5565
rect 7745 5556 7757 5559
rect 4488 5528 7757 5556
rect 4488 5516 4494 5528
rect 7745 5525 7757 5528
rect 7791 5525 7803 5559
rect 7745 5519 7803 5525
rect 7834 5516 7840 5568
rect 7892 5556 7898 5568
rect 11606 5556 11612 5568
rect 7892 5528 11612 5556
rect 7892 5516 7898 5528
rect 11606 5516 11612 5528
rect 11664 5516 11670 5568
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 10318 4700 10324 4752
rect 10376 4740 10382 4752
rect 15470 4740 15476 4752
rect 10376 4712 15476 4740
rect 10376 4700 10382 4712
rect 15470 4700 15476 4712
rect 15528 4700 15534 4752
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 9582 4156 9588 4208
rect 9640 4196 9646 4208
rect 9640 4168 10548 4196
rect 9640 4156 9646 4168
rect 5258 4088 5264 4140
rect 5316 4128 5322 4140
rect 9490 4128 9496 4140
rect 5316 4100 9496 4128
rect 5316 4088 5322 4100
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 10410 4060 10416 4072
rect 6328 4032 10416 4060
rect 6328 4020 6334 4032
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 10520 4060 10548 4168
rect 14274 4088 14280 4140
rect 14332 4128 14338 4140
rect 16298 4128 16304 4140
rect 14332 4100 16304 4128
rect 14332 4088 14338 4100
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 12894 4060 12900 4072
rect 10520 4032 12900 4060
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 13722 4020 13728 4072
rect 13780 4060 13786 4072
rect 15930 4060 15936 4072
rect 13780 4032 15936 4060
rect 13780 4020 13786 4032
rect 15930 4020 15936 4032
rect 15988 4020 15994 4072
rect 3142 3952 3148 4004
rect 3200 3992 3206 4004
rect 7558 3992 7564 4004
rect 3200 3964 7564 3992
rect 3200 3952 3206 3964
rect 7558 3952 7564 3964
rect 7616 3952 7622 4004
rect 7650 3952 7656 4004
rect 7708 3992 7714 4004
rect 9950 3992 9956 4004
rect 7708 3964 9956 3992
rect 7708 3952 7714 3964
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 8110 3924 8116 3936
rect 4028 3896 8116 3924
rect 4028 3884 4034 3896
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 9306 3884 9312 3936
rect 9364 3924 9370 3936
rect 11238 3924 11244 3936
rect 9364 3896 11244 3924
rect 9364 3884 9370 3896
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 9122 3720 9128 3732
rect 5592 3692 9128 3720
rect 5592 3680 5598 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 6914 3612 6920 3664
rect 6972 3652 6978 3664
rect 9490 3652 9496 3664
rect 6972 3624 9496 3652
rect 6972 3612 6978 3624
rect 9490 3612 9496 3624
rect 9548 3612 9554 3664
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 11606 3584 11612 3596
rect 8812 3556 11612 3584
rect 8812 3544 8818 3556
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 13170 3516 13176 3528
rect 10744 3488 13176 3516
rect 10744 3476 10750 3488
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 2314 3408 2320 3460
rect 2372 3448 2378 3460
rect 4614 3448 4620 3460
rect 2372 3420 4620 3448
rect 2372 3408 2378 3420
rect 4614 3408 4620 3420
rect 4672 3408 4678 3460
rect 6546 3408 6552 3460
rect 6604 3448 6610 3460
rect 9674 3448 9680 3460
rect 6604 3420 9680 3448
rect 6604 3408 6610 3420
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 566 3340 572 3392
rect 624 3380 630 3392
rect 4982 3380 4988 3392
rect 624 3352 4988 3380
rect 624 3340 630 3352
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 8202 3340 8208 3392
rect 8260 3380 8266 3392
rect 12710 3380 12716 3392
rect 8260 3352 12716 3380
rect 8260 3340 8266 3352
rect 12710 3340 12716 3352
rect 12768 3340 12774 3392
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 7098 3136 7104 3188
rect 7156 3176 7162 3188
rect 10686 3176 10692 3188
rect 7156 3148 10692 3176
rect 7156 3136 7162 3148
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 198 3068 204 3120
rect 256 3108 262 3120
rect 1394 3108 1400 3120
rect 256 3080 1400 3108
rect 256 3068 262 3080
rect 1394 3068 1400 3080
rect 1452 3068 1458 3120
rect 1854 3068 1860 3120
rect 1912 3108 1918 3120
rect 5350 3108 5356 3120
rect 1912 3080 5356 3108
rect 1912 3068 1918 3080
rect 5350 3068 5356 3080
rect 5408 3068 5414 3120
rect 8846 3068 8852 3120
rect 8904 3108 8910 3120
rect 12066 3108 12072 3120
rect 8904 3080 12072 3108
rect 8904 3068 8910 3080
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 2682 3000 2688 3052
rect 2740 3040 2746 3052
rect 4890 3040 4896 3052
rect 2740 3012 4896 3040
rect 2740 3000 2746 3012
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 10042 3000 10048 3052
rect 10100 3040 10106 3052
rect 12526 3040 12532 3052
rect 10100 3012 12532 3040
rect 10100 3000 10106 3012
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 1118 2932 1124 2984
rect 1176 2972 1182 2984
rect 2958 2972 2964 2984
rect 1176 2944 2964 2972
rect 1176 2932 1182 2944
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 1026 2864 1032 2916
rect 1084 2904 1090 2916
rect 4522 2904 4528 2916
rect 1084 2876 4528 2904
rect 1084 2864 1090 2876
rect 4522 2864 4528 2876
rect 4580 2864 4586 2916
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 5074 2836 5080 2848
rect 1452 2808 5080 2836
rect 1452 2796 1458 2808
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 3602 1436 3608 1488
rect 3660 1476 3666 1488
rect 7926 1476 7932 1488
rect 3660 1448 7932 1476
rect 3660 1436 3666 1448
rect 7926 1436 7932 1448
rect 7984 1436 7990 1488
rect 13998 552 14004 604
rect 14056 592 14062 604
rect 14642 592 14648 604
rect 14056 564 14648 592
rect 14056 552 14062 564
rect 14642 552 14648 564
rect 14700 552 14706 604
<< via1 >>
rect 3447 17382 3499 17434
rect 3511 17382 3563 17434
rect 3575 17382 3627 17434
rect 3639 17382 3691 17434
rect 8378 17382 8430 17434
rect 8442 17382 8494 17434
rect 8506 17382 8558 17434
rect 8570 17382 8622 17434
rect 13308 17382 13360 17434
rect 13372 17382 13424 17434
rect 13436 17382 13488 17434
rect 13500 17382 13552 17434
rect 9772 17008 9824 17060
rect 10968 17008 11020 17060
rect 5912 16838 5964 16890
rect 5976 16838 6028 16890
rect 6040 16838 6092 16890
rect 6104 16838 6156 16890
rect 10843 16838 10895 16890
rect 10907 16838 10959 16890
rect 10971 16838 11023 16890
rect 11035 16838 11087 16890
rect 4804 16396 4856 16448
rect 9312 16396 9364 16448
rect 3447 16294 3499 16346
rect 3511 16294 3563 16346
rect 3575 16294 3627 16346
rect 3639 16294 3691 16346
rect 8378 16294 8430 16346
rect 8442 16294 8494 16346
rect 8506 16294 8558 16346
rect 8570 16294 8622 16346
rect 13308 16294 13360 16346
rect 13372 16294 13424 16346
rect 13436 16294 13488 16346
rect 13500 16294 13552 16346
rect 3056 16192 3108 16244
rect 6460 16192 6512 16244
rect 9128 16192 9180 16244
rect 11336 16192 11388 16244
rect 5540 16124 5592 16176
rect 8208 16124 8260 16176
rect 6368 16056 6420 16108
rect 8116 16056 8168 16108
rect 3884 15988 3936 16040
rect 5632 15988 5684 16040
rect 6828 15988 6880 16040
rect 7840 15988 7892 16040
rect 8668 15988 8720 16040
rect 9588 15988 9640 16040
rect 14556 15988 14608 16040
rect 16304 15988 16356 16040
rect 3332 15920 3384 15972
rect 6368 15920 6420 15972
rect 7932 15920 7984 15972
rect 12624 15920 12676 15972
rect 4712 15852 4764 15904
rect 6828 15852 6880 15904
rect 8024 15852 8076 15904
rect 12164 15852 12216 15904
rect 5912 15750 5964 15802
rect 5976 15750 6028 15802
rect 6040 15750 6092 15802
rect 6104 15750 6156 15802
rect 10843 15750 10895 15802
rect 10907 15750 10959 15802
rect 10971 15750 11023 15802
rect 11035 15750 11087 15802
rect 1400 15648 1452 15700
rect 4712 15648 4764 15700
rect 6276 15648 6328 15700
rect 10048 15648 10100 15700
rect 9404 15580 9456 15632
rect 14280 15580 14332 15632
rect 1032 15444 1084 15496
rect 5080 15444 5132 15496
rect 9312 15444 9364 15496
rect 13176 15444 13228 15496
rect 14372 15444 14424 15496
rect 15936 15444 15988 15496
rect 2228 15376 2280 15428
rect 5540 15376 5592 15428
rect 7012 15376 7064 15428
rect 9680 15376 9732 15428
rect 204 15308 256 15360
rect 2872 15308 2924 15360
rect 7196 15308 7248 15360
rect 9496 15308 9548 15360
rect 3447 15206 3499 15258
rect 3511 15206 3563 15258
rect 3575 15206 3627 15258
rect 3639 15206 3691 15258
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 13308 15206 13360 15258
rect 13372 15206 13424 15258
rect 13436 15206 13488 15258
rect 13500 15206 13552 15258
rect 572 15104 624 15156
rect 4712 15147 4764 15156
rect 4712 15113 4721 15147
rect 4721 15113 4755 15147
rect 4755 15113 4764 15147
rect 4712 15104 4764 15113
rect 5540 15147 5592 15156
rect 5540 15113 5549 15147
rect 5549 15113 5583 15147
rect 5583 15113 5592 15147
rect 5540 15104 5592 15113
rect 6828 15104 6880 15156
rect 9496 15147 9548 15156
rect 9496 15113 9505 15147
rect 9505 15113 9539 15147
rect 9539 15113 9548 15147
rect 9496 15104 9548 15113
rect 6736 14968 6788 15020
rect 6552 14832 6604 14884
rect 8944 14900 8996 14952
rect 9864 14900 9916 14952
rect 8024 14832 8076 14884
rect 5912 14662 5964 14714
rect 5976 14662 6028 14714
rect 6040 14662 6092 14714
rect 6104 14662 6156 14714
rect 10843 14662 10895 14714
rect 10907 14662 10959 14714
rect 10971 14662 11023 14714
rect 11035 14662 11087 14714
rect 3447 14118 3499 14170
rect 3511 14118 3563 14170
rect 3575 14118 3627 14170
rect 3639 14118 3691 14170
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 13308 14118 13360 14170
rect 13372 14118 13424 14170
rect 13436 14118 13488 14170
rect 13500 14118 13552 14170
rect 7380 13948 7432 14000
rect 3792 13880 3844 13932
rect 4344 13855 4396 13864
rect 4344 13821 4353 13855
rect 4353 13821 4387 13855
rect 4387 13821 4396 13855
rect 4344 13812 4396 13821
rect 5912 13574 5964 13626
rect 5976 13574 6028 13626
rect 6040 13574 6092 13626
rect 6104 13574 6156 13626
rect 10843 13574 10895 13626
rect 10907 13574 10959 13626
rect 10971 13574 11023 13626
rect 11035 13574 11087 13626
rect 4344 13472 4396 13524
rect 13728 13472 13780 13524
rect 2872 13379 2924 13388
rect 2872 13345 2881 13379
rect 2881 13345 2915 13379
rect 2915 13345 2924 13379
rect 2872 13336 2924 13345
rect 7196 13336 7248 13388
rect 9220 13268 9272 13320
rect 3332 13175 3384 13184
rect 3332 13141 3341 13175
rect 3341 13141 3375 13175
rect 3375 13141 3384 13175
rect 3332 13132 3384 13141
rect 13820 13132 13872 13184
rect 3447 13030 3499 13082
rect 3511 13030 3563 13082
rect 3575 13030 3627 13082
rect 3639 13030 3691 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 13308 13030 13360 13082
rect 13372 13030 13424 13082
rect 13436 13030 13488 13082
rect 13500 13030 13552 13082
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 6736 12724 6788 12776
rect 6920 12724 6972 12776
rect 7012 12656 7064 12708
rect 6276 12588 6328 12640
rect 9220 12588 9272 12640
rect 13728 12588 13780 12640
rect 5912 12486 5964 12538
rect 5976 12486 6028 12538
rect 6040 12486 6092 12538
rect 6104 12486 6156 12538
rect 10843 12486 10895 12538
rect 10907 12486 10959 12538
rect 10971 12486 11023 12538
rect 11035 12486 11087 12538
rect 6644 12384 6696 12436
rect 8852 12384 8904 12436
rect 11152 12316 11204 12368
rect 9864 12248 9916 12300
rect 10508 12248 10560 12300
rect 8024 12180 8076 12232
rect 7288 12112 7340 12164
rect 7196 12044 7248 12096
rect 8760 12044 8812 12096
rect 3447 11942 3499 11994
rect 3511 11942 3563 11994
rect 3575 11942 3627 11994
rect 3639 11942 3691 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 13308 11942 13360 11994
rect 13372 11942 13424 11994
rect 13436 11942 13488 11994
rect 13500 11942 13552 11994
rect 8024 11840 8076 11892
rect 9220 11883 9272 11892
rect 7288 11772 7340 11824
rect 9220 11849 9229 11883
rect 9229 11849 9263 11883
rect 9263 11849 9272 11883
rect 9220 11840 9272 11849
rect 10232 11772 10284 11824
rect 6644 11636 6696 11688
rect 7288 11636 7340 11688
rect 6552 11568 6604 11620
rect 6736 11500 6788 11552
rect 7472 11500 7524 11552
rect 7656 11500 7708 11552
rect 8024 11568 8076 11620
rect 8944 11500 8996 11552
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 6104 11398 6156 11450
rect 10843 11398 10895 11450
rect 10907 11398 10959 11450
rect 10971 11398 11023 11450
rect 11035 11398 11087 11450
rect 6736 11339 6788 11348
rect 6736 11305 6745 11339
rect 6745 11305 6779 11339
rect 6779 11305 6788 11339
rect 6736 11296 6788 11305
rect 6276 11228 6328 11280
rect 7380 11228 7432 11280
rect 7288 11203 7340 11212
rect 7288 11169 7297 11203
rect 7297 11169 7331 11203
rect 7331 11169 7340 11203
rect 7288 11160 7340 11169
rect 7104 11024 7156 11076
rect 9036 11092 9088 11144
rect 12992 11296 13044 11348
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 10324 11160 10376 11212
rect 10876 11024 10928 11076
rect 8668 10999 8720 11008
rect 8668 10965 8677 10999
rect 8677 10965 8711 10999
rect 8711 10965 8720 10999
rect 8668 10956 8720 10965
rect 9680 10999 9732 11008
rect 9680 10965 9689 10999
rect 9689 10965 9723 10999
rect 9723 10965 9732 10999
rect 9680 10956 9732 10965
rect 3447 10854 3499 10906
rect 3511 10854 3563 10906
rect 3575 10854 3627 10906
rect 3639 10854 3691 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 13308 10854 13360 10906
rect 13372 10854 13424 10906
rect 13436 10854 13488 10906
rect 13500 10854 13552 10906
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 13636 10752 13688 10804
rect 13820 10752 13872 10804
rect 7288 10684 7340 10736
rect 1584 10548 1636 10600
rect 3332 10548 3384 10600
rect 7196 10548 7248 10600
rect 7748 10548 7800 10600
rect 9680 10616 9732 10668
rect 10876 10659 10928 10668
rect 10876 10625 10885 10659
rect 10885 10625 10919 10659
rect 10919 10625 10928 10659
rect 10876 10616 10928 10625
rect 10600 10548 10652 10600
rect 15476 10548 15528 10600
rect 8668 10480 8720 10532
rect 6736 10412 6788 10464
rect 9128 10412 9180 10464
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 10692 10455 10744 10464
rect 10692 10421 10701 10455
rect 10701 10421 10735 10455
rect 10735 10421 10744 10455
rect 10692 10412 10744 10421
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 6104 10310 6156 10362
rect 10843 10310 10895 10362
rect 10907 10310 10959 10362
rect 10971 10310 11023 10362
rect 11035 10310 11087 10362
rect 9312 10208 9364 10260
rect 10692 10208 10744 10260
rect 1584 10183 1636 10192
rect 1584 10149 1593 10183
rect 1593 10149 1627 10183
rect 1627 10149 1636 10183
rect 1584 10140 1636 10149
rect 2780 10140 2832 10192
rect 7748 10140 7800 10192
rect 7196 10072 7248 10124
rect 7288 10115 7340 10124
rect 7288 10081 7297 10115
rect 7297 10081 7331 10115
rect 7331 10081 7340 10115
rect 7288 10072 7340 10081
rect 2964 9936 3016 9988
rect 6276 9911 6328 9920
rect 6276 9877 6285 9911
rect 6285 9877 6319 9911
rect 6319 9877 6328 9911
rect 6276 9868 6328 9877
rect 8024 9868 8076 9920
rect 3447 9766 3499 9818
rect 3511 9766 3563 9818
rect 3575 9766 3627 9818
rect 3639 9766 3691 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 13308 9766 13360 9818
rect 13372 9766 13424 9818
rect 13436 9766 13488 9818
rect 13500 9766 13552 9818
rect 6920 9596 6972 9648
rect 7012 9596 7064 9648
rect 7104 9596 7156 9648
rect 6920 9460 6972 9512
rect 4344 9392 4396 9444
rect 8668 9596 8720 9648
rect 7840 9571 7892 9580
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 8760 9571 8812 9580
rect 7840 9528 7892 9537
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 7196 9324 7248 9376
rect 8852 9324 8904 9376
rect 9496 9324 9548 9376
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 6104 9222 6156 9274
rect 10843 9222 10895 9274
rect 10907 9222 10959 9274
rect 10971 9222 11023 9274
rect 11035 9222 11087 9274
rect 12532 9027 12584 9036
rect 12532 8993 12541 9027
rect 12541 8993 12575 9027
rect 12575 8993 12584 9027
rect 12532 8984 12584 8993
rect 11152 8916 11204 8968
rect 3447 8678 3499 8730
rect 3511 8678 3563 8730
rect 3575 8678 3627 8730
rect 3639 8678 3691 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 13308 8678 13360 8730
rect 13372 8678 13424 8730
rect 13436 8678 13488 8730
rect 13500 8678 13552 8730
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 6104 8134 6156 8186
rect 10843 8134 10895 8186
rect 10907 8134 10959 8186
rect 10971 8134 11023 8186
rect 11035 8134 11087 8186
rect 6460 8032 6512 8084
rect 9312 7896 9364 7948
rect 7472 7828 7524 7880
rect 11796 7828 11848 7880
rect 2688 7760 2740 7812
rect 6368 7760 6420 7812
rect 7656 7760 7708 7812
rect 10968 7760 11020 7812
rect 5172 7692 5224 7744
rect 9128 7692 9180 7744
rect 9588 7692 9640 7744
rect 12624 7692 12676 7744
rect 3447 7590 3499 7642
rect 3511 7590 3563 7642
rect 3575 7590 3627 7642
rect 3639 7590 3691 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 13308 7590 13360 7642
rect 13372 7590 13424 7642
rect 13436 7590 13488 7642
rect 13500 7590 13552 7642
rect 5080 7531 5132 7540
rect 5080 7497 5089 7531
rect 5089 7497 5123 7531
rect 5123 7497 5132 7531
rect 5080 7488 5132 7497
rect 6368 7531 6420 7540
rect 6368 7497 6377 7531
rect 6377 7497 6411 7531
rect 6411 7497 6420 7531
rect 6368 7488 6420 7497
rect 6460 7488 6512 7540
rect 8208 7488 8260 7540
rect 5632 7420 5684 7472
rect 8116 7420 8168 7472
rect 10968 7531 11020 7540
rect 10968 7497 10977 7531
rect 10977 7497 11011 7531
rect 11011 7497 11020 7531
rect 10968 7488 11020 7497
rect 11796 7531 11848 7540
rect 11796 7497 11805 7531
rect 11805 7497 11839 7531
rect 11839 7497 11848 7531
rect 11796 7488 11848 7497
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 6276 7352 6328 7404
rect 5540 7284 5592 7336
rect 3056 7216 3108 7268
rect 7104 7284 7156 7336
rect 10048 7352 10100 7404
rect 9496 7327 9548 7336
rect 7656 7216 7708 7268
rect 8852 7216 8904 7268
rect 9496 7293 9505 7327
rect 9505 7293 9539 7327
rect 9539 7293 9548 7327
rect 9496 7284 9548 7293
rect 14004 7420 14056 7472
rect 15016 7352 15068 7404
rect 10692 7216 10744 7268
rect 16856 7284 16908 7336
rect 13728 7216 13780 7268
rect 1860 7148 1912 7200
rect 8300 7148 8352 7200
rect 8484 7191 8536 7200
rect 8484 7157 8493 7191
rect 8493 7157 8527 7191
rect 8527 7157 8536 7191
rect 8484 7148 8536 7157
rect 9128 7191 9180 7200
rect 9128 7157 9137 7191
rect 9137 7157 9171 7191
rect 9171 7157 9180 7191
rect 9128 7148 9180 7157
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 6104 7046 6156 7098
rect 10843 7046 10895 7098
rect 10907 7046 10959 7098
rect 10971 7046 11023 7098
rect 11035 7046 11087 7098
rect 4436 6944 4488 6996
rect 8484 6944 8536 6996
rect 9496 6944 9548 6996
rect 13820 6944 13872 6996
rect 4804 6851 4856 6860
rect 4804 6817 4813 6851
rect 4813 6817 4847 6851
rect 4847 6817 4856 6851
rect 4804 6808 4856 6817
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 8208 6876 8260 6928
rect 6736 6808 6788 6860
rect 7932 6851 7984 6860
rect 4896 6740 4948 6792
rect 7932 6817 7941 6851
rect 7941 6817 7975 6851
rect 7975 6817 7984 6851
rect 7932 6808 7984 6817
rect 9404 6808 9456 6860
rect 4620 6672 4672 6724
rect 9220 6740 9272 6792
rect 9956 6851 10008 6860
rect 9956 6817 9965 6851
rect 9965 6817 9999 6851
rect 9999 6817 10008 6851
rect 9956 6808 10008 6817
rect 15108 6876 15160 6928
rect 11980 6851 12032 6860
rect 10416 6740 10468 6792
rect 11980 6817 11989 6851
rect 11989 6817 12023 6851
rect 12023 6817 12032 6851
rect 11980 6808 12032 6817
rect 16764 6808 16816 6860
rect 14556 6740 14608 6792
rect 10140 6715 10192 6724
rect 4988 6647 5040 6656
rect 4988 6613 4997 6647
rect 4997 6613 5031 6647
rect 5031 6613 5040 6647
rect 4988 6604 5040 6613
rect 5080 6604 5132 6656
rect 5908 6604 5960 6656
rect 7564 6647 7616 6656
rect 7564 6613 7573 6647
rect 7573 6613 7607 6647
rect 7607 6613 7616 6647
rect 7564 6604 7616 6613
rect 8116 6647 8168 6656
rect 8116 6613 8125 6647
rect 8125 6613 8159 6647
rect 8159 6613 8168 6647
rect 8116 6604 8168 6613
rect 8668 6647 8720 6656
rect 8668 6613 8677 6647
rect 8677 6613 8711 6647
rect 8711 6613 8720 6647
rect 8668 6604 8720 6613
rect 10140 6681 10149 6715
rect 10149 6681 10183 6715
rect 10183 6681 10192 6715
rect 10140 6672 10192 6681
rect 12164 6715 12216 6724
rect 12164 6681 12173 6715
rect 12173 6681 12207 6715
rect 12207 6681 12216 6715
rect 12164 6672 12216 6681
rect 9680 6604 9732 6656
rect 11612 6647 11664 6656
rect 11612 6613 11621 6647
rect 11621 6613 11655 6647
rect 11655 6613 11664 6647
rect 11612 6604 11664 6613
rect 12716 6647 12768 6656
rect 12716 6613 12725 6647
rect 12725 6613 12759 6647
rect 12759 6613 12768 6647
rect 12716 6604 12768 6613
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 4804 6400 4856 6452
rect 8668 6400 8720 6452
rect 4344 6239 4396 6248
rect 4344 6205 4353 6239
rect 4353 6205 4387 6239
rect 4387 6205 4396 6239
rect 4344 6196 4396 6205
rect 7840 6264 7892 6316
rect 8024 6332 8076 6384
rect 9864 6400 9916 6452
rect 11980 6400 12032 6452
rect 14280 6400 14332 6452
rect 9496 6332 9548 6384
rect 9956 6332 10008 6384
rect 14188 6332 14240 6384
rect 7748 6239 7800 6248
rect 7748 6205 7757 6239
rect 7757 6205 7791 6239
rect 7791 6205 7800 6239
rect 7748 6196 7800 6205
rect 7932 6196 7984 6248
rect 9404 6239 9456 6248
rect 9404 6205 9413 6239
rect 9413 6205 9447 6239
rect 9447 6205 9456 6239
rect 9404 6196 9456 6205
rect 14648 6264 14700 6316
rect 14372 6196 14424 6248
rect 6552 6128 6604 6180
rect 7380 6128 7432 6180
rect 1400 6060 1452 6112
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 5356 6103 5408 6112
rect 5356 6069 5365 6103
rect 5365 6069 5399 6103
rect 5399 6069 5408 6103
rect 5356 6060 5408 6069
rect 8208 6060 8260 6112
rect 9772 6060 9824 6112
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 7748 5788 7800 5840
rect 11888 5856 11940 5908
rect 9404 5788 9456 5840
rect 14096 5788 14148 5840
rect 9036 5720 9088 5772
rect 10600 5720 10652 5772
rect 5632 5652 5684 5704
rect 10508 5652 10560 5704
rect 7012 5584 7064 5636
rect 4436 5516 4488 5568
rect 7840 5516 7892 5568
rect 11612 5516 11664 5568
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 10324 4700 10376 4752
rect 15476 4700 15528 4752
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 9588 4156 9640 4208
rect 5264 4088 5316 4140
rect 9496 4088 9548 4140
rect 6276 4020 6328 4072
rect 10416 4020 10468 4072
rect 14280 4088 14332 4140
rect 16304 4088 16356 4140
rect 12900 4020 12952 4072
rect 13728 4020 13780 4072
rect 15936 4020 15988 4072
rect 3148 3952 3200 4004
rect 7564 3952 7616 4004
rect 7656 3952 7708 4004
rect 9956 3952 10008 4004
rect 3976 3884 4028 3936
rect 8116 3884 8168 3936
rect 9312 3884 9364 3936
rect 11244 3884 11296 3936
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 5540 3680 5592 3732
rect 9128 3680 9180 3732
rect 6920 3612 6972 3664
rect 9496 3612 9548 3664
rect 8760 3544 8812 3596
rect 11612 3544 11664 3596
rect 10692 3476 10744 3528
rect 13176 3476 13228 3528
rect 2320 3408 2372 3460
rect 4620 3408 4672 3460
rect 6552 3408 6604 3460
rect 9680 3408 9732 3460
rect 572 3340 624 3392
rect 4988 3340 5040 3392
rect 8208 3340 8260 3392
rect 12716 3340 12768 3392
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 7104 3136 7156 3188
rect 10692 3136 10744 3188
rect 204 3068 256 3120
rect 1400 3068 1452 3120
rect 1860 3068 1912 3120
rect 5356 3068 5408 3120
rect 8852 3068 8904 3120
rect 12072 3068 12124 3120
rect 2688 3000 2740 3052
rect 4896 3000 4948 3052
rect 10048 3000 10100 3052
rect 12532 3000 12584 3052
rect 1124 2932 1176 2984
rect 2964 2932 3016 2984
rect 1032 2864 1084 2916
rect 4528 2864 4580 2916
rect 1400 2796 1452 2848
rect 5080 2796 5132 2848
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 3608 1436 3660 1488
rect 7932 1436 7984 1488
rect 14004 552 14056 604
rect 14648 552 14700 604
<< metal2 >>
rect 202 19520 258 20000
rect 570 19520 626 20000
rect 1030 19520 1086 20000
rect 1398 19520 1454 20000
rect 1858 19520 1914 20000
rect 2226 19520 2282 20000
rect 2686 19520 2742 20000
rect 3054 19520 3110 20000
rect 3514 19520 3570 20000
rect 3882 19520 3938 20000
rect 4342 19520 4398 20000
rect 4710 19520 4766 20000
rect 5170 19520 5226 20000
rect 5538 19520 5594 20000
rect 5998 19520 6054 20000
rect 6366 19520 6422 20000
rect 6826 19520 6882 20000
rect 7194 19520 7250 20000
rect 7654 19520 7710 20000
rect 8022 19520 8078 20000
rect 8482 19520 8538 20000
rect 8850 19520 8906 20000
rect 9310 19520 9366 20000
rect 9678 19520 9734 20000
rect 10138 19520 10194 20000
rect 10506 19520 10562 20000
rect 10966 19520 11022 20000
rect 11334 19520 11390 20000
rect 11794 19520 11850 20000
rect 12162 19520 12218 20000
rect 12622 19520 12678 20000
rect 12990 19520 13046 20000
rect 13450 19520 13506 20000
rect 13818 19520 13874 20000
rect 14278 19520 14334 20000
rect 14646 19520 14702 20000
rect 15106 19520 15162 20000
rect 15474 19520 15530 20000
rect 15934 19520 15990 20000
rect 16302 19520 16358 20000
rect 16762 19520 16818 20000
rect 216 15366 244 19520
rect 204 15360 256 15366
rect 204 15302 256 15308
rect 584 15162 612 19520
rect 1044 15502 1072 19520
rect 1412 15706 1440 19520
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 1032 15496 1084 15502
rect 1032 15438 1084 15444
rect 572 15156 624 15162
rect 572 15098 624 15104
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1596 10198 1624 10542
rect 1584 10192 1636 10198
rect 1584 10134 1636 10140
rect 1596 8401 1624 10134
rect 1582 8392 1638 8401
rect 1582 8327 1638 8336
rect 1872 7206 1900 19520
rect 2240 15434 2268 19520
rect 2228 15428 2280 15434
rect 2228 15370 2280 15376
rect 2700 7818 2728 19520
rect 3068 16250 3096 19520
rect 3528 17626 3556 19520
rect 3790 18320 3846 18329
rect 3790 18255 3846 18264
rect 3344 17598 3556 17626
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 3344 15978 3372 17598
rect 3421 17436 3717 17456
rect 3477 17434 3501 17436
rect 3557 17434 3581 17436
rect 3637 17434 3661 17436
rect 3499 17382 3501 17434
rect 3563 17382 3575 17434
rect 3637 17382 3639 17434
rect 3477 17380 3501 17382
rect 3557 17380 3581 17382
rect 3637 17380 3661 17382
rect 3421 17360 3717 17380
rect 3421 16348 3717 16368
rect 3477 16346 3501 16348
rect 3557 16346 3581 16348
rect 3637 16346 3661 16348
rect 3499 16294 3501 16346
rect 3563 16294 3575 16346
rect 3637 16294 3639 16346
rect 3477 16292 3501 16294
rect 3557 16292 3581 16294
rect 3637 16292 3661 16294
rect 3421 16272 3717 16292
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 10198 2820 14991
rect 2884 13394 2912 15302
rect 3421 15260 3717 15280
rect 3477 15258 3501 15260
rect 3557 15258 3581 15260
rect 3637 15258 3661 15260
rect 3499 15206 3501 15258
rect 3563 15206 3575 15258
rect 3637 15206 3639 15258
rect 3477 15204 3501 15206
rect 3557 15204 3581 15206
rect 3637 15204 3661 15206
rect 3421 15184 3717 15204
rect 3421 14172 3717 14192
rect 3477 14170 3501 14172
rect 3557 14170 3581 14172
rect 3637 14170 3661 14172
rect 3499 14118 3501 14170
rect 3563 14118 3575 14170
rect 3637 14118 3639 14170
rect 3477 14116 3501 14118
rect 3557 14116 3581 14118
rect 3637 14116 3661 14118
rect 3421 14096 3717 14116
rect 3804 13938 3832 18255
rect 3896 16046 3924 19520
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 4356 13954 4384 19520
rect 4724 15910 4752 19520
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4724 15162 4752 15642
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 3792 13932 3844 13938
rect 4356 13926 4476 13954
rect 3792 13874 3844 13880
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 4356 13530 4384 13806
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3344 10606 3372 13126
rect 3421 13084 3717 13104
rect 3477 13082 3501 13084
rect 3557 13082 3581 13084
rect 3637 13082 3661 13084
rect 3499 13030 3501 13082
rect 3563 13030 3575 13082
rect 3637 13030 3639 13082
rect 3477 13028 3501 13030
rect 3557 13028 3581 13030
rect 3637 13028 3661 13030
rect 3421 13008 3717 13028
rect 3421 11996 3717 12016
rect 3477 11994 3501 11996
rect 3557 11994 3581 11996
rect 3637 11994 3661 11996
rect 3499 11942 3501 11994
rect 3563 11942 3575 11994
rect 3637 11942 3639 11994
rect 3477 11940 3501 11942
rect 3557 11940 3581 11942
rect 3637 11940 3661 11942
rect 3421 11920 3717 11940
rect 4066 11656 4122 11665
rect 4066 11591 4122 11600
rect 3421 10908 3717 10928
rect 3477 10906 3501 10908
rect 3557 10906 3581 10908
rect 3637 10906 3661 10908
rect 3499 10854 3501 10906
rect 3563 10854 3575 10906
rect 3637 10854 3639 10906
rect 3477 10852 3501 10854
rect 3557 10852 3581 10854
rect 3637 10852 3661 10854
rect 3421 10832 3717 10852
rect 4080 10674 4108 11591
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 572 3392 624 3398
rect 572 3334 624 3340
rect 204 3120 256 3126
rect 204 3062 256 3068
rect 216 480 244 3062
rect 584 480 612 3334
rect 1412 3126 1440 6054
rect 2320 3460 2372 3466
rect 2320 3402 2372 3408
rect 1400 3120 1452 3126
rect 1400 3062 1452 3068
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 1124 2984 1176 2990
rect 1124 2926 1176 2932
rect 1032 2916 1084 2922
rect 1032 2858 1084 2864
rect 1044 480 1072 2858
rect 1136 1737 1164 2926
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1122 1728 1178 1737
rect 1122 1663 1178 1672
rect 1412 480 1440 2790
rect 1872 480 1900 3062
rect 2332 480 2360 3402
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2700 480 2728 2994
rect 2976 2990 3004 9930
rect 3421 9820 3717 9840
rect 3477 9818 3501 9820
rect 3557 9818 3581 9820
rect 3637 9818 3661 9820
rect 3499 9766 3501 9818
rect 3563 9766 3575 9818
rect 3637 9766 3639 9818
rect 3477 9764 3501 9766
rect 3557 9764 3581 9766
rect 3637 9764 3661 9766
rect 3421 9744 3717 9764
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 3421 8732 3717 8752
rect 3477 8730 3501 8732
rect 3557 8730 3581 8732
rect 3637 8730 3661 8732
rect 3499 8678 3501 8730
rect 3563 8678 3575 8730
rect 3637 8678 3639 8730
rect 3477 8676 3501 8678
rect 3557 8676 3581 8678
rect 3637 8676 3661 8678
rect 3421 8656 3717 8676
rect 3421 7644 3717 7664
rect 3477 7642 3501 7644
rect 3557 7642 3581 7644
rect 3637 7642 3661 7644
rect 3499 7590 3501 7642
rect 3563 7590 3575 7642
rect 3637 7590 3639 7642
rect 3477 7588 3501 7590
rect 3557 7588 3581 7590
rect 3637 7588 3661 7590
rect 3421 7568 3717 7588
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 3068 5001 3096 7210
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 4356 6254 4384 9386
rect 4448 7002 4476 13926
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 4816 6866 4844 16390
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 5092 7546 5120 15438
rect 5184 7750 5212 19520
rect 5552 16182 5580 19520
rect 6012 17082 6040 19520
rect 6012 17054 6316 17082
rect 5886 16892 6182 16912
rect 5942 16890 5966 16892
rect 6022 16890 6046 16892
rect 6102 16890 6126 16892
rect 5964 16838 5966 16890
rect 6028 16838 6040 16890
rect 6102 16838 6104 16890
rect 5942 16836 5966 16838
rect 6022 16836 6046 16838
rect 6102 16836 6126 16838
rect 5886 16816 6182 16836
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5552 15162 5580 15370
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5644 7478 5672 15982
rect 5886 15804 6182 15824
rect 5942 15802 5966 15804
rect 6022 15802 6046 15804
rect 6102 15802 6126 15804
rect 5964 15750 5966 15802
rect 6028 15750 6040 15802
rect 6102 15750 6104 15802
rect 5942 15748 5966 15750
rect 6022 15748 6046 15750
rect 6102 15748 6126 15750
rect 5886 15728 6182 15748
rect 6288 15706 6316 17054
rect 6380 16114 6408 19520
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6368 15972 6420 15978
rect 6368 15914 6420 15920
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 5886 14716 6182 14736
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6126 14716
rect 5964 14662 5966 14714
rect 6028 14662 6040 14714
rect 6102 14662 6104 14714
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6126 14662
rect 5886 14640 6182 14660
rect 5886 13628 6182 13648
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6126 13628
rect 5964 13574 5966 13626
rect 6028 13574 6040 13626
rect 6102 13574 6104 13626
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6126 13574
rect 5886 13552 6182 13572
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 5886 12540 6182 12560
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6126 12540
rect 5964 12486 5966 12538
rect 6028 12486 6040 12538
rect 6102 12486 6104 12538
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6126 12486
rect 5886 12464 6182 12484
rect 5886 11452 6182 11472
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6126 11452
rect 5964 11398 5966 11450
rect 6028 11398 6040 11450
rect 6102 11398 6104 11450
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6126 11398
rect 5886 11376 6182 11396
rect 6288 11286 6316 12582
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 5886 10364 6182 10384
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6126 10364
rect 5964 10310 5966 10362
rect 6028 10310 6040 10362
rect 6102 10310 6104 10362
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6126 10310
rect 5886 10288 6182 10308
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 5886 9276 6182 9296
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6126 9276
rect 5964 9222 5966 9274
rect 6028 9222 6040 9274
rect 6102 9222 6104 9274
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6126 9222
rect 5886 9200 6182 9220
rect 5886 8188 6182 8208
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6126 8188
rect 5964 8134 5966 8186
rect 6028 8134 6040 8186
rect 6102 8134 6104 8186
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6126 8134
rect 5886 8112 6182 8132
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 6288 7410 6316 9862
rect 6380 7970 6408 15914
rect 6472 8090 6500 16186
rect 6840 16046 6868 19520
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 15162 6868 15846
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6564 11626 6592 14826
rect 6748 12782 6776 14962
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6656 11694 6684 12378
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6656 11506 6684 11630
rect 6564 11478 6684 11506
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6380 7942 6500 7970
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6380 7546 6408 7754
rect 6472 7546 6500 7942
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 3054 4992 3110 5001
rect 3054 4927 3110 4936
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 3160 480 3188 3946
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3421 3292 3717 3312
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3421 2128 3717 2148
rect 3608 1488 3660 1494
rect 3608 1430 3660 1436
rect 3620 480 3648 1430
rect 3988 480 4016 3878
rect 4448 480 4476 5510
rect 4540 2922 4568 6054
rect 4632 3466 4660 6666
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4528 2916 4580 2922
rect 4528 2858 4580 2864
rect 4816 480 4844 6394
rect 4908 3058 4936 6734
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5000 3398 5028 6598
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 5092 2854 5120 6598
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5276 480 5304 4082
rect 5368 3126 5396 6054
rect 5552 3738 5580 7278
rect 5886 7100 6182 7120
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6126 7100
rect 5964 7046 5966 7098
rect 6028 7046 6040 7098
rect 6102 7046 6104 7098
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6126 7046
rect 5886 7024 6182 7044
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5644 5710 5672 6802
rect 5908 6656 5960 6662
rect 5736 6616 5908 6644
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 5736 480 5764 6616
rect 5908 6598 5960 6604
rect 6564 6186 6592 11478
rect 6748 11354 6776 11494
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6748 6866 6776 10406
rect 6932 9654 6960 12718
rect 7024 12714 7052 15370
rect 7208 15366 7236 19520
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 7024 9654 7052 12650
rect 7208 12102 7236 13330
rect 7392 12850 7420 13942
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7392 12730 7420 12786
rect 7300 12702 7420 12730
rect 7300 12170 7328 12702
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7116 9654 7144 11018
rect 7208 10606 7236 12038
rect 7300 11830 7328 12106
rect 7288 11824 7340 11830
rect 7340 11772 7420 11778
rect 7288 11766 7420 11772
rect 7300 11750 7420 11766
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7300 11218 7328 11630
rect 7392 11286 7420 11750
rect 7668 11558 7696 19520
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7300 10742 7328 11154
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7300 10130 7328 10678
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 5886 3836 6182 3856
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 6288 1850 6316 4014
rect 6932 3670 6960 9454
rect 7208 9382 7236 10066
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7484 7886 7512 11494
rect 7852 10690 7880 15982
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 7668 10662 7880 10690
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7668 7818 7696 10662
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7760 10198 7788 10542
rect 7748 10192 7800 10198
rect 7800 10140 7880 10146
rect 7748 10134 7880 10140
rect 7760 10118 7880 10134
rect 7852 9586 7880 10118
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6104 1822 6316 1850
rect 6104 480 6132 1822
rect 6564 480 6592 3402
rect 7024 480 7052 5578
rect 7116 3194 7144 7278
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7392 480 7420 6122
rect 7576 4010 7604 6598
rect 7668 4010 7696 7210
rect 7944 6866 7972 15914
rect 8036 15910 8064 19520
rect 8496 17626 8524 19520
rect 8496 17598 8708 17626
rect 8352 17436 8648 17456
rect 8408 17434 8432 17436
rect 8488 17434 8512 17436
rect 8568 17434 8592 17436
rect 8430 17382 8432 17434
rect 8494 17382 8506 17434
rect 8568 17382 8570 17434
rect 8408 17380 8432 17382
rect 8488 17380 8512 17382
rect 8568 17380 8592 17382
rect 8352 17360 8648 17380
rect 8352 16348 8648 16368
rect 8408 16346 8432 16348
rect 8488 16346 8512 16348
rect 8568 16346 8592 16348
rect 8430 16294 8432 16346
rect 8494 16294 8506 16346
rect 8568 16294 8570 16346
rect 8408 16292 8432 16294
rect 8488 16292 8512 16294
rect 8568 16292 8592 16294
rect 8352 16272 8648 16292
rect 8208 16176 8260 16182
rect 8208 16118 8260 16124
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 8024 14884 8076 14890
rect 8024 14826 8076 14832
rect 8036 12238 8064 14826
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8036 11898 8064 12174
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 8036 9926 8064 11562
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8128 7478 8156 16050
rect 8220 7546 8248 16118
rect 8680 16046 8708 17598
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8352 15260 8648 15280
rect 8408 15258 8432 15260
rect 8488 15258 8512 15260
rect 8568 15258 8592 15260
rect 8430 15206 8432 15258
rect 8494 15206 8506 15258
rect 8568 15206 8570 15258
rect 8408 15204 8432 15206
rect 8488 15204 8512 15206
rect 8568 15204 8592 15206
rect 8352 15184 8648 15204
rect 8352 14172 8648 14192
rect 8408 14170 8432 14172
rect 8488 14170 8512 14172
rect 8568 14170 8592 14172
rect 8430 14118 8432 14170
rect 8494 14118 8506 14170
rect 8568 14118 8570 14170
rect 8408 14116 8432 14118
rect 8488 14116 8512 14118
rect 8568 14116 8592 14118
rect 8352 14096 8648 14116
rect 8352 13084 8648 13104
rect 8408 13082 8432 13084
rect 8488 13082 8512 13084
rect 8568 13082 8592 13084
rect 8430 13030 8432 13082
rect 8494 13030 8506 13082
rect 8568 13030 8570 13082
rect 8408 13028 8432 13030
rect 8488 13028 8512 13030
rect 8568 13028 8592 13030
rect 8352 13008 8648 13028
rect 8864 12442 8892 19520
rect 9324 16454 9352 19520
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8352 11996 8648 12016
rect 8408 11994 8432 11996
rect 8488 11994 8512 11996
rect 8568 11994 8592 11996
rect 8430 11942 8432 11994
rect 8494 11942 8506 11994
rect 8568 11942 8570 11994
rect 8408 11940 8432 11942
rect 8488 11940 8512 11942
rect 8568 11940 8592 11942
rect 8352 11920 8648 11940
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8352 10908 8648 10928
rect 8408 10906 8432 10908
rect 8488 10906 8512 10908
rect 8568 10906 8592 10908
rect 8430 10854 8432 10906
rect 8494 10854 8506 10906
rect 8568 10854 8570 10906
rect 8408 10852 8432 10854
rect 8488 10852 8512 10854
rect 8568 10852 8592 10854
rect 8352 10832 8648 10852
rect 8680 10538 8708 10950
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8352 9820 8648 9840
rect 8408 9818 8432 9820
rect 8488 9818 8512 9820
rect 8568 9818 8592 9820
rect 8430 9766 8432 9818
rect 8494 9766 8506 9818
rect 8568 9766 8570 9818
rect 8408 9764 8432 9766
rect 8488 9764 8512 9766
rect 8568 9764 8592 9766
rect 8352 9744 8648 9764
rect 8680 9654 8708 10474
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8772 9586 8800 12038
rect 8956 11642 8984 14894
rect 8864 11614 8984 11642
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8864 9382 8892 11614
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8352 8732 8648 8752
rect 8408 8730 8432 8732
rect 8488 8730 8512 8732
rect 8568 8730 8592 8732
rect 8430 8678 8432 8730
rect 8494 8678 8506 8730
rect 8568 8678 8570 8730
rect 8408 8676 8432 8678
rect 8488 8676 8512 8678
rect 8568 8676 8592 8678
rect 8352 8656 8648 8676
rect 8352 7644 8648 7664
rect 8408 7642 8432 7644
rect 8488 7642 8512 7644
rect 8568 7642 8592 7644
rect 8430 7590 8432 7642
rect 8494 7590 8506 7642
rect 8568 7590 8570 7642
rect 8408 7588 8432 7590
rect 8488 7588 8512 7590
rect 8568 7588 8592 7590
rect 8352 7568 8648 7588
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8024 6384 8076 6390
rect 7852 6332 8024 6338
rect 7852 6326 8076 6332
rect 7852 6322 8064 6326
rect 7840 6316 8064 6322
rect 7892 6310 8064 6316
rect 7840 6258 7892 6264
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7760 5846 7788 6190
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7852 480 7880 5510
rect 7944 1494 7972 6190
rect 8128 3942 8156 6598
rect 8220 6118 8248 6870
rect 8312 6746 8340 7142
rect 8496 7002 8524 7142
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8312 6718 8800 6746
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8352 6480 8648 6500
rect 8680 6458 8708 6598
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8352 5392 8648 5412
rect 8352 4380 8648 4400
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8772 3602 8800 6718
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 7932 1488 7984 1494
rect 7932 1430 7984 1436
rect 8220 480 8248 3334
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8352 3216 8648 3236
rect 8864 3126 8892 7210
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 8956 2938 8984 11494
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9048 5778 9076 11086
rect 9140 10470 9168 16186
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9404 15632 9456 15638
rect 9404 15574 9456 15580
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9232 12646 9260 13262
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9232 11898 9260 12582
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9324 10554 9352 15438
rect 9232 10526 9352 10554
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 7206 9168 7686
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9232 6798 9260 10526
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 10266 9352 10406
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9324 3942 9352 7890
rect 9416 6866 9444 15574
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9508 15162 9536 15302
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9508 7562 9536 9318
rect 9600 7750 9628 15982
rect 9692 15434 9720 19520
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9692 10674 9720 10950
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9508 7534 9628 7562
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9508 7002 9536 7278
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9416 5846 9444 6190
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 9508 4146 9536 6326
rect 9600 4214 9628 7534
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 8772 2910 8984 2938
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 8772 898 8800 2910
rect 8680 870 8800 898
rect 8680 480 8708 870
rect 9140 480 9168 3674
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9508 480 9536 3606
rect 9692 3466 9720 6598
rect 9784 6118 9812 17002
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9876 12730 9904 14894
rect 10060 12866 10088 15642
rect 10152 13002 10180 19520
rect 10152 12974 10272 13002
rect 10060 12838 10180 12866
rect 9876 12702 10088 12730
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9876 6458 9904 12242
rect 10060 11218 10088 12702
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9968 6390 9996 6802
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9968 480 9996 3946
rect 10060 3058 10088 7346
rect 10152 6730 10180 12838
rect 10244 11914 10272 12974
rect 10520 12306 10548 19520
rect 10980 17066 11008 19520
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10817 16892 11113 16912
rect 10873 16890 10897 16892
rect 10953 16890 10977 16892
rect 11033 16890 11057 16892
rect 10895 16838 10897 16890
rect 10959 16838 10971 16890
rect 11033 16838 11035 16890
rect 10873 16836 10897 16838
rect 10953 16836 10977 16838
rect 11033 16836 11057 16838
rect 10817 16816 11113 16836
rect 11348 16250 11376 19520
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 10817 15804 11113 15824
rect 10873 15802 10897 15804
rect 10953 15802 10977 15804
rect 11033 15802 11057 15804
rect 10895 15750 10897 15802
rect 10959 15750 10971 15802
rect 11033 15750 11035 15802
rect 10873 15748 10897 15750
rect 10953 15748 10977 15750
rect 11033 15748 11057 15750
rect 10817 15728 11113 15748
rect 10817 14716 11113 14736
rect 10873 14714 10897 14716
rect 10953 14714 10977 14716
rect 11033 14714 11057 14716
rect 10895 14662 10897 14714
rect 10959 14662 10971 14714
rect 11033 14662 11035 14714
rect 10873 14660 10897 14662
rect 10953 14660 10977 14662
rect 11033 14660 11057 14662
rect 10817 14640 11113 14660
rect 10817 13628 11113 13648
rect 10873 13626 10897 13628
rect 10953 13626 10977 13628
rect 11033 13626 11057 13628
rect 10895 13574 10897 13626
rect 10959 13574 10971 13626
rect 11033 13574 11035 13626
rect 10873 13572 10897 13574
rect 10953 13572 10977 13574
rect 11033 13572 11057 13574
rect 10817 13552 11113 13572
rect 10817 12540 11113 12560
rect 10873 12538 10897 12540
rect 10953 12538 10977 12540
rect 11033 12538 11057 12540
rect 10895 12486 10897 12538
rect 10959 12486 10971 12538
rect 11033 12486 11035 12538
rect 10873 12484 10897 12486
rect 10953 12484 10977 12486
rect 11033 12484 11057 12486
rect 10817 12464 11113 12484
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10244 11886 10548 11914
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10244 2802 10272 11766
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10336 4758 10364 11154
rect 10414 9480 10470 9489
rect 10414 9415 10470 9424
rect 10428 6798 10456 9415
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10428 4078 10456 6054
rect 10520 5710 10548 11886
rect 10817 11452 11113 11472
rect 10873 11450 10897 11452
rect 10953 11450 10977 11452
rect 11033 11450 11057 11452
rect 10895 11398 10897 11450
rect 10959 11398 10971 11450
rect 11033 11398 11035 11450
rect 10873 11396 10897 11398
rect 10953 11396 10977 11398
rect 11033 11396 11057 11398
rect 10817 11376 11113 11396
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10888 10674 10916 11018
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10612 5778 10640 10542
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10704 10266 10732 10406
rect 10817 10364 11113 10384
rect 10873 10362 10897 10364
rect 10953 10362 10977 10364
rect 11033 10362 11057 10364
rect 10895 10310 10897 10362
rect 10959 10310 10971 10362
rect 11033 10310 11035 10362
rect 10873 10308 10897 10310
rect 10953 10308 10977 10310
rect 11033 10308 11057 10310
rect 10817 10288 11113 10308
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10817 9276 11113 9296
rect 10873 9274 10897 9276
rect 10953 9274 10977 9276
rect 11033 9274 11057 9276
rect 10895 9222 10897 9274
rect 10959 9222 10971 9274
rect 11033 9222 11035 9274
rect 10873 9220 10897 9222
rect 10953 9220 10977 9222
rect 11033 9220 11057 9222
rect 10817 9200 11113 9220
rect 11164 8974 11192 12310
rect 11808 9761 11836 19520
rect 12176 15994 12204 19520
rect 12084 15966 12204 15994
rect 12636 15978 12664 19520
rect 12624 15972 12676 15978
rect 12084 12356 12112 15966
rect 12624 15914 12676 15920
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 11992 12328 12112 12356
rect 11794 9752 11850 9761
rect 11794 9687 11850 9696
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 10817 8188 11113 8208
rect 10873 8186 10897 8188
rect 10953 8186 10977 8188
rect 11033 8186 11057 8188
rect 10895 8134 10897 8186
rect 10959 8134 10971 8186
rect 11033 8134 11035 8186
rect 10873 8132 10897 8134
rect 10953 8132 10977 8134
rect 11033 8132 11057 8134
rect 10817 8112 11113 8132
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10980 7546 11008 7754
rect 11808 7546 11836 7822
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10704 3534 10732 7210
rect 10817 7100 11113 7120
rect 10873 7098 10897 7100
rect 10953 7098 10977 7100
rect 11033 7098 11057 7100
rect 10895 7046 10897 7098
rect 10959 7046 10971 7098
rect 11033 7046 11035 7098
rect 10873 7044 10897 7046
rect 10953 7044 10977 7046
rect 11033 7044 11057 7046
rect 10817 7024 11113 7044
rect 11992 7018 12020 12328
rect 11900 6990 12020 7018
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 11624 5574 11652 6598
rect 11900 5914 11928 6990
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11992 6458 12020 6802
rect 12176 6730 12204 15846
rect 13004 11354 13032 19520
rect 13464 17626 13492 19520
rect 13188 17598 13492 17626
rect 13188 15502 13216 17598
rect 13726 17504 13782 17513
rect 13282 17436 13578 17456
rect 13726 17439 13782 17448
rect 13338 17434 13362 17436
rect 13418 17434 13442 17436
rect 13498 17434 13522 17436
rect 13360 17382 13362 17434
rect 13424 17382 13436 17434
rect 13498 17382 13500 17434
rect 13338 17380 13362 17382
rect 13418 17380 13442 17382
rect 13498 17380 13522 17382
rect 13282 17360 13578 17380
rect 13282 16348 13578 16368
rect 13338 16346 13362 16348
rect 13418 16346 13442 16348
rect 13498 16346 13522 16348
rect 13360 16294 13362 16346
rect 13424 16294 13436 16346
rect 13498 16294 13500 16346
rect 13338 16292 13362 16294
rect 13418 16292 13442 16294
rect 13498 16292 13522 16294
rect 13282 16272 13578 16292
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13282 15260 13578 15280
rect 13338 15258 13362 15260
rect 13418 15258 13442 15260
rect 13498 15258 13522 15260
rect 13360 15206 13362 15258
rect 13424 15206 13436 15258
rect 13498 15206 13500 15258
rect 13338 15204 13362 15206
rect 13418 15204 13442 15206
rect 13498 15204 13522 15206
rect 13282 15184 13578 15204
rect 13282 14172 13578 14192
rect 13338 14170 13362 14172
rect 13418 14170 13442 14172
rect 13498 14170 13522 14172
rect 13360 14118 13362 14170
rect 13424 14118 13436 14170
rect 13498 14118 13500 14170
rect 13338 14116 13362 14118
rect 13418 14116 13442 14118
rect 13498 14116 13522 14118
rect 13282 14096 13578 14116
rect 13740 13530 13768 17439
rect 13832 15994 13860 19520
rect 13832 15966 14136 15994
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13282 13084 13578 13104
rect 13338 13082 13362 13084
rect 13418 13082 13442 13084
rect 13498 13082 13522 13084
rect 13360 13030 13362 13082
rect 13424 13030 13436 13082
rect 13498 13030 13500 13082
rect 13338 13028 13362 13030
rect 13418 13028 13442 13030
rect 13498 13028 13522 13030
rect 13282 13008 13578 13028
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13740 12481 13768 12582
rect 13726 12472 13782 12481
rect 13726 12407 13782 12416
rect 13282 11996 13578 12016
rect 13338 11994 13362 11996
rect 13418 11994 13442 11996
rect 13498 11994 13522 11996
rect 13360 11942 13362 11994
rect 13424 11942 13436 11994
rect 13498 11942 13500 11994
rect 13338 11940 13362 11942
rect 13418 11940 13442 11942
rect 13498 11940 13522 11942
rect 13282 11920 13578 11940
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13282 10908 13578 10928
rect 13338 10906 13362 10908
rect 13418 10906 13442 10908
rect 13498 10906 13522 10908
rect 13360 10854 13362 10906
rect 13424 10854 13436 10906
rect 13498 10854 13500 10906
rect 13338 10852 13362 10854
rect 13418 10852 13442 10854
rect 13498 10852 13522 10854
rect 13282 10832 13578 10852
rect 13832 10810 13860 13126
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13282 9820 13578 9840
rect 13338 9818 13362 9820
rect 13418 9818 13442 9820
rect 13498 9818 13522 9820
rect 13360 9766 13362 9818
rect 13424 9766 13436 9818
rect 13498 9766 13500 9818
rect 13338 9764 13362 9766
rect 13418 9764 13442 9766
rect 13498 9764 13522 9766
rect 13282 9744 13578 9764
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12544 7449 12572 8978
rect 13282 8732 13578 8752
rect 13338 8730 13362 8732
rect 13418 8730 13442 8732
rect 13498 8730 13522 8732
rect 13360 8678 13362 8730
rect 13424 8678 13436 8730
rect 13498 8678 13500 8730
rect 13338 8676 13362 8678
rect 13418 8676 13442 8678
rect 13498 8676 13522 8678
rect 13282 8656 13578 8676
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12636 7546 12664 7686
rect 13282 7644 13578 7664
rect 13338 7642 13362 7644
rect 13418 7642 13442 7644
rect 13498 7642 13522 7644
rect 13360 7590 13362 7642
rect 13424 7590 13436 7642
rect 13498 7590 13500 7642
rect 13338 7588 13362 7590
rect 13418 7588 13442 7590
rect 13498 7588 13522 7590
rect 13282 7568 13578 7588
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12530 7440 12586 7449
rect 12530 7375 12586 7384
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10817 4848 11113 4868
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10244 2774 10364 2802
rect 10336 2666 10364 2774
rect 10336 2638 10456 2666
rect 10428 480 10456 2638
rect 10704 2530 10732 3130
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10817 2672 11113 2692
rect 10704 2502 10824 2530
rect 10796 480 10824 2502
rect 11256 480 11284 3878
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11624 480 11652 3538
rect 12728 3398 12756 6598
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13282 4380 13578 4400
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12084 480 12112 3062
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12544 480 12572 2994
rect 12912 480 12940 4014
rect 13648 3890 13676 10746
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13740 4078 13768 7210
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13648 3862 13768 3890
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13188 1986 13216 3470
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 13740 2553 13768 3862
rect 13726 2544 13782 2553
rect 13726 2479 13782 2488
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 13188 1958 13400 1986
rect 13372 480 13400 1958
rect 13832 480 13860 6938
rect 14016 610 14044 7414
rect 14108 5846 14136 15966
rect 14292 15638 14320 19520
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14280 15632 14332 15638
rect 14280 15574 14332 15580
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 14004 604 14056 610
rect 14004 546 14056 552
rect 14200 480 14228 6326
rect 14292 4146 14320 6394
rect 14384 6254 14412 15438
rect 14568 6798 14596 15982
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14660 6322 14688 19520
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14648 604 14700 610
rect 14648 546 14700 552
rect 14660 480 14688 546
rect 15028 480 15056 7346
rect 15120 6934 15148 19520
rect 15488 10606 15516 19520
rect 15948 15502 15976 19520
rect 16316 16046 16344 19520
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 16776 6866 16804 19520
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 15488 480 15516 4694
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15948 480 15976 4014
rect 16316 480 16344 4082
rect 16868 2802 16896 7278
rect 16776 2774 16896 2802
rect 16776 480 16804 2774
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1398 0 1454 480
rect 1858 0 1914 480
rect 2318 0 2374 480
rect 2686 0 2742 480
rect 3146 0 3202 480
rect 3606 0 3662 480
rect 3974 0 4030 480
rect 4434 0 4490 480
rect 4802 0 4858 480
rect 5262 0 5318 480
rect 5722 0 5778 480
rect 6090 0 6146 480
rect 6550 0 6606 480
rect 7010 0 7066 480
rect 7378 0 7434 480
rect 7838 0 7894 480
rect 8206 0 8262 480
rect 8666 0 8722 480
rect 9126 0 9182 480
rect 9494 0 9550 480
rect 9954 0 10010 480
rect 10414 0 10470 480
rect 10782 0 10838 480
rect 11242 0 11298 480
rect 11610 0 11666 480
rect 12070 0 12126 480
rect 12530 0 12586 480
rect 12898 0 12954 480
rect 13358 0 13414 480
rect 13818 0 13874 480
rect 14186 0 14242 480
rect 14646 0 14702 480
rect 15014 0 15070 480
rect 15474 0 15530 480
rect 15934 0 15990 480
rect 16302 0 16358 480
rect 16762 0 16818 480
<< via2 >>
rect 1582 8336 1638 8392
rect 3790 18264 3846 18320
rect 3421 17434 3477 17436
rect 3501 17434 3557 17436
rect 3581 17434 3637 17436
rect 3661 17434 3717 17436
rect 3421 17382 3447 17434
rect 3447 17382 3477 17434
rect 3501 17382 3511 17434
rect 3511 17382 3557 17434
rect 3581 17382 3627 17434
rect 3627 17382 3637 17434
rect 3661 17382 3691 17434
rect 3691 17382 3717 17434
rect 3421 17380 3477 17382
rect 3501 17380 3557 17382
rect 3581 17380 3637 17382
rect 3661 17380 3717 17382
rect 3421 16346 3477 16348
rect 3501 16346 3557 16348
rect 3581 16346 3637 16348
rect 3661 16346 3717 16348
rect 3421 16294 3447 16346
rect 3447 16294 3477 16346
rect 3501 16294 3511 16346
rect 3511 16294 3557 16346
rect 3581 16294 3627 16346
rect 3627 16294 3637 16346
rect 3661 16294 3691 16346
rect 3691 16294 3717 16346
rect 3421 16292 3477 16294
rect 3501 16292 3557 16294
rect 3581 16292 3637 16294
rect 3661 16292 3717 16294
rect 2778 15000 2834 15056
rect 3421 15258 3477 15260
rect 3501 15258 3557 15260
rect 3581 15258 3637 15260
rect 3661 15258 3717 15260
rect 3421 15206 3447 15258
rect 3447 15206 3477 15258
rect 3501 15206 3511 15258
rect 3511 15206 3557 15258
rect 3581 15206 3627 15258
rect 3627 15206 3637 15258
rect 3661 15206 3691 15258
rect 3691 15206 3717 15258
rect 3421 15204 3477 15206
rect 3501 15204 3557 15206
rect 3581 15204 3637 15206
rect 3661 15204 3717 15206
rect 3421 14170 3477 14172
rect 3501 14170 3557 14172
rect 3581 14170 3637 14172
rect 3661 14170 3717 14172
rect 3421 14118 3447 14170
rect 3447 14118 3477 14170
rect 3501 14118 3511 14170
rect 3511 14118 3557 14170
rect 3581 14118 3627 14170
rect 3627 14118 3637 14170
rect 3661 14118 3691 14170
rect 3691 14118 3717 14170
rect 3421 14116 3477 14118
rect 3501 14116 3557 14118
rect 3581 14116 3637 14118
rect 3661 14116 3717 14118
rect 3421 13082 3477 13084
rect 3501 13082 3557 13084
rect 3581 13082 3637 13084
rect 3661 13082 3717 13084
rect 3421 13030 3447 13082
rect 3447 13030 3477 13082
rect 3501 13030 3511 13082
rect 3511 13030 3557 13082
rect 3581 13030 3627 13082
rect 3627 13030 3637 13082
rect 3661 13030 3691 13082
rect 3691 13030 3717 13082
rect 3421 13028 3477 13030
rect 3501 13028 3557 13030
rect 3581 13028 3637 13030
rect 3661 13028 3717 13030
rect 3421 11994 3477 11996
rect 3501 11994 3557 11996
rect 3581 11994 3637 11996
rect 3661 11994 3717 11996
rect 3421 11942 3447 11994
rect 3447 11942 3477 11994
rect 3501 11942 3511 11994
rect 3511 11942 3557 11994
rect 3581 11942 3627 11994
rect 3627 11942 3637 11994
rect 3661 11942 3691 11994
rect 3691 11942 3717 11994
rect 3421 11940 3477 11942
rect 3501 11940 3557 11942
rect 3581 11940 3637 11942
rect 3661 11940 3717 11942
rect 4066 11600 4122 11656
rect 3421 10906 3477 10908
rect 3501 10906 3557 10908
rect 3581 10906 3637 10908
rect 3661 10906 3717 10908
rect 3421 10854 3447 10906
rect 3447 10854 3477 10906
rect 3501 10854 3511 10906
rect 3511 10854 3557 10906
rect 3581 10854 3627 10906
rect 3627 10854 3637 10906
rect 3661 10854 3691 10906
rect 3691 10854 3717 10906
rect 3421 10852 3477 10854
rect 3501 10852 3557 10854
rect 3581 10852 3637 10854
rect 3661 10852 3717 10854
rect 1122 1672 1178 1728
rect 3421 9818 3477 9820
rect 3501 9818 3557 9820
rect 3581 9818 3637 9820
rect 3661 9818 3717 9820
rect 3421 9766 3447 9818
rect 3447 9766 3477 9818
rect 3501 9766 3511 9818
rect 3511 9766 3557 9818
rect 3581 9766 3627 9818
rect 3627 9766 3637 9818
rect 3661 9766 3691 9818
rect 3691 9766 3717 9818
rect 3421 9764 3477 9766
rect 3501 9764 3557 9766
rect 3581 9764 3637 9766
rect 3661 9764 3717 9766
rect 3421 8730 3477 8732
rect 3501 8730 3557 8732
rect 3581 8730 3637 8732
rect 3661 8730 3717 8732
rect 3421 8678 3447 8730
rect 3447 8678 3477 8730
rect 3501 8678 3511 8730
rect 3511 8678 3557 8730
rect 3581 8678 3627 8730
rect 3627 8678 3637 8730
rect 3661 8678 3691 8730
rect 3691 8678 3717 8730
rect 3421 8676 3477 8678
rect 3501 8676 3557 8678
rect 3581 8676 3637 8678
rect 3661 8676 3717 8678
rect 3421 7642 3477 7644
rect 3501 7642 3557 7644
rect 3581 7642 3637 7644
rect 3661 7642 3717 7644
rect 3421 7590 3447 7642
rect 3447 7590 3477 7642
rect 3501 7590 3511 7642
rect 3511 7590 3557 7642
rect 3581 7590 3627 7642
rect 3627 7590 3637 7642
rect 3661 7590 3691 7642
rect 3691 7590 3717 7642
rect 3421 7588 3477 7590
rect 3501 7588 3557 7590
rect 3581 7588 3637 7590
rect 3661 7588 3717 7590
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 5886 16890 5942 16892
rect 5966 16890 6022 16892
rect 6046 16890 6102 16892
rect 6126 16890 6182 16892
rect 5886 16838 5912 16890
rect 5912 16838 5942 16890
rect 5966 16838 5976 16890
rect 5976 16838 6022 16890
rect 6046 16838 6092 16890
rect 6092 16838 6102 16890
rect 6126 16838 6156 16890
rect 6156 16838 6182 16890
rect 5886 16836 5942 16838
rect 5966 16836 6022 16838
rect 6046 16836 6102 16838
rect 6126 16836 6182 16838
rect 5886 15802 5942 15804
rect 5966 15802 6022 15804
rect 6046 15802 6102 15804
rect 6126 15802 6182 15804
rect 5886 15750 5912 15802
rect 5912 15750 5942 15802
rect 5966 15750 5976 15802
rect 5976 15750 6022 15802
rect 6046 15750 6092 15802
rect 6092 15750 6102 15802
rect 6126 15750 6156 15802
rect 6156 15750 6182 15802
rect 5886 15748 5942 15750
rect 5966 15748 6022 15750
rect 6046 15748 6102 15750
rect 6126 15748 6182 15750
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 6126 14714 6182 14716
rect 5886 14662 5912 14714
rect 5912 14662 5942 14714
rect 5966 14662 5976 14714
rect 5976 14662 6022 14714
rect 6046 14662 6092 14714
rect 6092 14662 6102 14714
rect 6126 14662 6156 14714
rect 6156 14662 6182 14714
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 6126 14660 6182 14662
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 6126 13626 6182 13628
rect 5886 13574 5912 13626
rect 5912 13574 5942 13626
rect 5966 13574 5976 13626
rect 5976 13574 6022 13626
rect 6046 13574 6092 13626
rect 6092 13574 6102 13626
rect 6126 13574 6156 13626
rect 6156 13574 6182 13626
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 6126 13572 6182 13574
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 6126 12538 6182 12540
rect 5886 12486 5912 12538
rect 5912 12486 5942 12538
rect 5966 12486 5976 12538
rect 5976 12486 6022 12538
rect 6046 12486 6092 12538
rect 6092 12486 6102 12538
rect 6126 12486 6156 12538
rect 6156 12486 6182 12538
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 6126 12484 6182 12486
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 6126 11450 6182 11452
rect 5886 11398 5912 11450
rect 5912 11398 5942 11450
rect 5966 11398 5976 11450
rect 5976 11398 6022 11450
rect 6046 11398 6092 11450
rect 6092 11398 6102 11450
rect 6126 11398 6156 11450
rect 6156 11398 6182 11450
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 6126 11396 6182 11398
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 6126 10362 6182 10364
rect 5886 10310 5912 10362
rect 5912 10310 5942 10362
rect 5966 10310 5976 10362
rect 5976 10310 6022 10362
rect 6046 10310 6092 10362
rect 6092 10310 6102 10362
rect 6126 10310 6156 10362
rect 6156 10310 6182 10362
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 6126 10308 6182 10310
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 6126 9274 6182 9276
rect 5886 9222 5912 9274
rect 5912 9222 5942 9274
rect 5966 9222 5976 9274
rect 5976 9222 6022 9274
rect 6046 9222 6092 9274
rect 6092 9222 6102 9274
rect 6126 9222 6156 9274
rect 6156 9222 6182 9274
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 6126 9220 6182 9222
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 6126 8186 6182 8188
rect 5886 8134 5912 8186
rect 5912 8134 5942 8186
rect 5966 8134 5976 8186
rect 5976 8134 6022 8186
rect 6046 8134 6092 8186
rect 6092 8134 6102 8186
rect 6126 8134 6156 8186
rect 6156 8134 6182 8186
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 6126 8132 6182 8134
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 3054 4936 3110 4992
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 6126 7098 6182 7100
rect 5886 7046 5912 7098
rect 5912 7046 5942 7098
rect 5966 7046 5976 7098
rect 5976 7046 6022 7098
rect 6046 7046 6092 7098
rect 6092 7046 6102 7098
rect 6126 7046 6156 7098
rect 6156 7046 6182 7098
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 6126 7044 6182 7046
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 8352 17434 8408 17436
rect 8432 17434 8488 17436
rect 8512 17434 8568 17436
rect 8592 17434 8648 17436
rect 8352 17382 8378 17434
rect 8378 17382 8408 17434
rect 8432 17382 8442 17434
rect 8442 17382 8488 17434
rect 8512 17382 8558 17434
rect 8558 17382 8568 17434
rect 8592 17382 8622 17434
rect 8622 17382 8648 17434
rect 8352 17380 8408 17382
rect 8432 17380 8488 17382
rect 8512 17380 8568 17382
rect 8592 17380 8648 17382
rect 8352 16346 8408 16348
rect 8432 16346 8488 16348
rect 8512 16346 8568 16348
rect 8592 16346 8648 16348
rect 8352 16294 8378 16346
rect 8378 16294 8408 16346
rect 8432 16294 8442 16346
rect 8442 16294 8488 16346
rect 8512 16294 8558 16346
rect 8558 16294 8568 16346
rect 8592 16294 8622 16346
rect 8622 16294 8648 16346
rect 8352 16292 8408 16294
rect 8432 16292 8488 16294
rect 8512 16292 8568 16294
rect 8592 16292 8648 16294
rect 8352 15258 8408 15260
rect 8432 15258 8488 15260
rect 8512 15258 8568 15260
rect 8592 15258 8648 15260
rect 8352 15206 8378 15258
rect 8378 15206 8408 15258
rect 8432 15206 8442 15258
rect 8442 15206 8488 15258
rect 8512 15206 8558 15258
rect 8558 15206 8568 15258
rect 8592 15206 8622 15258
rect 8622 15206 8648 15258
rect 8352 15204 8408 15206
rect 8432 15204 8488 15206
rect 8512 15204 8568 15206
rect 8592 15204 8648 15206
rect 8352 14170 8408 14172
rect 8432 14170 8488 14172
rect 8512 14170 8568 14172
rect 8592 14170 8648 14172
rect 8352 14118 8378 14170
rect 8378 14118 8408 14170
rect 8432 14118 8442 14170
rect 8442 14118 8488 14170
rect 8512 14118 8558 14170
rect 8558 14118 8568 14170
rect 8592 14118 8622 14170
rect 8622 14118 8648 14170
rect 8352 14116 8408 14118
rect 8432 14116 8488 14118
rect 8512 14116 8568 14118
rect 8592 14116 8648 14118
rect 8352 13082 8408 13084
rect 8432 13082 8488 13084
rect 8512 13082 8568 13084
rect 8592 13082 8648 13084
rect 8352 13030 8378 13082
rect 8378 13030 8408 13082
rect 8432 13030 8442 13082
rect 8442 13030 8488 13082
rect 8512 13030 8558 13082
rect 8558 13030 8568 13082
rect 8592 13030 8622 13082
rect 8622 13030 8648 13082
rect 8352 13028 8408 13030
rect 8432 13028 8488 13030
rect 8512 13028 8568 13030
rect 8592 13028 8648 13030
rect 8352 11994 8408 11996
rect 8432 11994 8488 11996
rect 8512 11994 8568 11996
rect 8592 11994 8648 11996
rect 8352 11942 8378 11994
rect 8378 11942 8408 11994
rect 8432 11942 8442 11994
rect 8442 11942 8488 11994
rect 8512 11942 8558 11994
rect 8558 11942 8568 11994
rect 8592 11942 8622 11994
rect 8622 11942 8648 11994
rect 8352 11940 8408 11942
rect 8432 11940 8488 11942
rect 8512 11940 8568 11942
rect 8592 11940 8648 11942
rect 8352 10906 8408 10908
rect 8432 10906 8488 10908
rect 8512 10906 8568 10908
rect 8592 10906 8648 10908
rect 8352 10854 8378 10906
rect 8378 10854 8408 10906
rect 8432 10854 8442 10906
rect 8442 10854 8488 10906
rect 8512 10854 8558 10906
rect 8558 10854 8568 10906
rect 8592 10854 8622 10906
rect 8622 10854 8648 10906
rect 8352 10852 8408 10854
rect 8432 10852 8488 10854
rect 8512 10852 8568 10854
rect 8592 10852 8648 10854
rect 8352 9818 8408 9820
rect 8432 9818 8488 9820
rect 8512 9818 8568 9820
rect 8592 9818 8648 9820
rect 8352 9766 8378 9818
rect 8378 9766 8408 9818
rect 8432 9766 8442 9818
rect 8442 9766 8488 9818
rect 8512 9766 8558 9818
rect 8558 9766 8568 9818
rect 8592 9766 8622 9818
rect 8622 9766 8648 9818
rect 8352 9764 8408 9766
rect 8432 9764 8488 9766
rect 8512 9764 8568 9766
rect 8592 9764 8648 9766
rect 8352 8730 8408 8732
rect 8432 8730 8488 8732
rect 8512 8730 8568 8732
rect 8592 8730 8648 8732
rect 8352 8678 8378 8730
rect 8378 8678 8408 8730
rect 8432 8678 8442 8730
rect 8442 8678 8488 8730
rect 8512 8678 8558 8730
rect 8558 8678 8568 8730
rect 8592 8678 8622 8730
rect 8622 8678 8648 8730
rect 8352 8676 8408 8678
rect 8432 8676 8488 8678
rect 8512 8676 8568 8678
rect 8592 8676 8648 8678
rect 8352 7642 8408 7644
rect 8432 7642 8488 7644
rect 8512 7642 8568 7644
rect 8592 7642 8648 7644
rect 8352 7590 8378 7642
rect 8378 7590 8408 7642
rect 8432 7590 8442 7642
rect 8442 7590 8488 7642
rect 8512 7590 8558 7642
rect 8558 7590 8568 7642
rect 8592 7590 8622 7642
rect 8622 7590 8648 7642
rect 8352 7588 8408 7590
rect 8432 7588 8488 7590
rect 8512 7588 8568 7590
rect 8592 7588 8648 7590
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 10817 16890 10873 16892
rect 10897 16890 10953 16892
rect 10977 16890 11033 16892
rect 11057 16890 11113 16892
rect 10817 16838 10843 16890
rect 10843 16838 10873 16890
rect 10897 16838 10907 16890
rect 10907 16838 10953 16890
rect 10977 16838 11023 16890
rect 11023 16838 11033 16890
rect 11057 16838 11087 16890
rect 11087 16838 11113 16890
rect 10817 16836 10873 16838
rect 10897 16836 10953 16838
rect 10977 16836 11033 16838
rect 11057 16836 11113 16838
rect 10817 15802 10873 15804
rect 10897 15802 10953 15804
rect 10977 15802 11033 15804
rect 11057 15802 11113 15804
rect 10817 15750 10843 15802
rect 10843 15750 10873 15802
rect 10897 15750 10907 15802
rect 10907 15750 10953 15802
rect 10977 15750 11023 15802
rect 11023 15750 11033 15802
rect 11057 15750 11087 15802
rect 11087 15750 11113 15802
rect 10817 15748 10873 15750
rect 10897 15748 10953 15750
rect 10977 15748 11033 15750
rect 11057 15748 11113 15750
rect 10817 14714 10873 14716
rect 10897 14714 10953 14716
rect 10977 14714 11033 14716
rect 11057 14714 11113 14716
rect 10817 14662 10843 14714
rect 10843 14662 10873 14714
rect 10897 14662 10907 14714
rect 10907 14662 10953 14714
rect 10977 14662 11023 14714
rect 11023 14662 11033 14714
rect 11057 14662 11087 14714
rect 11087 14662 11113 14714
rect 10817 14660 10873 14662
rect 10897 14660 10953 14662
rect 10977 14660 11033 14662
rect 11057 14660 11113 14662
rect 10817 13626 10873 13628
rect 10897 13626 10953 13628
rect 10977 13626 11033 13628
rect 11057 13626 11113 13628
rect 10817 13574 10843 13626
rect 10843 13574 10873 13626
rect 10897 13574 10907 13626
rect 10907 13574 10953 13626
rect 10977 13574 11023 13626
rect 11023 13574 11033 13626
rect 11057 13574 11087 13626
rect 11087 13574 11113 13626
rect 10817 13572 10873 13574
rect 10897 13572 10953 13574
rect 10977 13572 11033 13574
rect 11057 13572 11113 13574
rect 10817 12538 10873 12540
rect 10897 12538 10953 12540
rect 10977 12538 11033 12540
rect 11057 12538 11113 12540
rect 10817 12486 10843 12538
rect 10843 12486 10873 12538
rect 10897 12486 10907 12538
rect 10907 12486 10953 12538
rect 10977 12486 11023 12538
rect 11023 12486 11033 12538
rect 11057 12486 11087 12538
rect 11087 12486 11113 12538
rect 10817 12484 10873 12486
rect 10897 12484 10953 12486
rect 10977 12484 11033 12486
rect 11057 12484 11113 12486
rect 10414 9424 10470 9480
rect 10817 11450 10873 11452
rect 10897 11450 10953 11452
rect 10977 11450 11033 11452
rect 11057 11450 11113 11452
rect 10817 11398 10843 11450
rect 10843 11398 10873 11450
rect 10897 11398 10907 11450
rect 10907 11398 10953 11450
rect 10977 11398 11023 11450
rect 11023 11398 11033 11450
rect 11057 11398 11087 11450
rect 11087 11398 11113 11450
rect 10817 11396 10873 11398
rect 10897 11396 10953 11398
rect 10977 11396 11033 11398
rect 11057 11396 11113 11398
rect 10817 10362 10873 10364
rect 10897 10362 10953 10364
rect 10977 10362 11033 10364
rect 11057 10362 11113 10364
rect 10817 10310 10843 10362
rect 10843 10310 10873 10362
rect 10897 10310 10907 10362
rect 10907 10310 10953 10362
rect 10977 10310 11023 10362
rect 11023 10310 11033 10362
rect 11057 10310 11087 10362
rect 11087 10310 11113 10362
rect 10817 10308 10873 10310
rect 10897 10308 10953 10310
rect 10977 10308 11033 10310
rect 11057 10308 11113 10310
rect 10817 9274 10873 9276
rect 10897 9274 10953 9276
rect 10977 9274 11033 9276
rect 11057 9274 11113 9276
rect 10817 9222 10843 9274
rect 10843 9222 10873 9274
rect 10897 9222 10907 9274
rect 10907 9222 10953 9274
rect 10977 9222 11023 9274
rect 11023 9222 11033 9274
rect 11057 9222 11087 9274
rect 11087 9222 11113 9274
rect 10817 9220 10873 9222
rect 10897 9220 10953 9222
rect 10977 9220 11033 9222
rect 11057 9220 11113 9222
rect 11794 9696 11850 9752
rect 10817 8186 10873 8188
rect 10897 8186 10953 8188
rect 10977 8186 11033 8188
rect 11057 8186 11113 8188
rect 10817 8134 10843 8186
rect 10843 8134 10873 8186
rect 10897 8134 10907 8186
rect 10907 8134 10953 8186
rect 10977 8134 11023 8186
rect 11023 8134 11033 8186
rect 11057 8134 11087 8186
rect 11087 8134 11113 8186
rect 10817 8132 10873 8134
rect 10897 8132 10953 8134
rect 10977 8132 11033 8134
rect 11057 8132 11113 8134
rect 10817 7098 10873 7100
rect 10897 7098 10953 7100
rect 10977 7098 11033 7100
rect 11057 7098 11113 7100
rect 10817 7046 10843 7098
rect 10843 7046 10873 7098
rect 10897 7046 10907 7098
rect 10907 7046 10953 7098
rect 10977 7046 11023 7098
rect 11023 7046 11033 7098
rect 11057 7046 11087 7098
rect 11087 7046 11113 7098
rect 10817 7044 10873 7046
rect 10897 7044 10953 7046
rect 10977 7044 11033 7046
rect 11057 7044 11113 7046
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 13726 17448 13782 17504
rect 13282 17434 13338 17436
rect 13362 17434 13418 17436
rect 13442 17434 13498 17436
rect 13522 17434 13578 17436
rect 13282 17382 13308 17434
rect 13308 17382 13338 17434
rect 13362 17382 13372 17434
rect 13372 17382 13418 17434
rect 13442 17382 13488 17434
rect 13488 17382 13498 17434
rect 13522 17382 13552 17434
rect 13552 17382 13578 17434
rect 13282 17380 13338 17382
rect 13362 17380 13418 17382
rect 13442 17380 13498 17382
rect 13522 17380 13578 17382
rect 13282 16346 13338 16348
rect 13362 16346 13418 16348
rect 13442 16346 13498 16348
rect 13522 16346 13578 16348
rect 13282 16294 13308 16346
rect 13308 16294 13338 16346
rect 13362 16294 13372 16346
rect 13372 16294 13418 16346
rect 13442 16294 13488 16346
rect 13488 16294 13498 16346
rect 13522 16294 13552 16346
rect 13552 16294 13578 16346
rect 13282 16292 13338 16294
rect 13362 16292 13418 16294
rect 13442 16292 13498 16294
rect 13522 16292 13578 16294
rect 13282 15258 13338 15260
rect 13362 15258 13418 15260
rect 13442 15258 13498 15260
rect 13522 15258 13578 15260
rect 13282 15206 13308 15258
rect 13308 15206 13338 15258
rect 13362 15206 13372 15258
rect 13372 15206 13418 15258
rect 13442 15206 13488 15258
rect 13488 15206 13498 15258
rect 13522 15206 13552 15258
rect 13552 15206 13578 15258
rect 13282 15204 13338 15206
rect 13362 15204 13418 15206
rect 13442 15204 13498 15206
rect 13522 15204 13578 15206
rect 13282 14170 13338 14172
rect 13362 14170 13418 14172
rect 13442 14170 13498 14172
rect 13522 14170 13578 14172
rect 13282 14118 13308 14170
rect 13308 14118 13338 14170
rect 13362 14118 13372 14170
rect 13372 14118 13418 14170
rect 13442 14118 13488 14170
rect 13488 14118 13498 14170
rect 13522 14118 13552 14170
rect 13552 14118 13578 14170
rect 13282 14116 13338 14118
rect 13362 14116 13418 14118
rect 13442 14116 13498 14118
rect 13522 14116 13578 14118
rect 13282 13082 13338 13084
rect 13362 13082 13418 13084
rect 13442 13082 13498 13084
rect 13522 13082 13578 13084
rect 13282 13030 13308 13082
rect 13308 13030 13338 13082
rect 13362 13030 13372 13082
rect 13372 13030 13418 13082
rect 13442 13030 13488 13082
rect 13488 13030 13498 13082
rect 13522 13030 13552 13082
rect 13552 13030 13578 13082
rect 13282 13028 13338 13030
rect 13362 13028 13418 13030
rect 13442 13028 13498 13030
rect 13522 13028 13578 13030
rect 13726 12416 13782 12472
rect 13282 11994 13338 11996
rect 13362 11994 13418 11996
rect 13442 11994 13498 11996
rect 13522 11994 13578 11996
rect 13282 11942 13308 11994
rect 13308 11942 13338 11994
rect 13362 11942 13372 11994
rect 13372 11942 13418 11994
rect 13442 11942 13488 11994
rect 13488 11942 13498 11994
rect 13522 11942 13552 11994
rect 13552 11942 13578 11994
rect 13282 11940 13338 11942
rect 13362 11940 13418 11942
rect 13442 11940 13498 11942
rect 13522 11940 13578 11942
rect 13282 10906 13338 10908
rect 13362 10906 13418 10908
rect 13442 10906 13498 10908
rect 13522 10906 13578 10908
rect 13282 10854 13308 10906
rect 13308 10854 13338 10906
rect 13362 10854 13372 10906
rect 13372 10854 13418 10906
rect 13442 10854 13488 10906
rect 13488 10854 13498 10906
rect 13522 10854 13552 10906
rect 13552 10854 13578 10906
rect 13282 10852 13338 10854
rect 13362 10852 13418 10854
rect 13442 10852 13498 10854
rect 13522 10852 13578 10854
rect 13282 9818 13338 9820
rect 13362 9818 13418 9820
rect 13442 9818 13498 9820
rect 13522 9818 13578 9820
rect 13282 9766 13308 9818
rect 13308 9766 13338 9818
rect 13362 9766 13372 9818
rect 13372 9766 13418 9818
rect 13442 9766 13488 9818
rect 13488 9766 13498 9818
rect 13522 9766 13552 9818
rect 13552 9766 13578 9818
rect 13282 9764 13338 9766
rect 13362 9764 13418 9766
rect 13442 9764 13498 9766
rect 13522 9764 13578 9766
rect 13282 8730 13338 8732
rect 13362 8730 13418 8732
rect 13442 8730 13498 8732
rect 13522 8730 13578 8732
rect 13282 8678 13308 8730
rect 13308 8678 13338 8730
rect 13362 8678 13372 8730
rect 13372 8678 13418 8730
rect 13442 8678 13488 8730
rect 13488 8678 13498 8730
rect 13522 8678 13552 8730
rect 13552 8678 13578 8730
rect 13282 8676 13338 8678
rect 13362 8676 13418 8678
rect 13442 8676 13498 8678
rect 13522 8676 13578 8678
rect 13282 7642 13338 7644
rect 13362 7642 13418 7644
rect 13442 7642 13498 7644
rect 13522 7642 13578 7644
rect 13282 7590 13308 7642
rect 13308 7590 13338 7642
rect 13362 7590 13372 7642
rect 13372 7590 13418 7642
rect 13442 7590 13488 7642
rect 13488 7590 13498 7642
rect 13522 7590 13552 7642
rect 13552 7590 13578 7642
rect 13282 7588 13338 7590
rect 13362 7588 13418 7590
rect 13442 7588 13498 7590
rect 13522 7588 13578 7590
rect 12530 7384 12586 7440
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 13726 2488 13782 2544
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
<< metal3 >>
rect 0 18322 480 18352
rect 3785 18322 3851 18325
rect 0 18320 3851 18322
rect 0 18264 3790 18320
rect 3846 18264 3851 18320
rect 0 18262 3851 18264
rect 0 18232 480 18262
rect 3785 18259 3851 18262
rect 13721 17506 13787 17509
rect 16520 17506 17000 17536
rect 13721 17504 17000 17506
rect 13721 17448 13726 17504
rect 13782 17448 17000 17504
rect 13721 17446 17000 17448
rect 13721 17443 13787 17446
rect 3409 17440 3729 17441
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 17375 3729 17376
rect 8340 17440 8660 17441
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 17375 8660 17376
rect 13270 17440 13590 17441
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 16520 17416 17000 17446
rect 13270 17375 13590 17376
rect 5874 16896 6194 16897
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6194 16896
rect 5874 16831 6194 16832
rect 10805 16896 11125 16897
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 16831 11125 16832
rect 3409 16352 3729 16353
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 16287 3729 16288
rect 8340 16352 8660 16353
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 16287 8660 16288
rect 13270 16352 13590 16353
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 16287 13590 16288
rect 5874 15808 6194 15809
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6194 15808
rect 5874 15743 6194 15744
rect 10805 15808 11125 15809
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 15743 11125 15744
rect 3409 15264 3729 15265
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 15199 3729 15200
rect 8340 15264 8660 15265
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 15199 8660 15200
rect 13270 15264 13590 15265
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 15199 13590 15200
rect 0 15058 480 15088
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14968 480 14998
rect 2773 14995 2839 14998
rect 5874 14720 6194 14721
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6194 14720
rect 5874 14655 6194 14656
rect 10805 14720 11125 14721
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 14655 11125 14656
rect 3409 14176 3729 14177
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 14111 3729 14112
rect 8340 14176 8660 14177
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 14111 8660 14112
rect 13270 14176 13590 14177
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 14111 13590 14112
rect 5874 13632 6194 13633
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6194 13632
rect 5874 13567 6194 13568
rect 10805 13632 11125 13633
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 13567 11125 13568
rect 3409 13088 3729 13089
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 13023 3729 13024
rect 8340 13088 8660 13089
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 13023 8660 13024
rect 13270 13088 13590 13089
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 13023 13590 13024
rect 5874 12544 6194 12545
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6194 12544
rect 5874 12479 6194 12480
rect 10805 12544 11125 12545
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 12479 11125 12480
rect 13721 12474 13787 12477
rect 16520 12474 17000 12504
rect 13721 12472 17000 12474
rect 13721 12416 13726 12472
rect 13782 12416 17000 12472
rect 13721 12414 17000 12416
rect 13721 12411 13787 12414
rect 16520 12384 17000 12414
rect 3409 12000 3729 12001
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 11935 3729 11936
rect 8340 12000 8660 12001
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 11935 8660 11936
rect 13270 12000 13590 12001
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 11935 13590 11936
rect 0 11658 480 11688
rect 4061 11658 4127 11661
rect 0 11656 4127 11658
rect 0 11600 4066 11656
rect 4122 11600 4127 11656
rect 0 11598 4127 11600
rect 0 11568 480 11598
rect 4061 11595 4127 11598
rect 5874 11456 6194 11457
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6194 11456
rect 5874 11391 6194 11392
rect 10805 11456 11125 11457
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 11391 11125 11392
rect 3409 10912 3729 10913
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 10847 3729 10848
rect 8340 10912 8660 10913
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 10847 8660 10848
rect 13270 10912 13590 10913
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 10847 13590 10848
rect 5874 10368 6194 10369
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6194 10368
rect 5874 10303 6194 10304
rect 10805 10368 11125 10369
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 10303 11125 10304
rect 3409 9824 3729 9825
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 9759 3729 9760
rect 8340 9824 8660 9825
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 9759 8660 9760
rect 13270 9824 13590 9825
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 9759 13590 9760
rect 11789 9754 11855 9757
rect 11286 9752 11855 9754
rect 11286 9696 11794 9752
rect 11850 9696 11855 9752
rect 11286 9694 11855 9696
rect 10409 9482 10475 9485
rect 11286 9482 11346 9694
rect 11789 9691 11855 9694
rect 10409 9480 11346 9482
rect 10409 9424 10414 9480
rect 10470 9424 11346 9480
rect 10409 9422 11346 9424
rect 10409 9419 10475 9422
rect 5874 9280 6194 9281
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6194 9280
rect 5874 9215 6194 9216
rect 10805 9280 11125 9281
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 9215 11125 9216
rect 3409 8736 3729 8737
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 8671 3729 8672
rect 8340 8736 8660 8737
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 8671 8660 8672
rect 13270 8736 13590 8737
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 8671 13590 8672
rect 0 8394 480 8424
rect 1577 8394 1643 8397
rect 0 8392 1643 8394
rect 0 8336 1582 8392
rect 1638 8336 1643 8392
rect 0 8334 1643 8336
rect 0 8304 480 8334
rect 1577 8331 1643 8334
rect 5874 8192 6194 8193
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6194 8192
rect 5874 8127 6194 8128
rect 10805 8192 11125 8193
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 8127 11125 8128
rect 3409 7648 3729 7649
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 7583 3729 7584
rect 8340 7648 8660 7649
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 7583 8660 7584
rect 13270 7648 13590 7649
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 7583 13590 7584
rect 12525 7442 12591 7445
rect 16520 7442 17000 7472
rect 12525 7440 17000 7442
rect 12525 7384 12530 7440
rect 12586 7384 17000 7440
rect 12525 7382 17000 7384
rect 12525 7379 12591 7382
rect 16520 7352 17000 7382
rect 5874 7104 6194 7105
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6194 7104
rect 5874 7039 6194 7040
rect 10805 7104 11125 7105
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 7039 11125 7040
rect 3409 6560 3729 6561
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 3409 5472 3729 5473
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 0 4994 480 5024
rect 3049 4994 3115 4997
rect 0 4992 3115 4994
rect 0 4936 3054 4992
rect 3110 4936 3115 4992
rect 0 4934 3115 4936
rect 0 4904 480 4934
rect 3049 4931 3115 4934
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 3409 4384 3729 4385
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 4319 13590 4320
rect 5874 3840 6194 3841
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 3231 13590 3232
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 13721 2546 13787 2549
rect 16520 2546 17000 2576
rect 13721 2544 17000 2546
rect 13721 2488 13726 2544
rect 13782 2488 17000 2544
rect 13721 2486 17000 2488
rect 13721 2483 13787 2486
rect 16520 2456 17000 2486
rect 3409 2208 3729 2209
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
rect 0 1730 480 1760
rect 1117 1730 1183 1733
rect 0 1728 1183 1730
rect 0 1672 1122 1728
rect 1178 1672 1183 1728
rect 0 1670 1183 1672
rect 0 1640 480 1670
rect 1117 1667 1183 1670
<< via3 >>
rect 3417 17436 3481 17440
rect 3417 17380 3421 17436
rect 3421 17380 3477 17436
rect 3477 17380 3481 17436
rect 3417 17376 3481 17380
rect 3497 17436 3561 17440
rect 3497 17380 3501 17436
rect 3501 17380 3557 17436
rect 3557 17380 3561 17436
rect 3497 17376 3561 17380
rect 3577 17436 3641 17440
rect 3577 17380 3581 17436
rect 3581 17380 3637 17436
rect 3637 17380 3641 17436
rect 3577 17376 3641 17380
rect 3657 17436 3721 17440
rect 3657 17380 3661 17436
rect 3661 17380 3717 17436
rect 3717 17380 3721 17436
rect 3657 17376 3721 17380
rect 8348 17436 8412 17440
rect 8348 17380 8352 17436
rect 8352 17380 8408 17436
rect 8408 17380 8412 17436
rect 8348 17376 8412 17380
rect 8428 17436 8492 17440
rect 8428 17380 8432 17436
rect 8432 17380 8488 17436
rect 8488 17380 8492 17436
rect 8428 17376 8492 17380
rect 8508 17436 8572 17440
rect 8508 17380 8512 17436
rect 8512 17380 8568 17436
rect 8568 17380 8572 17436
rect 8508 17376 8572 17380
rect 8588 17436 8652 17440
rect 8588 17380 8592 17436
rect 8592 17380 8648 17436
rect 8648 17380 8652 17436
rect 8588 17376 8652 17380
rect 13278 17436 13342 17440
rect 13278 17380 13282 17436
rect 13282 17380 13338 17436
rect 13338 17380 13342 17436
rect 13278 17376 13342 17380
rect 13358 17436 13422 17440
rect 13358 17380 13362 17436
rect 13362 17380 13418 17436
rect 13418 17380 13422 17436
rect 13358 17376 13422 17380
rect 13438 17436 13502 17440
rect 13438 17380 13442 17436
rect 13442 17380 13498 17436
rect 13498 17380 13502 17436
rect 13438 17376 13502 17380
rect 13518 17436 13582 17440
rect 13518 17380 13522 17436
rect 13522 17380 13578 17436
rect 13578 17380 13582 17436
rect 13518 17376 13582 17380
rect 5882 16892 5946 16896
rect 5882 16836 5886 16892
rect 5886 16836 5942 16892
rect 5942 16836 5946 16892
rect 5882 16832 5946 16836
rect 5962 16892 6026 16896
rect 5962 16836 5966 16892
rect 5966 16836 6022 16892
rect 6022 16836 6026 16892
rect 5962 16832 6026 16836
rect 6042 16892 6106 16896
rect 6042 16836 6046 16892
rect 6046 16836 6102 16892
rect 6102 16836 6106 16892
rect 6042 16832 6106 16836
rect 6122 16892 6186 16896
rect 6122 16836 6126 16892
rect 6126 16836 6182 16892
rect 6182 16836 6186 16892
rect 6122 16832 6186 16836
rect 10813 16892 10877 16896
rect 10813 16836 10817 16892
rect 10817 16836 10873 16892
rect 10873 16836 10877 16892
rect 10813 16832 10877 16836
rect 10893 16892 10957 16896
rect 10893 16836 10897 16892
rect 10897 16836 10953 16892
rect 10953 16836 10957 16892
rect 10893 16832 10957 16836
rect 10973 16892 11037 16896
rect 10973 16836 10977 16892
rect 10977 16836 11033 16892
rect 11033 16836 11037 16892
rect 10973 16832 11037 16836
rect 11053 16892 11117 16896
rect 11053 16836 11057 16892
rect 11057 16836 11113 16892
rect 11113 16836 11117 16892
rect 11053 16832 11117 16836
rect 3417 16348 3481 16352
rect 3417 16292 3421 16348
rect 3421 16292 3477 16348
rect 3477 16292 3481 16348
rect 3417 16288 3481 16292
rect 3497 16348 3561 16352
rect 3497 16292 3501 16348
rect 3501 16292 3557 16348
rect 3557 16292 3561 16348
rect 3497 16288 3561 16292
rect 3577 16348 3641 16352
rect 3577 16292 3581 16348
rect 3581 16292 3637 16348
rect 3637 16292 3641 16348
rect 3577 16288 3641 16292
rect 3657 16348 3721 16352
rect 3657 16292 3661 16348
rect 3661 16292 3717 16348
rect 3717 16292 3721 16348
rect 3657 16288 3721 16292
rect 8348 16348 8412 16352
rect 8348 16292 8352 16348
rect 8352 16292 8408 16348
rect 8408 16292 8412 16348
rect 8348 16288 8412 16292
rect 8428 16348 8492 16352
rect 8428 16292 8432 16348
rect 8432 16292 8488 16348
rect 8488 16292 8492 16348
rect 8428 16288 8492 16292
rect 8508 16348 8572 16352
rect 8508 16292 8512 16348
rect 8512 16292 8568 16348
rect 8568 16292 8572 16348
rect 8508 16288 8572 16292
rect 8588 16348 8652 16352
rect 8588 16292 8592 16348
rect 8592 16292 8648 16348
rect 8648 16292 8652 16348
rect 8588 16288 8652 16292
rect 13278 16348 13342 16352
rect 13278 16292 13282 16348
rect 13282 16292 13338 16348
rect 13338 16292 13342 16348
rect 13278 16288 13342 16292
rect 13358 16348 13422 16352
rect 13358 16292 13362 16348
rect 13362 16292 13418 16348
rect 13418 16292 13422 16348
rect 13358 16288 13422 16292
rect 13438 16348 13502 16352
rect 13438 16292 13442 16348
rect 13442 16292 13498 16348
rect 13498 16292 13502 16348
rect 13438 16288 13502 16292
rect 13518 16348 13582 16352
rect 13518 16292 13522 16348
rect 13522 16292 13578 16348
rect 13578 16292 13582 16348
rect 13518 16288 13582 16292
rect 5882 15804 5946 15808
rect 5882 15748 5886 15804
rect 5886 15748 5942 15804
rect 5942 15748 5946 15804
rect 5882 15744 5946 15748
rect 5962 15804 6026 15808
rect 5962 15748 5966 15804
rect 5966 15748 6022 15804
rect 6022 15748 6026 15804
rect 5962 15744 6026 15748
rect 6042 15804 6106 15808
rect 6042 15748 6046 15804
rect 6046 15748 6102 15804
rect 6102 15748 6106 15804
rect 6042 15744 6106 15748
rect 6122 15804 6186 15808
rect 6122 15748 6126 15804
rect 6126 15748 6182 15804
rect 6182 15748 6186 15804
rect 6122 15744 6186 15748
rect 10813 15804 10877 15808
rect 10813 15748 10817 15804
rect 10817 15748 10873 15804
rect 10873 15748 10877 15804
rect 10813 15744 10877 15748
rect 10893 15804 10957 15808
rect 10893 15748 10897 15804
rect 10897 15748 10953 15804
rect 10953 15748 10957 15804
rect 10893 15744 10957 15748
rect 10973 15804 11037 15808
rect 10973 15748 10977 15804
rect 10977 15748 11033 15804
rect 11033 15748 11037 15804
rect 10973 15744 11037 15748
rect 11053 15804 11117 15808
rect 11053 15748 11057 15804
rect 11057 15748 11113 15804
rect 11113 15748 11117 15804
rect 11053 15744 11117 15748
rect 3417 15260 3481 15264
rect 3417 15204 3421 15260
rect 3421 15204 3477 15260
rect 3477 15204 3481 15260
rect 3417 15200 3481 15204
rect 3497 15260 3561 15264
rect 3497 15204 3501 15260
rect 3501 15204 3557 15260
rect 3557 15204 3561 15260
rect 3497 15200 3561 15204
rect 3577 15260 3641 15264
rect 3577 15204 3581 15260
rect 3581 15204 3637 15260
rect 3637 15204 3641 15260
rect 3577 15200 3641 15204
rect 3657 15260 3721 15264
rect 3657 15204 3661 15260
rect 3661 15204 3717 15260
rect 3717 15204 3721 15260
rect 3657 15200 3721 15204
rect 8348 15260 8412 15264
rect 8348 15204 8352 15260
rect 8352 15204 8408 15260
rect 8408 15204 8412 15260
rect 8348 15200 8412 15204
rect 8428 15260 8492 15264
rect 8428 15204 8432 15260
rect 8432 15204 8488 15260
rect 8488 15204 8492 15260
rect 8428 15200 8492 15204
rect 8508 15260 8572 15264
rect 8508 15204 8512 15260
rect 8512 15204 8568 15260
rect 8568 15204 8572 15260
rect 8508 15200 8572 15204
rect 8588 15260 8652 15264
rect 8588 15204 8592 15260
rect 8592 15204 8648 15260
rect 8648 15204 8652 15260
rect 8588 15200 8652 15204
rect 13278 15260 13342 15264
rect 13278 15204 13282 15260
rect 13282 15204 13338 15260
rect 13338 15204 13342 15260
rect 13278 15200 13342 15204
rect 13358 15260 13422 15264
rect 13358 15204 13362 15260
rect 13362 15204 13418 15260
rect 13418 15204 13422 15260
rect 13358 15200 13422 15204
rect 13438 15260 13502 15264
rect 13438 15204 13442 15260
rect 13442 15204 13498 15260
rect 13498 15204 13502 15260
rect 13438 15200 13502 15204
rect 13518 15260 13582 15264
rect 13518 15204 13522 15260
rect 13522 15204 13578 15260
rect 13578 15204 13582 15260
rect 13518 15200 13582 15204
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 6122 14716 6186 14720
rect 6122 14660 6126 14716
rect 6126 14660 6182 14716
rect 6182 14660 6186 14716
rect 6122 14656 6186 14660
rect 10813 14716 10877 14720
rect 10813 14660 10817 14716
rect 10817 14660 10873 14716
rect 10873 14660 10877 14716
rect 10813 14656 10877 14660
rect 10893 14716 10957 14720
rect 10893 14660 10897 14716
rect 10897 14660 10953 14716
rect 10953 14660 10957 14716
rect 10893 14656 10957 14660
rect 10973 14716 11037 14720
rect 10973 14660 10977 14716
rect 10977 14660 11033 14716
rect 11033 14660 11037 14716
rect 10973 14656 11037 14660
rect 11053 14716 11117 14720
rect 11053 14660 11057 14716
rect 11057 14660 11113 14716
rect 11113 14660 11117 14716
rect 11053 14656 11117 14660
rect 3417 14172 3481 14176
rect 3417 14116 3421 14172
rect 3421 14116 3477 14172
rect 3477 14116 3481 14172
rect 3417 14112 3481 14116
rect 3497 14172 3561 14176
rect 3497 14116 3501 14172
rect 3501 14116 3557 14172
rect 3557 14116 3561 14172
rect 3497 14112 3561 14116
rect 3577 14172 3641 14176
rect 3577 14116 3581 14172
rect 3581 14116 3637 14172
rect 3637 14116 3641 14172
rect 3577 14112 3641 14116
rect 3657 14172 3721 14176
rect 3657 14116 3661 14172
rect 3661 14116 3717 14172
rect 3717 14116 3721 14172
rect 3657 14112 3721 14116
rect 8348 14172 8412 14176
rect 8348 14116 8352 14172
rect 8352 14116 8408 14172
rect 8408 14116 8412 14172
rect 8348 14112 8412 14116
rect 8428 14172 8492 14176
rect 8428 14116 8432 14172
rect 8432 14116 8488 14172
rect 8488 14116 8492 14172
rect 8428 14112 8492 14116
rect 8508 14172 8572 14176
rect 8508 14116 8512 14172
rect 8512 14116 8568 14172
rect 8568 14116 8572 14172
rect 8508 14112 8572 14116
rect 8588 14172 8652 14176
rect 8588 14116 8592 14172
rect 8592 14116 8648 14172
rect 8648 14116 8652 14172
rect 8588 14112 8652 14116
rect 13278 14172 13342 14176
rect 13278 14116 13282 14172
rect 13282 14116 13338 14172
rect 13338 14116 13342 14172
rect 13278 14112 13342 14116
rect 13358 14172 13422 14176
rect 13358 14116 13362 14172
rect 13362 14116 13418 14172
rect 13418 14116 13422 14172
rect 13358 14112 13422 14116
rect 13438 14172 13502 14176
rect 13438 14116 13442 14172
rect 13442 14116 13498 14172
rect 13498 14116 13502 14172
rect 13438 14112 13502 14116
rect 13518 14172 13582 14176
rect 13518 14116 13522 14172
rect 13522 14116 13578 14172
rect 13578 14116 13582 14172
rect 13518 14112 13582 14116
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 6122 13628 6186 13632
rect 6122 13572 6126 13628
rect 6126 13572 6182 13628
rect 6182 13572 6186 13628
rect 6122 13568 6186 13572
rect 10813 13628 10877 13632
rect 10813 13572 10817 13628
rect 10817 13572 10873 13628
rect 10873 13572 10877 13628
rect 10813 13568 10877 13572
rect 10893 13628 10957 13632
rect 10893 13572 10897 13628
rect 10897 13572 10953 13628
rect 10953 13572 10957 13628
rect 10893 13568 10957 13572
rect 10973 13628 11037 13632
rect 10973 13572 10977 13628
rect 10977 13572 11033 13628
rect 11033 13572 11037 13628
rect 10973 13568 11037 13572
rect 11053 13628 11117 13632
rect 11053 13572 11057 13628
rect 11057 13572 11113 13628
rect 11113 13572 11117 13628
rect 11053 13568 11117 13572
rect 3417 13084 3481 13088
rect 3417 13028 3421 13084
rect 3421 13028 3477 13084
rect 3477 13028 3481 13084
rect 3417 13024 3481 13028
rect 3497 13084 3561 13088
rect 3497 13028 3501 13084
rect 3501 13028 3557 13084
rect 3557 13028 3561 13084
rect 3497 13024 3561 13028
rect 3577 13084 3641 13088
rect 3577 13028 3581 13084
rect 3581 13028 3637 13084
rect 3637 13028 3641 13084
rect 3577 13024 3641 13028
rect 3657 13084 3721 13088
rect 3657 13028 3661 13084
rect 3661 13028 3717 13084
rect 3717 13028 3721 13084
rect 3657 13024 3721 13028
rect 8348 13084 8412 13088
rect 8348 13028 8352 13084
rect 8352 13028 8408 13084
rect 8408 13028 8412 13084
rect 8348 13024 8412 13028
rect 8428 13084 8492 13088
rect 8428 13028 8432 13084
rect 8432 13028 8488 13084
rect 8488 13028 8492 13084
rect 8428 13024 8492 13028
rect 8508 13084 8572 13088
rect 8508 13028 8512 13084
rect 8512 13028 8568 13084
rect 8568 13028 8572 13084
rect 8508 13024 8572 13028
rect 8588 13084 8652 13088
rect 8588 13028 8592 13084
rect 8592 13028 8648 13084
rect 8648 13028 8652 13084
rect 8588 13024 8652 13028
rect 13278 13084 13342 13088
rect 13278 13028 13282 13084
rect 13282 13028 13338 13084
rect 13338 13028 13342 13084
rect 13278 13024 13342 13028
rect 13358 13084 13422 13088
rect 13358 13028 13362 13084
rect 13362 13028 13418 13084
rect 13418 13028 13422 13084
rect 13358 13024 13422 13028
rect 13438 13084 13502 13088
rect 13438 13028 13442 13084
rect 13442 13028 13498 13084
rect 13498 13028 13502 13084
rect 13438 13024 13502 13028
rect 13518 13084 13582 13088
rect 13518 13028 13522 13084
rect 13522 13028 13578 13084
rect 13578 13028 13582 13084
rect 13518 13024 13582 13028
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 6122 12540 6186 12544
rect 6122 12484 6126 12540
rect 6126 12484 6182 12540
rect 6182 12484 6186 12540
rect 6122 12480 6186 12484
rect 10813 12540 10877 12544
rect 10813 12484 10817 12540
rect 10817 12484 10873 12540
rect 10873 12484 10877 12540
rect 10813 12480 10877 12484
rect 10893 12540 10957 12544
rect 10893 12484 10897 12540
rect 10897 12484 10953 12540
rect 10953 12484 10957 12540
rect 10893 12480 10957 12484
rect 10973 12540 11037 12544
rect 10973 12484 10977 12540
rect 10977 12484 11033 12540
rect 11033 12484 11037 12540
rect 10973 12480 11037 12484
rect 11053 12540 11117 12544
rect 11053 12484 11057 12540
rect 11057 12484 11113 12540
rect 11113 12484 11117 12540
rect 11053 12480 11117 12484
rect 3417 11996 3481 12000
rect 3417 11940 3421 11996
rect 3421 11940 3477 11996
rect 3477 11940 3481 11996
rect 3417 11936 3481 11940
rect 3497 11996 3561 12000
rect 3497 11940 3501 11996
rect 3501 11940 3557 11996
rect 3557 11940 3561 11996
rect 3497 11936 3561 11940
rect 3577 11996 3641 12000
rect 3577 11940 3581 11996
rect 3581 11940 3637 11996
rect 3637 11940 3641 11996
rect 3577 11936 3641 11940
rect 3657 11996 3721 12000
rect 3657 11940 3661 11996
rect 3661 11940 3717 11996
rect 3717 11940 3721 11996
rect 3657 11936 3721 11940
rect 8348 11996 8412 12000
rect 8348 11940 8352 11996
rect 8352 11940 8408 11996
rect 8408 11940 8412 11996
rect 8348 11936 8412 11940
rect 8428 11996 8492 12000
rect 8428 11940 8432 11996
rect 8432 11940 8488 11996
rect 8488 11940 8492 11996
rect 8428 11936 8492 11940
rect 8508 11996 8572 12000
rect 8508 11940 8512 11996
rect 8512 11940 8568 11996
rect 8568 11940 8572 11996
rect 8508 11936 8572 11940
rect 8588 11996 8652 12000
rect 8588 11940 8592 11996
rect 8592 11940 8648 11996
rect 8648 11940 8652 11996
rect 8588 11936 8652 11940
rect 13278 11996 13342 12000
rect 13278 11940 13282 11996
rect 13282 11940 13338 11996
rect 13338 11940 13342 11996
rect 13278 11936 13342 11940
rect 13358 11996 13422 12000
rect 13358 11940 13362 11996
rect 13362 11940 13418 11996
rect 13418 11940 13422 11996
rect 13358 11936 13422 11940
rect 13438 11996 13502 12000
rect 13438 11940 13442 11996
rect 13442 11940 13498 11996
rect 13498 11940 13502 11996
rect 13438 11936 13502 11940
rect 13518 11996 13582 12000
rect 13518 11940 13522 11996
rect 13522 11940 13578 11996
rect 13578 11940 13582 11996
rect 13518 11936 13582 11940
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 6122 11452 6186 11456
rect 6122 11396 6126 11452
rect 6126 11396 6182 11452
rect 6182 11396 6186 11452
rect 6122 11392 6186 11396
rect 10813 11452 10877 11456
rect 10813 11396 10817 11452
rect 10817 11396 10873 11452
rect 10873 11396 10877 11452
rect 10813 11392 10877 11396
rect 10893 11452 10957 11456
rect 10893 11396 10897 11452
rect 10897 11396 10953 11452
rect 10953 11396 10957 11452
rect 10893 11392 10957 11396
rect 10973 11452 11037 11456
rect 10973 11396 10977 11452
rect 10977 11396 11033 11452
rect 11033 11396 11037 11452
rect 10973 11392 11037 11396
rect 11053 11452 11117 11456
rect 11053 11396 11057 11452
rect 11057 11396 11113 11452
rect 11113 11396 11117 11452
rect 11053 11392 11117 11396
rect 3417 10908 3481 10912
rect 3417 10852 3421 10908
rect 3421 10852 3477 10908
rect 3477 10852 3481 10908
rect 3417 10848 3481 10852
rect 3497 10908 3561 10912
rect 3497 10852 3501 10908
rect 3501 10852 3557 10908
rect 3557 10852 3561 10908
rect 3497 10848 3561 10852
rect 3577 10908 3641 10912
rect 3577 10852 3581 10908
rect 3581 10852 3637 10908
rect 3637 10852 3641 10908
rect 3577 10848 3641 10852
rect 3657 10908 3721 10912
rect 3657 10852 3661 10908
rect 3661 10852 3717 10908
rect 3717 10852 3721 10908
rect 3657 10848 3721 10852
rect 8348 10908 8412 10912
rect 8348 10852 8352 10908
rect 8352 10852 8408 10908
rect 8408 10852 8412 10908
rect 8348 10848 8412 10852
rect 8428 10908 8492 10912
rect 8428 10852 8432 10908
rect 8432 10852 8488 10908
rect 8488 10852 8492 10908
rect 8428 10848 8492 10852
rect 8508 10908 8572 10912
rect 8508 10852 8512 10908
rect 8512 10852 8568 10908
rect 8568 10852 8572 10908
rect 8508 10848 8572 10852
rect 8588 10908 8652 10912
rect 8588 10852 8592 10908
rect 8592 10852 8648 10908
rect 8648 10852 8652 10908
rect 8588 10848 8652 10852
rect 13278 10908 13342 10912
rect 13278 10852 13282 10908
rect 13282 10852 13338 10908
rect 13338 10852 13342 10908
rect 13278 10848 13342 10852
rect 13358 10908 13422 10912
rect 13358 10852 13362 10908
rect 13362 10852 13418 10908
rect 13418 10852 13422 10908
rect 13358 10848 13422 10852
rect 13438 10908 13502 10912
rect 13438 10852 13442 10908
rect 13442 10852 13498 10908
rect 13498 10852 13502 10908
rect 13438 10848 13502 10852
rect 13518 10908 13582 10912
rect 13518 10852 13522 10908
rect 13522 10852 13578 10908
rect 13578 10852 13582 10908
rect 13518 10848 13582 10852
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 6122 10364 6186 10368
rect 6122 10308 6126 10364
rect 6126 10308 6182 10364
rect 6182 10308 6186 10364
rect 6122 10304 6186 10308
rect 10813 10364 10877 10368
rect 10813 10308 10817 10364
rect 10817 10308 10873 10364
rect 10873 10308 10877 10364
rect 10813 10304 10877 10308
rect 10893 10364 10957 10368
rect 10893 10308 10897 10364
rect 10897 10308 10953 10364
rect 10953 10308 10957 10364
rect 10893 10304 10957 10308
rect 10973 10364 11037 10368
rect 10973 10308 10977 10364
rect 10977 10308 11033 10364
rect 11033 10308 11037 10364
rect 10973 10304 11037 10308
rect 11053 10364 11117 10368
rect 11053 10308 11057 10364
rect 11057 10308 11113 10364
rect 11113 10308 11117 10364
rect 11053 10304 11117 10308
rect 3417 9820 3481 9824
rect 3417 9764 3421 9820
rect 3421 9764 3477 9820
rect 3477 9764 3481 9820
rect 3417 9760 3481 9764
rect 3497 9820 3561 9824
rect 3497 9764 3501 9820
rect 3501 9764 3557 9820
rect 3557 9764 3561 9820
rect 3497 9760 3561 9764
rect 3577 9820 3641 9824
rect 3577 9764 3581 9820
rect 3581 9764 3637 9820
rect 3637 9764 3641 9820
rect 3577 9760 3641 9764
rect 3657 9820 3721 9824
rect 3657 9764 3661 9820
rect 3661 9764 3717 9820
rect 3717 9764 3721 9820
rect 3657 9760 3721 9764
rect 8348 9820 8412 9824
rect 8348 9764 8352 9820
rect 8352 9764 8408 9820
rect 8408 9764 8412 9820
rect 8348 9760 8412 9764
rect 8428 9820 8492 9824
rect 8428 9764 8432 9820
rect 8432 9764 8488 9820
rect 8488 9764 8492 9820
rect 8428 9760 8492 9764
rect 8508 9820 8572 9824
rect 8508 9764 8512 9820
rect 8512 9764 8568 9820
rect 8568 9764 8572 9820
rect 8508 9760 8572 9764
rect 8588 9820 8652 9824
rect 8588 9764 8592 9820
rect 8592 9764 8648 9820
rect 8648 9764 8652 9820
rect 8588 9760 8652 9764
rect 13278 9820 13342 9824
rect 13278 9764 13282 9820
rect 13282 9764 13338 9820
rect 13338 9764 13342 9820
rect 13278 9760 13342 9764
rect 13358 9820 13422 9824
rect 13358 9764 13362 9820
rect 13362 9764 13418 9820
rect 13418 9764 13422 9820
rect 13358 9760 13422 9764
rect 13438 9820 13502 9824
rect 13438 9764 13442 9820
rect 13442 9764 13498 9820
rect 13498 9764 13502 9820
rect 13438 9760 13502 9764
rect 13518 9820 13582 9824
rect 13518 9764 13522 9820
rect 13522 9764 13578 9820
rect 13578 9764 13582 9820
rect 13518 9760 13582 9764
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 6122 9276 6186 9280
rect 6122 9220 6126 9276
rect 6126 9220 6182 9276
rect 6182 9220 6186 9276
rect 6122 9216 6186 9220
rect 10813 9276 10877 9280
rect 10813 9220 10817 9276
rect 10817 9220 10873 9276
rect 10873 9220 10877 9276
rect 10813 9216 10877 9220
rect 10893 9276 10957 9280
rect 10893 9220 10897 9276
rect 10897 9220 10953 9276
rect 10953 9220 10957 9276
rect 10893 9216 10957 9220
rect 10973 9276 11037 9280
rect 10973 9220 10977 9276
rect 10977 9220 11033 9276
rect 11033 9220 11037 9276
rect 10973 9216 11037 9220
rect 11053 9276 11117 9280
rect 11053 9220 11057 9276
rect 11057 9220 11113 9276
rect 11113 9220 11117 9276
rect 11053 9216 11117 9220
rect 3417 8732 3481 8736
rect 3417 8676 3421 8732
rect 3421 8676 3477 8732
rect 3477 8676 3481 8732
rect 3417 8672 3481 8676
rect 3497 8732 3561 8736
rect 3497 8676 3501 8732
rect 3501 8676 3557 8732
rect 3557 8676 3561 8732
rect 3497 8672 3561 8676
rect 3577 8732 3641 8736
rect 3577 8676 3581 8732
rect 3581 8676 3637 8732
rect 3637 8676 3641 8732
rect 3577 8672 3641 8676
rect 3657 8732 3721 8736
rect 3657 8676 3661 8732
rect 3661 8676 3717 8732
rect 3717 8676 3721 8732
rect 3657 8672 3721 8676
rect 8348 8732 8412 8736
rect 8348 8676 8352 8732
rect 8352 8676 8408 8732
rect 8408 8676 8412 8732
rect 8348 8672 8412 8676
rect 8428 8732 8492 8736
rect 8428 8676 8432 8732
rect 8432 8676 8488 8732
rect 8488 8676 8492 8732
rect 8428 8672 8492 8676
rect 8508 8732 8572 8736
rect 8508 8676 8512 8732
rect 8512 8676 8568 8732
rect 8568 8676 8572 8732
rect 8508 8672 8572 8676
rect 8588 8732 8652 8736
rect 8588 8676 8592 8732
rect 8592 8676 8648 8732
rect 8648 8676 8652 8732
rect 8588 8672 8652 8676
rect 13278 8732 13342 8736
rect 13278 8676 13282 8732
rect 13282 8676 13338 8732
rect 13338 8676 13342 8732
rect 13278 8672 13342 8676
rect 13358 8732 13422 8736
rect 13358 8676 13362 8732
rect 13362 8676 13418 8732
rect 13418 8676 13422 8732
rect 13358 8672 13422 8676
rect 13438 8732 13502 8736
rect 13438 8676 13442 8732
rect 13442 8676 13498 8732
rect 13498 8676 13502 8732
rect 13438 8672 13502 8676
rect 13518 8732 13582 8736
rect 13518 8676 13522 8732
rect 13522 8676 13578 8732
rect 13578 8676 13582 8732
rect 13518 8672 13582 8676
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 6122 8188 6186 8192
rect 6122 8132 6126 8188
rect 6126 8132 6182 8188
rect 6182 8132 6186 8188
rect 6122 8128 6186 8132
rect 10813 8188 10877 8192
rect 10813 8132 10817 8188
rect 10817 8132 10873 8188
rect 10873 8132 10877 8188
rect 10813 8128 10877 8132
rect 10893 8188 10957 8192
rect 10893 8132 10897 8188
rect 10897 8132 10953 8188
rect 10953 8132 10957 8188
rect 10893 8128 10957 8132
rect 10973 8188 11037 8192
rect 10973 8132 10977 8188
rect 10977 8132 11033 8188
rect 11033 8132 11037 8188
rect 10973 8128 11037 8132
rect 11053 8188 11117 8192
rect 11053 8132 11057 8188
rect 11057 8132 11113 8188
rect 11113 8132 11117 8188
rect 11053 8128 11117 8132
rect 3417 7644 3481 7648
rect 3417 7588 3421 7644
rect 3421 7588 3477 7644
rect 3477 7588 3481 7644
rect 3417 7584 3481 7588
rect 3497 7644 3561 7648
rect 3497 7588 3501 7644
rect 3501 7588 3557 7644
rect 3557 7588 3561 7644
rect 3497 7584 3561 7588
rect 3577 7644 3641 7648
rect 3577 7588 3581 7644
rect 3581 7588 3637 7644
rect 3637 7588 3641 7644
rect 3577 7584 3641 7588
rect 3657 7644 3721 7648
rect 3657 7588 3661 7644
rect 3661 7588 3717 7644
rect 3717 7588 3721 7644
rect 3657 7584 3721 7588
rect 8348 7644 8412 7648
rect 8348 7588 8352 7644
rect 8352 7588 8408 7644
rect 8408 7588 8412 7644
rect 8348 7584 8412 7588
rect 8428 7644 8492 7648
rect 8428 7588 8432 7644
rect 8432 7588 8488 7644
rect 8488 7588 8492 7644
rect 8428 7584 8492 7588
rect 8508 7644 8572 7648
rect 8508 7588 8512 7644
rect 8512 7588 8568 7644
rect 8568 7588 8572 7644
rect 8508 7584 8572 7588
rect 8588 7644 8652 7648
rect 8588 7588 8592 7644
rect 8592 7588 8648 7644
rect 8648 7588 8652 7644
rect 8588 7584 8652 7588
rect 13278 7644 13342 7648
rect 13278 7588 13282 7644
rect 13282 7588 13338 7644
rect 13338 7588 13342 7644
rect 13278 7584 13342 7588
rect 13358 7644 13422 7648
rect 13358 7588 13362 7644
rect 13362 7588 13418 7644
rect 13418 7588 13422 7644
rect 13358 7584 13422 7588
rect 13438 7644 13502 7648
rect 13438 7588 13442 7644
rect 13442 7588 13498 7644
rect 13498 7588 13502 7644
rect 13438 7584 13502 7588
rect 13518 7644 13582 7648
rect 13518 7588 13522 7644
rect 13522 7588 13578 7644
rect 13578 7588 13582 7644
rect 13518 7584 13582 7588
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 6122 7100 6186 7104
rect 6122 7044 6126 7100
rect 6126 7044 6182 7100
rect 6182 7044 6186 7100
rect 6122 7040 6186 7044
rect 10813 7100 10877 7104
rect 10813 7044 10817 7100
rect 10817 7044 10873 7100
rect 10873 7044 10877 7100
rect 10813 7040 10877 7044
rect 10893 7100 10957 7104
rect 10893 7044 10897 7100
rect 10897 7044 10953 7100
rect 10953 7044 10957 7100
rect 10893 7040 10957 7044
rect 10973 7100 11037 7104
rect 10973 7044 10977 7100
rect 10977 7044 11033 7100
rect 11033 7044 11037 7100
rect 10973 7040 11037 7044
rect 11053 7100 11117 7104
rect 11053 7044 11057 7100
rect 11057 7044 11113 7100
rect 11113 7044 11117 7100
rect 11053 7040 11117 7044
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
<< metal4 >>
rect 3409 17440 3729 17456
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 16352 3729 17376
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 15264 3729 16288
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 14176 3729 15200
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 13088 3729 14112
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 12000 3729 13024
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 10912 3729 11936
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 9824 3729 10848
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 8736 3729 9760
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 7648 3729 8672
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 6560 3729 7584
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 5472 3729 6496
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 3296 3729 4320
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 2208 3729 3232
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 5874 16896 6195 17456
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6195 16896
rect 5874 15808 6195 16832
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6195 15808
rect 5874 14720 6195 15744
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6195 14720
rect 5874 13632 6195 14656
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6195 13632
rect 5874 12544 6195 13568
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6195 12544
rect 5874 11456 6195 12480
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6195 11456
rect 5874 10368 6195 11392
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6195 10368
rect 5874 9280 6195 10304
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6195 9280
rect 5874 8192 6195 9216
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6195 8192
rect 5874 7104 6195 8128
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6195 7104
rect 5874 6016 6195 7040
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5874 3840 6195 4864
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5874 2752 6195 3776
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 5874 2128 6195 2688
rect 8340 17440 8660 17456
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 16352 8660 17376
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 15264 8660 16288
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 14176 8660 15200
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 13088 8660 14112
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 12000 8660 13024
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 10912 8660 11936
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 9824 8660 10848
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 8736 8660 9760
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 7648 8660 8672
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 6560 8660 7584
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 5472 8660 6496
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 3296 8660 4320
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 2208 8660 3232
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 10805 16896 11125 17456
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 15808 11125 16832
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 14720 11125 15744
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 13632 11125 14656
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 12544 11125 13568
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 11456 11125 12480
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 10368 11125 11392
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 9280 11125 10304
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 8192 11125 9216
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 7104 11125 8128
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 6016 11125 7040
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 3840 11125 4864
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 2752 11125 3776
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2128 11125 2688
rect 13270 17440 13590 17456
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 13270 16352 13590 17376
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 15264 13590 16288
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 14176 13590 15200
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 13088 13590 14112
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 12000 13590 13024
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 10912 13590 11936
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 9824 13590 10848
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 8736 13590 9760
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 7648 13590 8672
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 6560 13590 7584
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 5472 13590 6496
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 3296 13590 4320
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 2208 13590 3232
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2128 13590 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606821651
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606821651
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1606821651
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1606821651
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606821651
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606821651
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1606821651
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606821651
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1606821651
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1606821651
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1606821651
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1606821651
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1606821651
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1606821651
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1606821651
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1606821651
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_147
timestamp 1606821651
transform 1 0 14628 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1606821651
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606821651
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606821651
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606821651
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1606821651
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1606821651
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1606821651
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1606821651
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1606821651
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1606821651
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1606821651
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606821651
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606821651
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606821651
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606821651
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606821651
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1606821651
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1606821651
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1606821651
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1606821651
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1606821651
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_147
timestamp 1606821651
transform 1 0 14628 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_155
timestamp 1606821651
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606821651
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606821651
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606821651
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1606821651
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1606821651
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1606821651
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1606821651
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1606821651
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1606821651
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1606821651
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606821651
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606821651
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606821651
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606821651
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606821651
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1606821651
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1606821651
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1606821651
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1606821651
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1606821651
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_147
timestamp 1606821651
transform 1 0 14628 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_155
timestamp 1606821651
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606821651
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606821651
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _37_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 4324 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1606821651
transform 1 0 3680 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606821651
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_27
timestamp 1606821651
transform 1 0 3588 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_32
timestamp 1606821651
transform 1 0 4048 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_39
timestamp 1606821651
transform 1 0 4692 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1606821651
transform 1 0 5152 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1606821651
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1606821651
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_43
timestamp 1606821651
transform 1 0 5060 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_48
timestamp 1606821651
transform 1 0 5520 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1606821651
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1606821651
transform 1 0 7544 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1606821651
transform 1 0 7728 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_68
timestamp 1606821651
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1606821651
transform 1 0 7912 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_70
timestamp 1606821651
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_76
timestamp 1606821651
transform 1 0 8096 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_88
timestamp 1606821651
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_86
timestamp 1606821651
transform 1 0 9016 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1606821651
transform 1 0 9384 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_103
timestamp 1606821651
transform 1 0 10580 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_98
timestamp 1606821651
transform 1 0 10120 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_94
timestamp 1606821651
transform 1 0 9752 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1606821651
transform 1 0 10212 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1606821651
transform 1 0 10028 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1606821651
transform 1 0 11500 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1606821651
transform 1 0 11132 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1606821651
transform 1 0 12236 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_111
timestamp 1606821651
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1606821651
transform 1 0 11868 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1606821651
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_133
timestamp 1606821651
transform 1 0 13340 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_145
timestamp 1606821651
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1606821651
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_147
timestamp 1606821651
transform 1 0 14628 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1606821651
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606821651
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1606821651
transform 1 0 4784 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606821651
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_32
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1606821651
transform 1 0 6808 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1606821651
transform 1 0 6256 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1606821651
transform 1 0 5612 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_44
timestamp 1606821651
transform 1 0 5152 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_48
timestamp 1606821651
transform 1 0 5520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp 1606821651
transform 1 0 5980 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_60
timestamp 1606821651
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1606821651
transform 1 0 8464 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1606821651
transform 1 0 7912 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1606821651
transform 1 0 7360 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_66
timestamp 1606821651
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_72
timestamp 1606821651
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_78
timestamp 1606821651
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _05_
timestamp 1606821651
transform 1 0 9936 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1606821651
transform 1 0 10672 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1606821651
transform 1 0 9016 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1606821651
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1606821651
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_100
timestamp 1606821651
transform 1 0 10304 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1606821651
transform 1 0 12512 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1606821651
transform 1 0 11408 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1606821651
transform 1 0 11960 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_108
timestamp 1606821651
transform 1 0 11040 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_116
timestamp 1606821651
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_122
timestamp 1606821651
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_128
timestamp 1606821651
transform 1 0 12880 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_140
timestamp 1606821651
transform 1 0 13984 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1606821651
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1606821651
transform 1 0 2484 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1606821651
transform 1 0 4876 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3220 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_29
timestamp 1606821651
transform 1 0 3772 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1606821651
transform 1 0 6164 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _15_
timestamp 1606821651
transform 1 0 5612 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1606821651
transform 1 0 5244 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1606821651
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606821651
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _09_
timestamp 1606821651
transform 1 0 8280 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _10_
timestamp 1606821651
transform 1 0 7728 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _11_
timestamp 1606821651
transform 1 0 7176 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_70
timestamp 1606821651
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_76
timestamp 1606821651
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_82
timestamp 1606821651
transform 1 0 8648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _04_
timestamp 1606821651
transform 1 0 10212 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _06_
timestamp 1606821651
transform 1 0 9476 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _07_
timestamp 1606821651
transform 1 0 8924 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_89
timestamp 1606821651
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1606821651
transform 1 0 9844 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_103
timestamp 1606821651
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _03_
timestamp 1606821651
transform 1 0 10764 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1606821651
transform 1 0 11592 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_109
timestamp 1606821651
transform 1 0 11132 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1606821651
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1606821651
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1606821651
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1606821651
transform 1 0 13892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_151
timestamp 1606821651
transform 1 0 14996 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606821651
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606821651
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1606821651
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_56
timestamp 1606821651
transform 1 0 6256 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1606821651
transform 1 0 6992 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1606821651
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1606821651
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1606821651
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1606821651
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1606821651
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1606821651
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1606821651
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1606821651
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1606821651
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1606821651
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606821651
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1606821651
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1606821651
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1606821651
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1606821651
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1606821651
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_147
timestamp 1606821651
transform 1 0 14628 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1606821651
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1606821651
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1606821651
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1606821651
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1606821651
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1606821651
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1606821651
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 12328 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1606821651
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_117
timestamp 1606821651
transform 1 0 11868 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_121
timestamp 1606821651
transform 1 0 12236 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_134
timestamp 1606821651
transform 1 0 13432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1606821651
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1606821651
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1606821651
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_16
timestamp 1606821651
transform 1 0 2576 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1606821651
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1606821651
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_28
timestamp 1606821651
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6256 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1606821651
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606821651
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1606821651
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 7268 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8280 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 7268 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_66
timestamp 1606821651
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_76
timestamp 1606821651
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_65
timestamp 1606821651
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_83
timestamp 1606821651
transform 1 0 8740 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _01_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_87
timestamp 1606821651
transform 1 0 9108 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_99
timestamp 1606821651
transform 1 0 10212 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1606821651
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_96
timestamp 1606821651
transform 1 0 9936 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_111
timestamp 1606821651
transform 1 0 11316 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1606821651
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_108
timestamp 1606821651
transform 1 0 11040 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_120
timestamp 1606821651
transform 1 0 12144 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1606821651
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_132
timestamp 1606821651
transform 1 0 13248 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_144
timestamp 1606821651
transform 1 0 14352 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_147
timestamp 1606821651
transform 1 0 14628 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1606821651
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1606821651
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_15
timestamp 1606821651
transform 1 0 2484 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3128 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606821651
transform 1 0 3956 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_15_21
timestamp 1606821651
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_25
timestamp 1606821651
transform 1 0 3404 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1606821651
transform 1 0 5152 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_56
timestamp 1606821651
transform 1 0 6256 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1606821651
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_62
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7636 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 7360 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 10304 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 9292 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_87
timestamp 1606821651
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1606821651
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_109
timestamp 1606821651
transform 1 0 11132 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1606821651
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1606821651
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_147
timestamp 1606821651
transform 1 0 14628 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1606821651
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1606821651
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606821651
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6256 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1606821651
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7268 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_65
timestamp 1606821651
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_83
timestamp 1606821651
transform 1 0 8740 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1606821651
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_102
timestamp 1606821651
transform 1 0 10488 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_114
timestamp 1606821651
transform 1 0 11592 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_126
timestamp 1606821651
transform 1 0 12696 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_138
timestamp 1606821651
transform 1 0 13800 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1606821651
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1606821651
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1606821651
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1606821651
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1606821651
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606821651
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7820 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1606821651
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_89
timestamp 1606821651
transform 1 0 9292 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_101
timestamp 1606821651
transform 1 0 10396 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1606821651
transform 1 0 11500 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1606821651
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1606821651
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_147
timestamp 1606821651
transform 1 0 14628 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1606821651
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606821651
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606821651
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6072 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_18_44
timestamp 1606821651
transform 1 0 5152 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1606821651
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 7912 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_83
timestamp 1606821651
transform 1 0 8740 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1606821651
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1606821651
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1606821651
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1606821651
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1606821651
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2852 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1606821651
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_15
timestamp 1606821651
transform 1 0 2484 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1606821651
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1606821651
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1606821651
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_32
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_40
timestamp 1606821651
transform 1 0 4784 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1606821651
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606821651
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1606821651
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1606821651
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_71
timestamp 1606821651
transform 1 0 7636 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_83
timestamp 1606821651
transform 1 0 8740 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1606821651
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1606821651
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_95
timestamp 1606821651
transform 1 0 9844 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_107
timestamp 1606821651
transform 1 0 10948 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_119
timestamp 1606821651
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1606821651
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1606821651
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1606821651
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1606821651
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1606821651
transform 1 0 14076 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1606821651
transform 1 0 14628 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_147
timestamp 1606821651
transform 1 0 14628 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1606821651
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1606821651
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1606821651
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4324 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_27
timestamp 1606821651
transform 1 0 3588 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1606821651
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606821651
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1606821651
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1606821651
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1606821651
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1606821651
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1606821651
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_147
timestamp 1606821651
transform 1 0 14628 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_155
timestamp 1606821651
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1606821651
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606821651
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1606821651
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1606821651
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1606821651
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1606821651
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1606821651
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1606821651
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1606821651
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1606821651
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1606821651
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1606821651
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1606821651
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1606821651
transform 1 0 4508 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1606821651
transform 1 0 3772 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_27
timestamp 1606821651
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_33
timestamp 1606821651
transform 1 0 4140 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_41
timestamp 1606821651
transform 1 0 4876 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1606821651
transform 1 0 5336 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_45
timestamp 1606821651
transform 1 0 5244 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_50
timestamp 1606821651
transform 1 0 5704 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_58
timestamp 1606821651
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_62
timestamp 1606821651
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1606821651
transform 1 0 7084 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1606821651
transform 1 0 7452 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1606821651
transform 1 0 8556 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _02_
timestamp 1606821651
transform 1 0 9292 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1606821651
transform 1 0 9660 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_105
timestamp 1606821651
transform 1 0 10764 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1606821651
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1606821651
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1606821651
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1606821651
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp 1606821651
transform 1 0 14628 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1606821651
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1606821651
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1606821651
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1606821651
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1606821651
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1606821651
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1606821651
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1606821651
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1606821651
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1606821651
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1606821651
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1606821651
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1606821651
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1606821651
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1606821651
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1606821651
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1606821651
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1606821651
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1606821651
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1606821651
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606821651
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1606821651
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1606821651
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1606821651
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1606821651
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1606821651
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1606821651
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1606821651
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_147
timestamp 1606821651
transform 1 0 14628 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1606821651
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1606821651
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1606821651
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1606821651
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1606821651
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1606821651
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1606821651
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1606821651
transform 1 0 3588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1606821651
transform 1 0 4048 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1606821651
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1606821651
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1606821651
transform 1 0 5152 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_56
timestamp 1606821651
transform 1 0 6256 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1606821651
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1606821651
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_63
timestamp 1606821651
transform 1 0 6900 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_75
timestamp 1606821651
transform 1 0 8004 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1606821651
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_87
timestamp 1606821651
transform 1 0 9108 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1606821651
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1606821651
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1606821651
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_106
timestamp 1606821651
transform 1 0 10856 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_118
timestamp 1606821651
transform 1 0 11960 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1606821651
transform 1 0 12604 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1606821651
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1606821651
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1606821651
transform 1 0 13708 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 15824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 15824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1606821651
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_149
timestamp 1606821651
transform 1 0 14812 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1606821651
transform 1 0 15456 0 1 16864
box -38 -48 130 592
<< labels >>
rlabel metal2 s 202 19520 258 20000 6 IO_ISOL_N
port 0 nsew default input
rlabel metal3 s 0 18232 480 18352 6 ccff_head
port 1 nsew default input
rlabel metal3 s 16520 12384 17000 12504 6 ccff_tail
port 2 nsew default tristate
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[0]
port 3 nsew default input
rlabel metal2 s 12898 0 12954 480 6 chany_bottom_in[10]
port 4 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[11]
port 5 nsew default input
rlabel metal2 s 13818 0 13874 480 6 chany_bottom_in[12]
port 6 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[13]
port 7 nsew default input
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_in[14]
port 8 nsew default input
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_in[15]
port 9 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_in[16]
port 10 nsew default input
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_in[17]
port 11 nsew default input
rlabel metal2 s 16302 0 16358 480 6 chany_bottom_in[18]
port 12 nsew default input
rlabel metal2 s 16762 0 16818 480 6 chany_bottom_in[19]
port 13 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[1]
port 14 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[2]
port 15 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[3]
port 16 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[4]
port 17 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[5]
port 18 nsew default input
rlabel metal2 s 11242 0 11298 480 6 chany_bottom_in[6]
port 19 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_in[7]
port 20 nsew default input
rlabel metal2 s 12070 0 12126 480 6 chany_bottom_in[8]
port 21 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[9]
port 22 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 23 nsew default tristate
rlabel metal2 s 4434 0 4490 480 6 chany_bottom_out[10]
port 24 nsew default tristate
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_out[11]
port 25 nsew default tristate
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_out[12]
port 26 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[13]
port 27 nsew default tristate
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_out[14]
port 28 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[15]
port 29 nsew default tristate
rlabel metal2 s 7010 0 7066 480 6 chany_bottom_out[16]
port 30 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[17]
port 31 nsew default tristate
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_out[18]
port 32 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_out[19]
port 33 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 34 nsew default tristate
rlabel metal2 s 1030 0 1086 480 6 chany_bottom_out[2]
port 35 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 36 nsew default tristate
rlabel metal2 s 1858 0 1914 480 6 chany_bottom_out[4]
port 37 nsew default tristate
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_out[5]
port 38 nsew default tristate
rlabel metal2 s 2686 0 2742 480 6 chany_bottom_out[6]
port 39 nsew default tristate
rlabel metal2 s 3146 0 3202 480 6 chany_bottom_out[7]
port 40 nsew default tristate
rlabel metal2 s 3606 0 3662 480 6 chany_bottom_out[8]
port 41 nsew default tristate
rlabel metal2 s 3974 0 4030 480 6 chany_bottom_out[9]
port 42 nsew default tristate
rlabel metal2 s 8850 19520 8906 20000 6 chany_top_in[0]
port 43 nsew default input
rlabel metal2 s 12990 19520 13046 20000 6 chany_top_in[10]
port 44 nsew default input
rlabel metal2 s 13450 19520 13506 20000 6 chany_top_in[11]
port 45 nsew default input
rlabel metal2 s 13818 19520 13874 20000 6 chany_top_in[12]
port 46 nsew default input
rlabel metal2 s 14278 19520 14334 20000 6 chany_top_in[13]
port 47 nsew default input
rlabel metal2 s 14646 19520 14702 20000 6 chany_top_in[14]
port 48 nsew default input
rlabel metal2 s 15106 19520 15162 20000 6 chany_top_in[15]
port 49 nsew default input
rlabel metal2 s 15474 19520 15530 20000 6 chany_top_in[16]
port 50 nsew default input
rlabel metal2 s 15934 19520 15990 20000 6 chany_top_in[17]
port 51 nsew default input
rlabel metal2 s 16302 19520 16358 20000 6 chany_top_in[18]
port 52 nsew default input
rlabel metal2 s 16762 19520 16818 20000 6 chany_top_in[19]
port 53 nsew default input
rlabel metal2 s 9310 19520 9366 20000 6 chany_top_in[1]
port 54 nsew default input
rlabel metal2 s 9678 19520 9734 20000 6 chany_top_in[2]
port 55 nsew default input
rlabel metal2 s 10138 19520 10194 20000 6 chany_top_in[3]
port 56 nsew default input
rlabel metal2 s 10506 19520 10562 20000 6 chany_top_in[4]
port 57 nsew default input
rlabel metal2 s 10966 19520 11022 20000 6 chany_top_in[5]
port 58 nsew default input
rlabel metal2 s 11334 19520 11390 20000 6 chany_top_in[6]
port 59 nsew default input
rlabel metal2 s 11794 19520 11850 20000 6 chany_top_in[7]
port 60 nsew default input
rlabel metal2 s 12162 19520 12218 20000 6 chany_top_in[8]
port 61 nsew default input
rlabel metal2 s 12622 19520 12678 20000 6 chany_top_in[9]
port 62 nsew default input
rlabel metal2 s 570 19520 626 20000 6 chany_top_out[0]
port 63 nsew default tristate
rlabel metal2 s 4710 19520 4766 20000 6 chany_top_out[10]
port 64 nsew default tristate
rlabel metal2 s 5170 19520 5226 20000 6 chany_top_out[11]
port 65 nsew default tristate
rlabel metal2 s 5538 19520 5594 20000 6 chany_top_out[12]
port 66 nsew default tristate
rlabel metal2 s 5998 19520 6054 20000 6 chany_top_out[13]
port 67 nsew default tristate
rlabel metal2 s 6366 19520 6422 20000 6 chany_top_out[14]
port 68 nsew default tristate
rlabel metal2 s 6826 19520 6882 20000 6 chany_top_out[15]
port 69 nsew default tristate
rlabel metal2 s 7194 19520 7250 20000 6 chany_top_out[16]
port 70 nsew default tristate
rlabel metal2 s 7654 19520 7710 20000 6 chany_top_out[17]
port 71 nsew default tristate
rlabel metal2 s 8022 19520 8078 20000 6 chany_top_out[18]
port 72 nsew default tristate
rlabel metal2 s 8482 19520 8538 20000 6 chany_top_out[19]
port 73 nsew default tristate
rlabel metal2 s 1030 19520 1086 20000 6 chany_top_out[1]
port 74 nsew default tristate
rlabel metal2 s 1398 19520 1454 20000 6 chany_top_out[2]
port 75 nsew default tristate
rlabel metal2 s 1858 19520 1914 20000 6 chany_top_out[3]
port 76 nsew default tristate
rlabel metal2 s 2226 19520 2282 20000 6 chany_top_out[4]
port 77 nsew default tristate
rlabel metal2 s 2686 19520 2742 20000 6 chany_top_out[5]
port 78 nsew default tristate
rlabel metal2 s 3054 19520 3110 20000 6 chany_top_out[6]
port 79 nsew default tristate
rlabel metal2 s 3514 19520 3570 20000 6 chany_top_out[7]
port 80 nsew default tristate
rlabel metal2 s 3882 19520 3938 20000 6 chany_top_out[8]
port 81 nsew default tristate
rlabel metal2 s 4342 19520 4398 20000 6 chany_top_out[9]
port 82 nsew default tristate
rlabel metal3 s 0 8304 480 8424 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 83 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 84 nsew default input
rlabel metal3 s 0 14968 480 15088 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 85 nsew default tristate
rlabel metal3 s 0 4904 480 5024 6 left_grid_pin_0_
port 86 nsew default tristate
rlabel metal3 s 16520 7352 17000 7472 6 prog_clk_0_E_in
port 87 nsew default input
rlabel metal3 s 0 1640 480 1760 6 right_width_0_height_0__pin_0_
port 88 nsew default input
rlabel metal3 s 16520 2456 17000 2576 6 right_width_0_height_0__pin_1_lower
port 89 nsew default tristate
rlabel metal3 s 16520 17416 17000 17536 6 right_width_0_height_0__pin_1_upper
port 90 nsew default tristate
rlabel metal4 s 3409 2128 3729 17456 6 VPWR
port 91 nsew default input
rlabel metal4 s 5875 2128 6195 17456 6 VGND
port 92 nsew default input
<< properties >>
string FIXED_BBOX 0 0 17000 20000
<< end >>
