* NGSPICE file created from grid_io_bottom.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_1 abstract view
.subckt scs8hd_ebufn_1 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_and4_4 abstract view
.subckt scs8hd_and4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

.subckt grid_io_bottom address[0] address[1] address[2] address[3] data_in enable
+ gfpga_pad_GPIO_PAD[0] gfpga_pad_GPIO_PAD[1] gfpga_pad_GPIO_PAD[2] gfpga_pad_GPIO_PAD[3]
+ gfpga_pad_GPIO_PAD[4] gfpga_pad_GPIO_PAD[5] gfpga_pad_GPIO_PAD[6] gfpga_pad_GPIO_PAD[7]
+ top_width_0_height_0__pin_0_ top_width_0_height_0__pin_10_ top_width_0_height_0__pin_11_
+ top_width_0_height_0__pin_12_ top_width_0_height_0__pin_13_ top_width_0_height_0__pin_14_
+ top_width_0_height_0__pin_15_ top_width_0_height_0__pin_1_ top_width_0_height_0__pin_2_
+ top_width_0_height_0__pin_3_ top_width_0_height_0__pin_4_ top_width_0_height_0__pin_5_
+ top_width_0_height_0__pin_6_ top_width_0_height_0__pin_7_ top_width_0_height_0__pin_8_
+ top_width_0_height_0__pin_9_ vpwr vgnd
XFILLER_7_1880 vgnd vpwr scs8hd_decap_8
XFILLER_3_2489 vgnd vpwr scs8hd_decap_12
XFILLER_3_1733 vgnd vpwr scs8hd_decap_12
XFILLER_8_3057 vgnd vpwr scs8hd_decap_12
XFILLER_8_2301 vgnd vpwr scs8hd_decap_12
XFILLER_8_2345 vgnd vpwr scs8hd_decap_4
XFILLER_8_1666 vgnd vpwr scs8hd_decap_12
XFILLER_5_3978 vgnd vpwr scs8hd_decap_12
XFILLER_4_1508 vgnd vpwr scs8hd_decap_12
XFILLER_3_2990 vgnd vpwr scs8hd_decap_12
XFILLER_2_1276 vgnd vpwr scs8hd_decap_12
XFILLER_9_137 vgnd vpwr scs8hd_decap_12
XFILLER_6_800 vgnd vpwr scs8hd_decap_12
XFILLER_9_2109 vgnd vpwr scs8hd_decap_12
XFILLER_9_1408 vgnd vpwr scs8hd_decap_12
XFILLER_5_354 vgnd vpwr scs8hd_decap_12
XFILLER_4_4167 vgnd vpwr scs8hd_decap_12
XFILLER_4_3411 vgnd vpwr scs8hd_decap_12
XFILLER_0_2629 vgnd vpwr scs8hd_decap_6
XFILLER_9_4012 vgnd vpwr scs8hd_decap_12
XFILLER_9_3311 vgnd vpwr scs8hd_decap_6
XFILLER_9_2698 vgnd vpwr scs8hd_decap_12
XFILLER_9_1997 vgnd vpwr scs8hd_decap_12
XFILLER_9_1931 vgnd vpwr scs8hd_decap_12
XFILLER_5_1806 vgnd vpwr scs8hd_decap_12
XPHY_905 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_2297 vpwr vgnd scs8hd_fill_2
XFILLER_3_1574 vgnd vpwr scs8hd_decap_12
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XFILLER_8_2142 vgnd vpwr scs8hd_decap_12
XFILLER_5_4454 vgnd vpwr scs8hd_decap_12
XFILLER_1_4307 vgnd vpwr scs8hd_decap_12
XFILLER_2_324 vgnd vpwr scs8hd_decap_12
XFILLER_8_1496 vgnd vpwr scs8hd_decap_12
XFILLER_4_1349 vgnd vpwr scs8hd_decap_12
XFILLER_1_2916 vgnd vpwr scs8hd_decap_12
XFILLER_6_2838 vgnd vpwr scs8hd_decap_12
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XFILLER_4_3252 vgnd vpwr scs8hd_decap_12
XFILLER_9_3163 vgnd vpwr scs8hd_decap_12
XFILLER_9_2462 vgnd vpwr scs8hd_decap_12
XFILLER_9_490 vgnd vpwr scs8hd_decap_6
XFILLER_5_3038 vgnd vpwr scs8hd_decap_12
XFILLER_9_1761 vgnd vpwr scs8hd_decap_6
XFILLER_3_2050 vgnd vpwr scs8hd_decap_12
XFILLER_0_4384 vgnd vpwr scs8hd_decap_12
XFILLER_2_3948 vgnd vpwr scs8hd_decap_12
XPHY_768 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_757 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_746 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_735 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_724 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_713 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_702 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_3683 vgnd vpwr scs8hd_decap_6
XPHY_779 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4527 vgnd vpwr scs8hd_decap_12
XFILLER_3_611 vgnd vpwr scs8hd_decap_12
XFILLER_5_4295 vgnd vpwr scs8hd_decap_12
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XFILLER_1_2746 vgnd vpwr scs8hd_decap_12
XFILLER_9_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_471 vgnd vpwr scs8hd_decap_12
XFILLER_9_1079 vgnd vpwr scs8hd_decap_6
XFILLER_9_1024 vgnd vpwr scs8hd_decap_12
XFILLER_6_2679 vgnd vpwr scs8hd_decap_12
XFILLER_6_1923 vgnd vpwr scs8hd_decap_12
XFILLER_4_3082 vgnd vpwr scs8hd_decap_12
XFILLER_4_1691 vgnd vpwr scs8hd_decap_12
XFILLER_0_1544 vgnd vpwr scs8hd_decap_6
XFILLER_0_2245 vgnd vpwr scs8hd_decap_12
XFILLER_7_1709 vgnd vpwr scs8hd_decap_12
XFILLER_5_2123 vgnd vpwr scs8hd_decap_12
XFILLER_2_4424 vgnd vpwr scs8hd_decap_12
XFILLER_0_614 vgnd vpwr scs8hd_decap_6
XFILLER_5_1477 vgnd vpwr scs8hd_decap_12
XFILLER_2_3789 vgnd vpwr scs8hd_decap_12
XFILLER_8_703 vgnd vpwr scs8hd_decap_12
XPHY_598 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_587 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_576 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_565 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_554 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_543 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_532 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_521 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_510 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4368 vgnd vpwr scs8hd_decap_12
XFILLER_7_3612 vgnd vpwr scs8hd_decap_12
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XFILLER_3_452 vgnd vpwr scs8hd_decap_12
XFILLER_7_2977 vgnd vpwr scs8hd_decap_12
XFILLER_5_3380 vgnd vpwr scs8hd_decap_12
XFILLER_3_2819 vgnd vpwr scs8hd_decap_12
XFILLER_1_1831 vgnd vpwr scs8hd_decap_12
XFILLER_1_2587 vgnd vpwr scs8hd_decap_12
XFILLER_6_3155 vgnd vpwr scs8hd_decap_12
XFILLER_2_3008 vgnd vpwr scs8hd_decap_12
XFILLER_6_1764 vgnd vpwr scs8hd_decap_12
XFILLER_1_4490 vgnd vpwr scs8hd_decap_12
XFILLER_0_1396 vgnd vpwr scs8hd_decap_12
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_2_4265 vgnd vpwr scs8hd_decap_12
XFILLER_1_989 vgnd vpwr scs8hd_decap_12
XFILLER_0_466 vgnd vpwr scs8hd_decap_12
XFILLER_2_2874 vgnd vpwr scs8hd_decap_12
XFILLER_8_544 vgnd vpwr scs8hd_decap_12
XPHY_395 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_384 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_373 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_362 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_351 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_340 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3453 vgnd vpwr scs8hd_decap_12
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XFILLER_3_293 vgnd vpwr scs8hd_decap_12
XFILLER_3_1904 vgnd vpwr scs8hd_decap_12
XFILLER_1_2362 vgnd vpwr scs8hd_decap_8
XFILLER_1_3063 vgnd vpwr scs8hd_decap_12
XFILLER_1_1672 vgnd vpwr scs8hd_decap_12
XFILLER_8_3228 vgnd vpwr scs8hd_decap_12
XFILLER_8_1837 vgnd vpwr scs8hd_decap_4
XFILLER_6_2240 vgnd vpwr scs8hd_decap_12
XFILLER_3_4563 vgnd vpwr scs8hd_decap_12
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_1160 vgnd vpwr scs8hd_decap_12
XFILLER_2_1447 vgnd vpwr scs8hd_decap_12
XFILLER_8_4485 vgnd vpwr scs8hd_decap_12
XFILLER_8_3740 vgnd vpwr scs8hd_decap_12
XFILLER_7_2026 vgnd vpwr scs8hd_decap_12
XFILLER_5_525 vgnd vpwr scs8hd_decap_12
XFILLER_4_4338 vgnd vpwr scs8hd_decap_12
XFILLER_1_720 vgnd vpwr scs8hd_decap_12
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XFILLER_4_2947 vgnd vpwr scs8hd_decap_12
XFILLER_2_3350 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3504 vgnd vpwr scs8hd_decap_12
XFILLER_9_2803 vgnd vpwr scs8hd_decap_12
XFILLER_9_831 vgnd vpwr scs8hd_decap_6
XFILLER_8_385 vgnd vpwr scs8hd_decap_12
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3559 vgnd vpwr scs8hd_decap_6
XFILLER_3_3136 vgnd vpwr scs8hd_decap_12
XFILLER_7_1892 vgnd vpwr scs8hd_decap_12
XFILLER_3_1745 vgnd vpwr scs8hd_decap_12
XFILLER_8_3069 vgnd vpwr scs8hd_decap_12
XFILLER_8_2313 vgnd vpwr scs8hd_decap_12
XFILLER_6_2081 vgnd vpwr scs8hd_decap_12
XFILLER_3_4393 vgnd vpwr scs8hd_decap_12
XFILLER_2_1288 vgnd vpwr scs8hd_decap_12
XFILLER_9_149 vgnd vpwr scs8hd_decap_6
XFILLER_6_812 vgnd vpwr scs8hd_decap_12
XFILLER_8_3570 vgnd vpwr scs8hd_decap_12
XFILLER_7_1111 vgnd vpwr scs8hd_decap_12
XFILLER_4_3423 vgnd vpwr scs8hd_decap_12
XFILLER_1_550 vgnd vpwr scs8hd_decap_12
XFILLER_4_2777 vgnd vpwr scs8hd_decap_12
XFILLER_2_3191 vgnd vpwr scs8hd_decap_12
XFILLER_9_4024 vgnd vpwr scs8hd_decap_6
XFILLER_9_683 vgnd vpwr scs8hd_decap_12
XFILLER_5_3209 vgnd vpwr scs8hd_decap_12
XFILLER_9_1954 vgnd vpwr scs8hd_decap_12
XFILLER_9_1943 vgnd vpwr scs8hd_decap_8
XFILLER_5_1818 vgnd vpwr scs8hd_decap_12
XFILLER_3_2221 vgnd vpwr scs8hd_decap_12
XPHY_906 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_3876 vgnd vpwr scs8hd_decap_12
XFILLER_8_2154 vgnd vpwr scs8hd_decap_12
XFILLER_5_4466 vgnd vpwr scs8hd_decap_12
XFILLER_1_4319 vgnd vpwr scs8hd_decap_12
XFILLER_6_642 vgnd vpwr scs8hd_decap_12
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XFILLER_1_391 vgnd vpwr scs8hd_decap_12
XFILLER_4_1862 vgnd vpwr scs8hd_decap_12
XFILLER_0_1737 vgnd vpwr scs8hd_decap_12
XFILLER_9_3175 vgnd vpwr scs8hd_decap_12
XFILLER_9_2485 vpwr vgnd scs8hd_fill_2
XFILLER_9_2474 vgnd vpwr scs8hd_decap_6
XFILLER_0_807 vgnd vpwr scs8hd_decap_12
XFILLER_5_1648 vgnd vpwr scs8hd_decap_12
XFILLER_3_2062 vgnd vpwr scs8hd_decap_12
XFILLER_0_3640 vgnd vpwr scs8hd_decap_12
XFILLER_0_4341 vgnd vpwr scs8hd_decap_12
XFILLER_0_4396 vgnd vpwr scs8hd_decap_6
XPHY_769 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_758 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_747 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_736 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_725 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_714 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_703 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4539 vgnd vpwr scs8hd_decap_12
XFILLER_7_428 vgnd vpwr scs8hd_decap_12
XFILLER_3_623 vgnd vpwr scs8hd_decap_12
XFILLER_5_3551 vgnd vpwr scs8hd_decap_12
XFILLER_1_3404 vgnd vpwr scs8hd_decap_12
XFILLER_1_4149 vgnd vpwr scs8hd_decap_12
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XFILLER_1_2758 vgnd vpwr scs8hd_decap_12
XFILLER_9_56 vgnd vpwr scs8hd_decap_6
XFILLER_7_940 vgnd vpwr scs8hd_decap_6
XFILLER_9_1036 vgnd vpwr scs8hd_decap_12
XFILLER_6_3326 vgnd vpwr scs8hd_decap_12
XFILLER_7_973 vgnd vpwr scs8hd_decap_3
XFILLER_6_483 vgnd vpwr scs8hd_decap_12
XFILLER_6_1935 vgnd vpwr scs8hd_decap_12
XFILLER_4_3094 vgnd vpwr scs8hd_decap_12
XFILLER_0_1501 vgnd vpwr scs8hd_decap_12
XFILLER_0_2202 vgnd vpwr scs8hd_decap_12
XFILLER_0_2257 vgnd vpwr scs8hd_decap_6
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _10_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_4436 vgnd vpwr scs8hd_decap_12
XPHY_500 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_1489 vgnd vpwr scs8hd_decap_12
XFILLER_0_2791 vgnd vpwr scs8hd_decap_12
XFILLER_8_715 vgnd vpwr scs8hd_decap_12
XPHY_599 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_588 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_577 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_566 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_555 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_544 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_533 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_522 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_511 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3624 vgnd vpwr scs8hd_decap_12
XFILLER_7_269 vgnd vpwr scs8hd_decap_12
XFILLER_4_910 vgnd vpwr scs8hd_decap_12
XFILLER_3_464 vgnd vpwr scs8hd_decap_12
XFILLER_5_3392 vgnd vpwr scs8hd_decap_12
XFILLER_1_3234 vgnd vpwr scs8hd_decap_12
XFILLER_1_1843 vgnd vpwr scs8hd_decap_12
XFILLER_1_2599 vgnd vpwr scs8hd_decap_12
XFILLER_7_781 vgnd vpwr scs8hd_decap_12
XFILLER_6_3167 vgnd vpwr scs8hd_decap_12
XFILLER_6_2411 vgnd vpwr scs8hd_decap_12
XFILLER_6_1776 vgnd vpwr scs8hd_decap_12
XFILLER_2_1618 vgnd vpwr scs8hd_decap_12
XFILLER_8_3911 vgnd vpwr scs8hd_decap_12
XFILLER_4_4509 vgnd vpwr scs8hd_decap_12
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_9_2090 vgnd vpwr scs8hd_decap_12
XFILLER_2_4277 vgnd vpwr scs8hd_decap_12
XFILLER_0_478 vgnd vpwr scs8hd_decap_12
XFILLER_2_3521 vgnd vpwr scs8hd_decap_12
XPHY_352 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_341 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_330 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_2886 vgnd vpwr scs8hd_decap_12
XFILLER_8_556 vgnd vpwr scs8hd_decap_12
XFILLER_7_4100 vgnd vpwr scs8hd_decap_12
XPHY_396 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_385 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_374 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_363 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3465 vgnd vpwr scs8hd_decap_12
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XFILLER_4_751 vgnd vpwr scs8hd_decap_12
XFILLER_3_3307 vgnd vpwr scs8hd_decap_12
XFILLER_3_1916 vgnd vpwr scs8hd_decap_12
XFILLER_1_3075 vgnd vpwr scs8hd_decap_12
XFILLER_1_1684 vgnd vpwr scs8hd_decap_12
XFILLER_6_2252 vgnd vpwr scs8hd_decap_12
XFILLER_0_1172 vgnd vpwr scs8hd_decap_6
XFILLER_2_1459 vgnd vpwr scs8hd_decap_12
XFILLER_5_537 vgnd vpwr scs8hd_decap_12
XFILLER_8_4497 vgnd vpwr scs8hd_decap_12
XFILLER_7_2038 vgnd vpwr scs8hd_decap_12
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XFILLER_5_1050 vgnd vpwr scs8hd_decap_12
XFILLER_2_1971 vgnd vpwr scs8hd_decap_12
XFILLER_2_3362 vgnd vpwr scs8hd_decap_12
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_4217 vgnd vpwr scs8hd_decap_12
XFILLER_9_3516 vgnd vpwr scs8hd_decap_12
XFILLER_9_2815 vgnd vpwr scs8hd_decap_6
XFILLER_7_3295 vgnd vpwr scs8hd_decap_12
XFILLER_7_2550 vgnd vpwr scs8hd_decap_12
XFILLER_4_581 vgnd vpwr scs8hd_decap_12
XFILLER_3_3148 vgnd vpwr scs8hd_decap_12
XFILLER_3_1757 vgnd vpwr scs8hd_decap_12
XFILLER_1_2160 vgnd vpwr scs8hd_decap_12
XFILLER_8_2325 vgnd vpwr scs8hd_decap_6
XFILLER_2_507 vgnd vpwr scs8hd_decap_12
XFILLER_8_1679 vgnd vpwr scs8hd_decap_12
XFILLER_6_2093 vgnd vpwr scs8hd_decap_12
XFILLER_9_106 vgnd vpwr scs8hd_decap_12
XFILLER_5_367 vgnd vpwr scs8hd_decap_12
XFILLER_8_3582 vgnd vpwr scs8hd_decap_12
XFILLER_7_1123 vgnd vpwr scs8hd_decap_12
XFILLER_4_3435 vgnd vpwr scs8hd_decap_12
XFILLER_1_562 vgnd vpwr scs8hd_decap_12
XFILLER_4_2789 vgnd vpwr scs8hd_decap_12
XFILLER_9_695 vgnd vpwr scs8hd_decap_12
XFILLER_9_2667 vgnd vpwr scs8hd_decap_12
XFILLER_9_1966 vgnd vpwr scs8hd_decap_12
XFILLER_7_2380 vgnd vpwr scs8hd_decap_12
XFILLER_3_2233 vgnd vpwr scs8hd_decap_12
XFILLER_0_3888 vgnd vpwr scs8hd_decap_12
XFILLER_0_4578 vgnd vpwr scs8hd_decap_3
XPHY_907 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1587 vgnd vpwr scs8hd_decap_12
XFILLER_9_4570 vgnd vpwr scs8hd_decap_8
XFILLER_8_1410 vgnd vpwr scs8hd_decap_12
XFILLER_5_4478 vgnd vpwr scs8hd_decap_12
XFILLER_5_3722 vgnd vpwr scs8hd_decap_12
XFILLER_4_2008 vgnd vpwr scs8hd_decap_12
XFILLER_2_337 vgnd vpwr scs8hd_decap_12
XFILLER_3_3490 vgnd vpwr scs8hd_decap_12
XFILLER_1_2929 vgnd vpwr scs8hd_decap_12
XFILLER_2_1020 vgnd vpwr scs8hd_decap_12
XFILLER_6_654 vgnd vpwr scs8hd_decap_12
XFILLER_4_3265 vgnd vpwr scs8hd_decap_12
XFILLER_4_2520 vgnd vpwr scs8hd_decap_12
XFILLER_0_2417 vgnd vpwr scs8hd_fill_1
XFILLER_4_1874 vgnd vpwr scs8hd_decap_12
XFILLER_0_1749 vgnd vpwr scs8hd_decap_12
XFILLER_9_3187 vgnd vpwr scs8hd_decap_6
XFILLER_9_3132 vgnd vpwr scs8hd_decap_12
XFILLER_9_2431 vgnd vpwr scs8hd_decap_12
XFILLER_9_1730 vgnd vpwr scs8hd_decap_6
XFILLER_5_2306 vgnd vpwr scs8hd_decap_8
XFILLER_0_819 vgnd vpwr scs8hd_decap_12
XFILLER_0_3652 vgnd vpwr scs8hd_decap_6
XFILLER_0_4353 vgnd vpwr scs8hd_decap_12
XPHY_759 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_748 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_737 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_726 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_715 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_704 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_635 vgnd vpwr scs8hd_decap_12
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_3563 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_9_1048 vgnd vpwr scs8hd_decap_6
XFILLER_9_1004 vgnd vpwr scs8hd_decap_12
XFILLER_6_3338 vgnd vpwr scs8hd_decap_12
XFILLER_6_495 vgnd vpwr scs8hd_decap_12
XFILLER_2_690 vgnd vpwr scs8hd_decap_12
XFILLER_6_1947 vgnd vpwr scs8hd_decap_12
XFILLER_4_2350 vgnd vpwr scs8hd_decap_6
XFILLER_0_1513 vgnd vpwr scs8hd_decap_6
XFILLER_0_2214 vgnd vpwr scs8hd_decap_12
XFILLER_9_1582 vgnd vpwr scs8hd_decap_12
XFILLER_6_3850 vgnd vpwr scs8hd_decap_12
XFILLER_5_2136 vgnd vpwr scs8hd_decap_12
XFILLER_2_4448 vgnd vpwr scs8hd_decap_12
XPHY_534 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_523 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_512 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_501 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_727 vgnd vpwr scs8hd_decap_12
XPHY_589 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_578 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_567 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_556 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_545 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3636 vgnd vpwr scs8hd_decap_12
XFILLER_4_922 vgnd vpwr scs8hd_decap_12
XFILLER_3_476 vgnd vpwr scs8hd_decap_12
XFILLER_8_1081 vgnd vpwr scs8hd_decap_12
XFILLER_1_3246 vgnd vpwr scs8hd_decap_12
XFILLER_1_1855 vgnd vpwr scs8hd_decap_12
XFILLER_6_3179 vgnd vpwr scs8hd_decap_12
XFILLER_6_2423 vgnd vpwr scs8hd_decap_12
XFILLER_6_1788 vgnd vpwr scs8hd_decap_12
XFILLER_4_2191 vgnd vpwr scs8hd_decap_12
XFILLER_0_1365 vgnd vpwr scs8hd_decap_12
XFILLER_5_708 vgnd vpwr scs8hd_decap_12
XFILLER_8_3923 vgnd vpwr scs8hd_decap_12
XFILLER_7_2209 vgnd vpwr scs8hd_decap_12
XFILLER_1_903 vgnd vpwr scs8hd_decap_12
XFILLER_0_435 vgnd vpwr scs8hd_decap_12
XFILLER_5_1221 vgnd vpwr scs8hd_decap_12
XFILLER_2_4289 vgnd vpwr scs8hd_decap_12
XFILLER_2_3533 vgnd vpwr scs8hd_decap_12
XPHY_386 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_375 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_364 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_353 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_342 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_331 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_320 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_568 vgnd vpwr scs8hd_decap_12
XFILLER_7_4112 vgnd vpwr scs8hd_decap_12
XPHY_397 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_2721 vgnd vpwr scs8hd_decap_12
XFILLER_3_3319 vgnd vpwr scs8hd_decap_12
XFILLER_3_1928 vgnd vpwr scs8hd_decap_12
XFILLER_1_1696 vgnd vpwr scs8hd_decap_12
XFILLER_1_2375 vpwr vgnd scs8hd_fill_2
XFILLER_1_3087 vgnd vpwr scs8hd_decap_12
XFILLER_6_2264 vgnd vpwr scs8hd_decap_12
XFILLER_3_4576 vgnd vpwr scs8hd_decap_4
XFILLER_3_3831 vgnd vpwr scs8hd_decap_12
XFILLER_2_2106 vgnd vpwr scs8hd_decap_12
XANTENNA__04__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_8_3753 vgnd vpwr scs8hd_decap_12
XFILLER_4_3606 vgnd vpwr scs8hd_decap_12
XFILLER_1_733 vgnd vpwr scs8hd_decap_12
XFILLER_5_1062 vgnd vpwr scs8hd_decap_12
XFILLER_2_3374 vgnd vpwr scs8hd_decap_12
XFILLER_9_800 vgnd vpwr scs8hd_decap_6
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_4229 vgnd vpwr scs8hd_decap_12
XFILLER_9_3528 vgnd vpwr scs8hd_decap_6
XFILLER_8_398 vgnd vpwr scs8hd_decap_12
XFILLER_4_593 vgnd vpwr scs8hd_decap_12
XFILLER_3_2404 vgnd vpwr scs8hd_decap_12
XFILLER_1_2172 vgnd vpwr scs8hd_decap_12
XFILLER_3_3661 vgnd vpwr scs8hd_decap_12
XFILLER_9_118 vgnd vpwr scs8hd_decap_6
XFILLER_6_825 vgnd vpwr scs8hd_decap_12
XFILLER_5_379 vgnd vpwr scs8hd_decap_12
XFILLER_8_3594 vgnd vpwr scs8hd_decap_12
XFILLER_7_1135 vgnd vpwr scs8hd_decap_12
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_574 vgnd vpwr scs8hd_decap_12
XFILLER_9_652 vgnd vpwr scs8hd_decap_12
XFILLER_9_2679 vgnd vpwr scs8hd_decap_12
XFILLER_5_891 vgnd vpwr scs8hd_decap_12
XFILLER_9_1978 vgnd vpwr scs8hd_decap_6
XFILLER_7_2392 vgnd vpwr scs8hd_decap_12
XFILLER_3_2245 vgnd vpwr scs8hd_decap_12
XFILLER_3_1599 vgnd vpwr scs8hd_decap_12
XFILLER_0_3845 vgnd vpwr scs8hd_decap_12
XPHY_908 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_806 vgnd vpwr scs8hd_decap_12
XFILLER_8_2167 vgnd vpwr scs8hd_decap_12
XFILLER_8_1422 vgnd vpwr scs8hd_decap_12
XFILLER_5_3734 vgnd vpwr scs8hd_decap_12
XFILLER_2_349 vgnd vpwr scs8hd_decap_12
XFILLER_2_1032 vgnd vpwr scs8hd_decap_12
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XFILLER_8_4070 vgnd vpwr scs8hd_decap_12
XFILLER_6_3509 vgnd vpwr scs8hd_decap_12
XFILLER_6_666 vgnd vpwr scs8hd_decap_12
XFILLER_2_861 vgnd vpwr scs8hd_decap_12
XFILLER_4_3277 vgnd vpwr scs8hd_decap_12
XFILLER_4_1886 vgnd vpwr scs8hd_decap_12
XFILLER_0_1706 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ top_width_0_height_0__pin_8_ logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[4] vgnd vpwr scs8hd_ebufn_1
XFILLER_9_3144 vgnd vpwr scs8hd_decap_12
XFILLER_9_2443 vgnd vpwr scs8hd_decap_6
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XFILLER_0_4310 vgnd vpwr scs8hd_decap_12
XFILLER_0_4365 vgnd vpwr scs8hd_decap_6
XPHY_727 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_716 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_705 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_2075 vgnd vpwr scs8hd_decap_12
XFILLER_3_1330 vgnd vpwr scs8hd_decap_12
XPHY_749 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_738 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3807 vgnd vpwr scs8hd_decap_12
XFILLER_5_4210 vgnd vpwr scs8hd_decap_12
XFILLER_3_647 vgnd vpwr scs8hd_decap_12
XANTENNA__12__A _10_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_1252 vgnd vpwr scs8hd_decap_12
XFILLER_5_3575 vgnd vpwr scs8hd_decap_12
XFILLER_4_1105 vgnd vpwr scs8hd_decap_12
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_3417 vgnd vpwr scs8hd_decap_12
XFILLER_7_953 vgnd vpwr scs8hd_decap_12
XFILLER_9_1016 vgnd vpwr scs8hd_decap_6
XFILLER_6_1959 vgnd vpwr scs8hd_decap_12
XFILLER_4_2384 vgnd vpwr scs8hd_fill_1
XFILLER_0_2226 vgnd vpwr scs8hd_decap_6
XFILLER_9_2295 vgnd vpwr scs8hd_decap_12
XFILLER_9_1594 vgnd vpwr scs8hd_decap_12
XFILLER_6_3862 vgnd vpwr scs8hd_decap_12
XFILLER_5_2148 vgnd vpwr scs8hd_decap_12
XFILLER_2_3704 vgnd vpwr scs8hd_decap_12
XPHY_568 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_557 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_546 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_535 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_524 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_513 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_502 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__07__A _13_/C vgnd vpwr scs8hd_diode_2
XFILLER_3_1160 vgnd vpwr scs8hd_decap_12
XFILLER_0_2760 vgnd vpwr scs8hd_decap_12
XFILLER_8_739 vgnd vpwr scs8hd_decap_12
XPHY_579 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_934 vgnd vpwr scs8hd_decap_12
XFILLER_7_3648 vgnd vpwr scs8hd_decap_12
XFILLER_5_4051 vgnd vpwr scs8hd_decap_12
XFILLER_8_1093 vgnd vpwr scs8hd_decap_12
XFILLER_5_2660 vgnd vpwr scs8hd_decap_12
XFILLER_1_1867 vgnd vpwr scs8hd_decap_12
XFILLER_1_2502 vgnd vpwr scs8hd_decap_12
XFILLER_1_3258 vgnd vpwr scs8hd_decap_12
XFILLER_7_794 vgnd vpwr scs8hd_decap_12
XFILLER_6_2435 vgnd vpwr scs8hd_decap_12
XFILLER_1_3770 vgnd vpwr scs8hd_decap_12
XFILLER_0_1377 vgnd vpwr scs8hd_decap_12
XFILLER_0_2078 vgnd vpwr scs8hd_decap_12
XFILLER_6_3692 vgnd vpwr scs8hd_decap_12
XFILLER_0_447 vgnd vpwr scs8hd_decap_12
XFILLER_5_1233 vgnd vpwr scs8hd_decap_12
XFILLER_0_3280 vgnd vpwr scs8hd_decap_6
XFILLER_2_2899 vgnd vpwr scs8hd_decap_12
XFILLER_2_3545 vgnd vpwr scs8hd_decap_12
XPHY_398 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_387 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_376 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_365 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_354 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_343 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_332 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_321 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_310 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4124 vgnd vpwr scs8hd_decap_12
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_764 vgnd vpwr scs8hd_decap_12
XFILLER_7_3478 vgnd vpwr scs8hd_decap_12
XFILLER_7_2733 vgnd vpwr scs8hd_decap_12
XFILLER_6_1008 vgnd vpwr scs8hd_decap_12
XFILLER_1_2354 vpwr vgnd scs8hd_fill_2
XFILLER_1_3099 vgnd vpwr scs8hd_decap_12
XFILLER_8_2508 vgnd vpwr scs8hd_decap_12
XFILLER_7_3990 vgnd vpwr scs8hd_decap_12
XFILLER_6_2276 vgnd vpwr scs8hd_decap_12
XFILLER_6_1520 vgnd vpwr scs8hd_decap_12
XFILLER_2_2118 vgnd vpwr scs8hd_decap_12
XFILLER_0_1141 vgnd vpwr scs8hd_decap_6
XFILLER_8_4411 vgnd vpwr scs8hd_decap_12
XANTENNA__20__A gfpga_pad_GPIO_PAD[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_3765 vgnd vpwr scs8hd_decap_12
XFILLER_7_1306 vgnd vpwr scs8hd_decap_12
XFILLER_4_3618 vgnd vpwr scs8hd_decap_12
XFILLER_1_745 vgnd vpwr scs8hd_decap_12
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XFILLER_2_2630 vgnd vpwr scs8hd_decap_12
XFILLER_2_4021 vgnd vpwr scs8hd_decap_12
XFILLER_5_1074 vgnd vpwr scs8hd_decap_12
XFILLER_2_1984 vgnd vpwr scs8hd_decap_12
XFILLER_8_300 vgnd vpwr scs8hd_decap_12
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_2563 vgnd vpwr scs8hd_decap_12
XFILLER_3_2416 vgnd vpwr scs8hd_decap_12
XFILLER_1_2184 vgnd vpwr scs8hd_decap_12
XFILLER_5_3905 vgnd vpwr scs8hd_decap_12
XFILLER_3_3673 vgnd vpwr scs8hd_decap_12
XFILLER_6_1361 vgnd vpwr scs8hd_decap_12
XFILLER_2_1203 vgnd vpwr scs8hd_decap_12
XFILLER_6_837 vgnd vpwr scs8hd_decap_12
XANTENNA__15__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_4241 vgnd vpwr scs8hd_decap_12
XFILLER_8_2850 vgnd vpwr scs8hd_decap_12
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_7_1147 vgnd vpwr scs8hd_decap_12
XFILLER_4_3448 vgnd vpwr scs8hd_decap_12
XFILLER_4_2703 vgnd vpwr scs8hd_decap_12
XFILLER_1_586 vgnd vpwr scs8hd_decap_12
XFILLER_9_664 vgnd vpwr scs8hd_decap_12
XFILLER_8_141 vgnd vpwr scs8hd_decap_12
XFILLER_9_2636 vgnd vpwr scs8hd_decap_12
XFILLER_4_3960 vgnd vpwr scs8hd_decap_12
XFILLER_0_4558 vgnd vpwr scs8hd_decap_12
XPHY_909 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1501 vgnd vpwr scs8hd_decap_12
XFILLER_0_3857 vgnd vpwr scs8hd_decap_12
XFILLER_3_818 vgnd vpwr scs8hd_decap_12
XFILLER_8_2179 vgnd vpwr scs8hd_decap_12
XFILLER_6_1191 vgnd vpwr scs8hd_decap_12
XFILLER_5_3746 vgnd vpwr scs8hd_decap_12
XFILLER_2_1044 vgnd vpwr scs8hd_decap_12
XFILLER_6_678 vgnd vpwr scs8hd_decap_12
XFILLER_8_4082 vgnd vpwr scs8hd_decap_12
XFILLER_8_2691 vgnd vpwr scs8hd_decap_12
XFILLER_2_873 vgnd vpwr scs8hd_decap_12
XFILLER_4_3289 vgnd vpwr scs8hd_decap_12
XFILLER_4_2533 vgnd vpwr scs8hd_decap_12
XFILLER_4_1898 vgnd vpwr scs8hd_decap_12
XFILLER_0_1718 vgnd vpwr scs8hd_decap_12
XFILLER_0_2419 vgnd vpwr scs8hd_decap_12
XFILLER_9_3156 vgnd vpwr scs8hd_decap_6
XFILLER_9_3101 vgnd vpwr scs8hd_decap_12
XFILLER_9_2400 vgnd vpwr scs8hd_decap_12
XFILLER_5_2319 vgnd vpwr scs8hd_decap_4
Xlogical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _12_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_3621 vgnd vpwr scs8hd_decap_6
XFILLER_0_4322 vgnd vpwr scs8hd_decap_12
XPHY_739 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_728 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_717 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_706 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_2087 vgnd vpwr scs8hd_decap_12
XANTENNA__12__B _11_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_3690 vgnd vpwr scs8hd_decap_12
XFILLER_7_3819 vgnd vpwr scs8hd_decap_12
XFILLER_5_4222 vgnd vpwr scs8hd_decap_12
XFILLER_5_2831 vgnd vpwr scs8hd_decap_12
XFILLER_3_659 vgnd vpwr scs8hd_decap_12
XFILLER_8_1264 vgnd vpwr scs8hd_decap_12
XFILLER_5_3587 vgnd vpwr scs8hd_decap_12
XFILLER_4_1117 vgnd vpwr scs8hd_decap_12
XFILLER_1_3429 vgnd vpwr scs8hd_decap_12
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_965 vgnd vpwr scs8hd_decap_8
XFILLER_6_2606 vgnd vpwr scs8hd_decap_12
XFILLER_1_3941 vgnd vpwr scs8hd_decap_12
XFILLER_9_280 vgnd vpwr scs8hd_decap_12
XFILLER_9_1551 vgnd vpwr scs8hd_decap_12
XFILLER_5_1404 vgnd vpwr scs8hd_decap_12
XFILLER_3_1172 vgnd vpwr scs8hd_decap_12
XFILLER_0_3473 vgnd vpwr scs8hd_decap_12
XFILLER_2_3716 vgnd vpwr scs8hd_decap_12
XPHY_569 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_558 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_547 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_536 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_525 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_514 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_503 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__07__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_2772 vgnd vpwr scs8hd_decap_12
XANTENNA__23__A gfpga_pad_GPIO_PAD[4] vgnd vpwr scs8hd_diode_2
XFILLER_7_2904 vgnd vpwr scs8hd_decap_12
XFILLER_5_4063 vgnd vpwr scs8hd_decap_12
XFILLER_5_2672 vgnd vpwr scs8hd_decap_12
XFILLER_3_489 vgnd vpwr scs8hd_decap_12
XFILLER_1_2514 vgnd vpwr scs8hd_decap_12
XFILLER_1_1879 vgnd vpwr scs8hd_decap_12
XFILLER_6_2447 vgnd vpwr scs8hd_decap_12
XFILLER_0_1389 vgnd vpwr scs8hd_decap_6
XFILLER_0_1334 vgnd vpwr scs8hd_decap_12
XFILLER_9_2071 vgnd vpwr scs8hd_decap_6
XFILLER_8_3936 vgnd vpwr scs8hd_decap_12
XFILLER_6_4350 vgnd vpwr scs8hd_decap_12
XFILLER_1_916 vgnd vpwr scs8hd_decap_12
XFILLER_0_459 vgnd vpwr scs8hd_decap_6
XFILLER_0_404 vgnd vpwr scs8hd_decap_12
XFILLER_2_2801 vgnd vpwr scs8hd_decap_12
XFILLER_2_3557 vgnd vpwr scs8hd_decap_12
XANTENNA__18__A gfpga_pad_GPIO_PAD[7] vgnd vpwr scs8hd_diode_2
XFILLER_5_1245 vgnd vpwr scs8hd_decap_12
XPHY_300 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_399 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_388 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_377 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_366 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_355 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_344 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_333 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_322 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_311 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4136 vgnd vpwr scs8hd_decap_12
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_4_776 vgnd vpwr scs8hd_decap_12
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XFILLER_0_993 vgnd vpwr scs8hd_decap_12
XFILLER_1_2322 vgnd vpwr scs8hd_decap_4
XFILLER_6_1532 vgnd vpwr scs8hd_decap_12
XFILLER_3_3844 vgnd vpwr scs8hd_decap_12
XFILLER_8_3777 vgnd vpwr scs8hd_decap_12
XFILLER_6_4180 vgnd vpwr scs8hd_decap_12
XFILLER_7_1318 vgnd vpwr scs8hd_decap_12
XFILLER_5_1020 vgnd vpwr scs8hd_decap_12
XFILLER_1_757 vgnd vpwr scs8hd_decap_12
XFILLER_2_2642 vgnd vpwr scs8hd_decap_12
XFILLER_2_3387 vgnd vpwr scs8hd_decap_12
XFILLER_2_4033 vgnd vpwr scs8hd_decap_12
XFILLER_5_1086 vgnd vpwr scs8hd_decap_12
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_1996 vgnd vpwr scs8hd_decap_12
XFILLER_8_312 vgnd vpwr scs8hd_decap_12
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3221 vgnd vpwr scs8hd_decap_12
XFILLER_7_2575 vgnd vpwr scs8hd_decap_12
XFILLER_3_2428 vgnd vpwr scs8hd_decap_12
XFILLER_1_1440 vgnd vpwr scs8hd_decap_12
XFILLER_5_3917 vgnd vpwr scs8hd_decap_12
XFILLER_8_1605 vgnd vpwr scs8hd_decap_12
XFILLER_3_3685 vgnd vpwr scs8hd_decap_12
XFILLER_2_1215 vgnd vpwr scs8hd_decap_12
XFILLER_6_849 vgnd vpwr scs8hd_decap_12
XANTENNA__15__B _11_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_4253 vgnd vpwr scs8hd_decap_12
XFILLER_8_2862 vgnd vpwr scs8hd_decap_12
XFILLER_4_4106 vgnd vpwr scs8hd_decap_12
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_598 vgnd vpwr scs8hd_decap_12
XFILLER_2_2472 vgnd vpwr scs8hd_decap_12
XFILLER_9_621 vgnd vpwr scs8hd_decap_12
XFILLER_9_3349 vgnd vpwr scs8hd_decap_12
XFILLER_9_676 vgnd vpwr scs8hd_decap_6
XFILLER_9_2648 vgnd vpwr scs8hd_decap_12
XFILLER_7_3051 vgnd vpwr scs8hd_decap_12
XFILLER_7_1660 vgnd vpwr scs8hd_decap_12
XFILLER_4_3972 vgnd vpwr scs8hd_decap_12
XFILLER_3_2258 vgnd vpwr scs8hd_decap_12
XFILLER_3_1513 vgnd vpwr scs8hd_decap_12
XFILLER_0_3814 vgnd vpwr scs8hd_decap_12
XFILLER_0_3869 vgnd vpwr scs8hd_decap_6
XFILLER_9_4551 vgnd vpwr scs8hd_decap_6
XFILLER_5_3758 vgnd vpwr scs8hd_decap_12
XFILLER_8_1435 vgnd vpwr scs8hd_decap_12
XFILLER_3_4161 vgnd vpwr scs8hd_decap_12
XFILLER_3_2770 vgnd vpwr scs8hd_decap_12
XFILLER_2_1056 vgnd vpwr scs8hd_decap_12
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XFILLER_8_4094 vgnd vpwr scs8hd_decap_12
XFILLER_4_2545 vgnd vpwr scs8hd_decap_12
XFILLER_9_3113 vgnd vpwr scs8hd_decap_12
XFILLER_9_2412 vgnd vpwr scs8hd_decap_6
XFILLER_9_2489 vgnd vpwr scs8hd_decap_12
XFILLER_9_1799 vgnd vpwr scs8hd_decap_12
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_3_2099 vgnd vpwr scs8hd_decap_12
XFILLER_3_1343 vgnd vpwr scs8hd_decap_12
XFILLER_0_4334 vgnd vpwr scs8hd_decap_6
XPHY_729 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_718 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_707 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__12__C _13_/C vgnd vpwr scs8hd_diode_2
XFILLER_8_1276 vgnd vpwr scs8hd_decap_12
XFILLER_5_4234 vgnd vpwr scs8hd_decap_12
XFILLER_5_2843 vgnd vpwr scs8hd_decap_12
XFILLER_9_27 vgnd vpwr scs8hd_decap_4
XFILLER_6_410 vgnd vpwr scs8hd_decap_12
XFILLER_6_4009 vgnd vpwr scs8hd_decap_12
XFILLER_7_977 vgnd vpwr scs8hd_decap_12
XFILLER_6_2618 vgnd vpwr scs8hd_decap_12
XFILLER_4_3021 vgnd vpwr scs8hd_decap_12
XFILLER_4_2320 vpwr vgnd scs8hd_fill_2
XFILLER_4_1630 vgnd vpwr scs8hd_decap_12
XFILLER_1_3953 vgnd vpwr scs8hd_decap_12
XFILLER_9_292 vgnd vpwr scs8hd_decap_12
XFILLER_9_2264 vgnd vpwr scs8hd_decap_12
XFILLER_9_1563 vgnd vpwr scs8hd_decap_12
XFILLER_6_4521 vgnd vpwr scs8hd_decap_12
XFILLER_6_3875 vgnd vpwr scs8hd_decap_12
XFILLER_5_1416 vgnd vpwr scs8hd_decap_12
XFILLER_2_3728 vgnd vpwr scs8hd_decap_12
XANTENNA__07__C _10_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_1184 vgnd vpwr scs8hd_decap_12
XFILLER_0_2784 vgnd vpwr scs8hd_decap_6
XFILLER_0_3485 vgnd vpwr scs8hd_decap_12
XFILLER_0_4186 vgnd vpwr scs8hd_decap_12
XPHY_559 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_548 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_537 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_526 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_515 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_504 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4307 vgnd vpwr scs8hd_decap_12
XFILLER_7_2916 vgnd vpwr scs8hd_decap_12
XFILLER_4_947 vgnd vpwr scs8hd_decap_12
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_4075 vgnd vpwr scs8hd_decap_12
XFILLER_1_2526 vgnd vpwr scs8hd_decap_12
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
XFILLER_6_2459 vgnd vpwr scs8hd_decap_12
XFILLER_6_1703 vgnd vpwr scs8hd_decap_12
XFILLER_4_1471 vgnd vpwr scs8hd_decap_12
XFILLER_0_1346 vgnd vpwr scs8hd_decap_12
XFILLER_0_2047 vgnd vpwr scs8hd_decap_12
XFILLER_1_3783 vgnd vpwr scs8hd_decap_12
XFILLER_8_3948 vgnd vpwr scs8hd_decap_12
XFILLER_6_2960 vgnd vpwr scs8hd_decap_12
XFILLER_5_1257 vgnd vpwr scs8hd_decap_12
XFILLER_1_928 vgnd vpwr scs8hd_decap_12
XFILLER_0_416 vgnd vpwr scs8hd_decap_12
XFILLER_2_2813 vgnd vpwr scs8hd_decap_12
XFILLER_2_4204 vgnd vpwr scs8hd_decap_12
XPHY_334 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_323 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_312 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_301 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_389 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_378 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_367 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_356 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_345 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_2746 vgnd vpwr scs8hd_decap_12
XFILLER_4_788 vgnd vpwr scs8hd_decap_12
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
XFILLER_5_3160 vgnd vpwr scs8hd_decap_12
XFILLER_1_1611 vgnd vpwr scs8hd_decap_12
XFILLER_1_2312 vpwr vgnd scs8hd_fill_2
XFILLER_1_3002 vgnd vpwr scs8hd_decap_12
XPHY_890 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_2289 vgnd vpwr scs8hd_decap_12
XFILLER_6_1544 vgnd vpwr scs8hd_decap_12
XFILLER_3_4502 vgnd vpwr scs8hd_decap_12
XFILLER_3_3856 vgnd vpwr scs8hd_decap_12
XFILLER_0_1110 vgnd vpwr scs8hd_decap_6
XFILLER_8_4424 vgnd vpwr scs8hd_decap_12
XFILLER_8_3789 vgnd vpwr scs8hd_decap_12
XFILLER_6_4192 vgnd vpwr scs8hd_decap_12
XFILLER_1_769 vgnd vpwr scs8hd_decap_12
XFILLER_5_1032 vgnd vpwr scs8hd_decap_4
XFILLER_2_3399 vgnd vpwr scs8hd_decap_12
XFILLER_2_4045 vgnd vpwr scs8hd_decap_12
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_869 vgnd vpwr scs8hd_decap_12
XFILLER_8_324 vgnd vpwr scs8hd_decap_12
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_2587 vgnd vpwr scs8hd_decap_12
XFILLER_7_1831 vgnd vpwr scs8hd_decap_8
XFILLER_1_1452 vgnd vpwr scs8hd_decap_12
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_1_2197 vgnd vpwr scs8hd_decap_12
XFILLER_8_3008 vgnd vpwr scs8hd_decap_12
XFILLER_7_4490 vgnd vpwr scs8hd_decap_12
XFILLER_5_3929 vgnd vpwr scs8hd_decap_12
XFILLER_3_4332 vgnd vpwr scs8hd_decap_12
XFILLER_6_2020 vgnd vpwr scs8hd_decap_12
XFILLER_6_1374 vgnd vpwr scs8hd_decap_12
XFILLER_3_3697 vgnd vpwr scs8hd_decap_12
XFILLER_3_2941 vgnd vpwr scs8hd_decap_12
XFILLER_2_1227 vgnd vpwr scs8hd_decap_12
XANTENNA__15__C _13_/C vgnd vpwr scs8hd_diode_2
XFILLER_8_4265 vgnd vpwr scs8hd_decap_12
XFILLER_8_2874 vgnd vpwr scs8hd_decap_12
XFILLER_4_2716 vgnd vpwr scs8hd_decap_12
XFILLER_2_3130 vgnd vpwr scs8hd_decap_12
XFILLER_2_2484 vgnd vpwr scs8hd_decap_12
XFILLER_9_633 vgnd vpwr scs8hd_decap_12
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XFILLER_9_2605 vgnd vpwr scs8hd_decap_12
XFILLER_9_1904 vgnd vpwr scs8hd_decap_12
XFILLER_7_3063 vgnd vpwr scs8hd_decap_12
XFILLER_7_2351 vgnd vpwr scs8hd_decap_12
XFILLER_7_1672 vgnd vpwr scs8hd_decap_12
XFILLER_4_3984 vgnd vpwr scs8hd_decap_12
XFILLER_0_3826 vgnd vpwr scs8hd_decap_12
XFILLER_0_4527 vgnd vpwr scs8hd_decap_12
XFILLER_1_1282 vgnd vpwr scs8hd_decap_12
XFILLER_8_1447 vgnd vpwr scs8hd_decap_12
XFILLER_5_4405 vgnd vpwr scs8hd_decap_12
XFILLER_3_4173 vgnd vpwr scs8hd_decap_12
XFILLER_3_2782 vgnd vpwr scs8hd_decap_12
XFILLER_8_3350 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
XFILLER_4_2557 vgnd vpwr scs8hd_decap_12
XFILLER_4_1801 vgnd vpwr scs8hd_decap_12
XFILLER_1_330 vgnd vpwr scs8hd_decap_12
XFILLER_2_886 vgnd vpwr scs8hd_decap_12
XFILLER_9_3125 vgnd vpwr scs8hd_decap_6
XFILLER_4_4460 vgnd vpwr scs8hd_decap_12
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_3_2001 vgnd vpwr scs8hd_decap_12
XFILLER_3_1355 vgnd vpwr scs8hd_decap_12
XFILLER_0_2977 vgnd vpwr scs8hd_decap_12
XPHY_719 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_708 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__12__D _10_/D vgnd vpwr scs8hd_diode_2
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XFILLER_8_1288 vgnd vpwr scs8hd_decap_12
XFILLER_5_4246 vgnd vpwr scs8hd_decap_12
XFILLER_5_2855 vgnd vpwr scs8hd_decap_12
XFILLER_6_422 vgnd vpwr scs8hd_decap_12
XFILLER_8_3191 vgnd vpwr scs8hd_decap_12
XFILLER_7_989 vgnd vpwr scs8hd_decap_12
XFILLER_4_3033 vgnd vpwr scs8hd_decap_12
XFILLER_4_2387 vgnd vpwr scs8hd_decap_12
XFILLER_4_2343 vgnd vpwr scs8hd_fill_1
XFILLER_4_1642 vgnd vpwr scs8hd_decap_12
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XFILLER_6_4533 vgnd vpwr scs8hd_decap_12
XFILLER_9_2276 vgnd vpwr scs8hd_decap_12
XFILLER_9_1575 vgnd vpwr scs8hd_decap_6
XFILLER_9_1520 vgnd vpwr scs8hd_decap_12
XFILLER_6_3887 vgnd vpwr scs8hd_decap_12
XFILLER_5_1428 vgnd vpwr scs8hd_decap_12
XPHY_516 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_505 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1196 vgnd vpwr scs8hd_decap_12
XFILLER_0_2741 vgnd vpwr scs8hd_decap_12
XFILLER_0_3442 vgnd vpwr scs8hd_decap_12
XFILLER_0_3497 vgnd vpwr scs8hd_decap_6
XFILLER_0_4198 vgnd vpwr scs8hd_decap_12
XANTENNA__07__D enable vgnd vpwr scs8hd_diode_2
XPHY_549 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
XPHY_538 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_527 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4319 vgnd vpwr scs8hd_decap_12
XFILLER_5_3331 vgnd vpwr scs8hd_decap_12
XFILLER_4_959 vgnd vpwr scs8hd_decap_12
XFILLER_3_403 vgnd vpwr scs8hd_decap_12
XFILLER_5_2685 vgnd vpwr scs8hd_decap_12
XFILLER_5_1940 vgnd vpwr scs8hd_decap_12
XFILLER_1_2538 vgnd vpwr scs8hd_decap_12
XFILLER_7_720 vgnd vpwr scs8hd_decap_12
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_3106 vgnd vpwr scs8hd_decap_12
XFILLER_6_1715 vgnd vpwr scs8hd_decap_12
XFILLER_1_4441 vgnd vpwr scs8hd_decap_12
XFILLER_4_1483 vgnd vpwr scs8hd_decap_12
XFILLER_0_1358 vgnd vpwr scs8hd_decap_6
XFILLER_0_1303 vgnd vpwr scs8hd_decap_12
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_0_2059 vgnd vpwr scs8hd_decap_12
XFILLER_1_3795 vgnd vpwr scs8hd_decap_12
XFILLER_9_2040 vgnd vpwr scs8hd_decap_6
XFILLER_6_4363 vgnd vpwr scs8hd_decap_12
XFILLER_0_428 vgnd vpwr scs8hd_decap_6
XFILLER_2_4216 vgnd vpwr scs8hd_decap_12
XFILLER_6_2972 vgnd vpwr scs8hd_decap_12
XFILLER_5_1269 vgnd vpwr scs8hd_decap_12
XFILLER_2_2825 vgnd vpwr scs8hd_decap_12
XPHY_368 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_357 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_346 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_335 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_324 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_313 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_1892 vgnd vpwr scs8hd_decap_12
XPHY_302 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_379 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4149 vgnd vpwr scs8hd_decap_12
XFILLER_7_3404 vgnd vpwr scs8hd_decap_12
XFILLER_7_2758 vgnd vpwr scs8hd_decap_12
XFILLER_0_962 vgnd vpwr scs8hd_decap_12
XFILLER_1_3014 vgnd vpwr scs8hd_decap_12
XFILLER_5_1770 vgnd vpwr scs8hd_decap_12
XFILLER_1_1623 vgnd vpwr scs8hd_decap_12
XPHY_891 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_880 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_550 vgnd vpwr scs8hd_decap_12
XFILLER_3_3868 vgnd vpwr scs8hd_decap_12
XFILLER_1_4271 vgnd vpwr scs8hd_decap_12
X_09_ address[1] enable address[3] _10_/D _09_/X vgnd vpwr scs8hd_and4_4
XFILLER_1_2880 vgnd vpwr scs8hd_decap_12
XFILLER_8_4436 vgnd vpwr scs8hd_decap_12
XFILLER_2_3301 vgnd vpwr scs8hd_decap_12
XFILLER_9_1191 vgnd vpwr scs8hd_decap_12
XFILLER_5_1099 vgnd vpwr scs8hd_decap_12
XFILLER_2_1910 vgnd vpwr scs8hd_decap_12
XFILLER_2_2655 vgnd vpwr scs8hd_decap_12
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3234 vgnd vpwr scs8hd_decap_12
XFILLER_4_520 vgnd vpwr scs8hd_decap_12
XFILLER_7_2599 vgnd vpwr scs8hd_decap_12
XFILLER_5_2290 vgnd vpwr scs8hd_decap_3
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_8_1618 vgnd vpwr scs8hd_decap_12
XFILLER_6_2032 vgnd vpwr scs8hd_decap_12
XFILLER_7_391 vgnd vpwr scs8hd_decap_12
XFILLER_3_4344 vgnd vpwr scs8hd_decap_12
XFILLER_6_1386 vgnd vpwr scs8hd_decap_12
XFILLER_3_2953 vgnd vpwr scs8hd_decap_12
XFILLER_2_1239 vgnd vpwr scs8hd_decap_12
XANTENNA__15__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_8_4277 vgnd vpwr scs8hd_decap_12
XFILLER_8_3521 vgnd vpwr scs8hd_decap_12
XFILLER_5_306 vgnd vpwr scs8hd_decap_12
XFILLER_4_4119 vgnd vpwr scs8hd_decap_12
XFILLER_1_501 vgnd vpwr scs8hd_decap_12
XFILLER_8_2886 vgnd vpwr scs8hd_decap_12
XFILLER_4_2728 vgnd vpwr scs8hd_decap_12
XFILLER_2_1740 vgnd vpwr scs8hd_decap_12
XFILLER_2_2496 vgnd vpwr scs8hd_decap_12
XFILLER_9_645 vgnd vpwr scs8hd_decap_6
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XFILLER_9_3318 vgnd vpwr scs8hd_decap_12
XFILLER_9_2617 vgnd vpwr scs8hd_decap_12
XFILLER_9_1927 vpwr vgnd scs8hd_fill_2
XFILLER_9_1916 vgnd vpwr scs8hd_decap_6
XFILLER_7_3075 vgnd vpwr scs8hd_decap_12
XFILLER_4_361 vgnd vpwr scs8hd_decap_12
XFILLER_7_2363 vgnd vpwr scs8hd_decap_12
XFILLER_7_1684 vgnd vpwr scs8hd_decap_12
XFILLER_3_1526 vgnd vpwr scs8hd_decap_12
XFILLER_0_3805 vpwr vgnd scs8hd_fill_2
XFILLER_0_3838 vgnd vpwr scs8hd_decap_6
XFILLER_0_4539 vgnd vpwr scs8hd_decap_12
XFILLER_1_1294 vgnd vpwr scs8hd_decap_12
XFILLER_9_4520 vgnd vpwr scs8hd_decap_6
XFILLER_5_4417 vgnd vpwr scs8hd_decap_12
XFILLER_8_1459 vgnd vpwr scs8hd_decap_12
XFILLER_3_4185 vgnd vpwr scs8hd_decap_12
XFILLER_3_2794 vgnd vpwr scs8hd_decap_12
XFILLER_2_1069 vgnd vpwr scs8hd_decap_12
XFILLER_8_3362 vgnd vpwr scs8hd_decap_12
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XFILLER_4_3204 vgnd vpwr scs8hd_decap_12
XFILLER_1_342 vgnd vpwr scs8hd_decap_12
XFILLER_8_1971 vgnd vpwr scs8hd_decap_12
XFILLER_4_2569 vgnd vpwr scs8hd_decap_12
XFILLER_4_1813 vgnd vpwr scs8hd_decap_12
XFILLER_2_898 vgnd vpwr scs8hd_decap_12
XFILLER_2_1581 vgnd vpwr scs8hd_decap_12
XFILLER_9_497 vgnd vpwr scs8hd_decap_12
XFILLER_9_1768 vgnd vpwr scs8hd_decap_12
XFILLER_7_2160 vgnd vpwr scs8hd_decap_12
XFILLER_4_4472 vgnd vpwr scs8hd_decap_12
XFILLER_0_4303 vgnd vpwr scs8hd_decap_6
XPHY_709 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1367 vgnd vpwr scs8hd_decap_12
XFILLER_0_2989 vgnd vpwr scs8hd_decap_12
XFILLER_9_4372 vgnd vpwr scs8hd_decap_12
XFILLER_9_3671 vgnd vpwr scs8hd_decap_12
XFILLER_5_4258 vgnd vpwr scs8hd_decap_12
XFILLER_5_3502 vgnd vpwr scs8hd_decap_12
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XFILLER_9_2970 vgnd vpwr scs8hd_decap_6
XFILLER_3_3270 vgnd vpwr scs8hd_decap_12
XFILLER_1_2709 vgnd vpwr scs8hd_decap_12
XFILLER_7_946 vgnd vpwr scs8hd_fill_1
XFILLER_6_434 vgnd vpwr scs8hd_decap_12
XFILLER_4_3045 vgnd vpwr scs8hd_decap_12
XFILLER_4_2399 vgnd vpwr scs8hd_decap_8
XFILLER_4_1654 vgnd vpwr scs8hd_decap_12
XFILLER_1_3966 vgnd vpwr scs8hd_decap_12
XFILLER_9_261 vgnd vpwr scs8hd_decap_12
XFILLER_9_2233 vgnd vpwr scs8hd_decap_12
XFILLER_9_2288 vgnd vpwr scs8hd_decap_6
XFILLER_9_1532 vgnd vpwr scs8hd_decap_12
XFILLER_6_4578 vgnd vpwr scs8hd_decap_3
XFILLER_6_3899 vgnd vpwr scs8hd_decap_12
XFILLER_0_3454 vgnd vpwr scs8hd_decap_12
XFILLER_0_4155 vgnd vpwr scs8hd_decap_12
XPHY_539 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_528 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_517 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_506 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_2753 vgnd vpwr scs8hd_decap_6
XFILLER_8_1020 vgnd vpwr scs8hd_decap_12
XFILLER_7_2929 vgnd vpwr scs8hd_decap_12
XFILLER_5_4088 vgnd vpwr scs8hd_decap_12
XFILLER_5_3343 vgnd vpwr scs8hd_decap_12
XFILLER_3_415 vgnd vpwr scs8hd_decap_12
XFILLER_5_2697 vgnd vpwr scs8hd_decap_12
XFILLER_6_3118 vgnd vpwr scs8hd_decap_12
XFILLER_6_2406 vgnd vpwr scs8hd_decap_4
XFILLER_6_1727 vgnd vpwr scs8hd_decap_12
XFILLER_4_2130 vgnd vpwr scs8hd_decap_12
XFILLER_0_1315 vgnd vpwr scs8hd_decap_12
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XFILLER_0_2016 vgnd vpwr scs8hd_decap_12
XFILLER_6_4375 vgnd vpwr scs8hd_decap_12
XFILLER_2_4228 vgnd vpwr scs8hd_decap_12
XFILLER_6_2984 vgnd vpwr scs8hd_decap_12
XFILLER_8_507 vgnd vpwr scs8hd_decap_12
XPHY_369 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_358 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_347 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_336 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_325 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_314 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_303 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_3173 vgnd vpwr scs8hd_decap_12
XFILLER_0_974 vgnd vpwr scs8hd_decap_12
XFILLER_1_3026 vgnd vpwr scs8hd_decap_12
XFILLER_5_1782 vgnd vpwr scs8hd_decap_12
XFILLER_1_1635 vgnd vpwr scs8hd_decap_12
XFILLER_1_2358 vpwr vgnd scs8hd_fill_2
XPHY_892 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_881 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_870 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xlogical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ top_width_0_height_0__pin_10_ logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[5] vgnd vpwr scs8hd_ebufn_1
XFILLER_6_2203 vgnd vpwr scs8hd_decap_12
XFILLER_7_562 vgnd vpwr scs8hd_decap_12
XFILLER_3_4515 vgnd vpwr scs8hd_decap_12
XFILLER_6_1557 vgnd vpwr scs8hd_decap_12
XFILLER_1_4283 vgnd vpwr scs8hd_decap_12
X_08_ address[2] _10_/D vgnd vpwr scs8hd_inv_8
XFILLER_1_2892 vgnd vpwr scs8hd_decap_12
XFILLER_8_4448 vgnd vpwr scs8hd_decap_12
XFILLER_6_3460 vgnd vpwr scs8hd_decap_12
XFILLER_2_3313 vgnd vpwr scs8hd_decap_12
XFILLER_2_4058 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ top_width_0_height_0__pin_14_ vgnd vpwr scs8hd_diode_2
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_3070 vgnd vpwr scs8hd_decap_12
XFILLER_2_2667 vgnd vpwr scs8hd_decap_12
XFILLER_9_838 vgnd vpwr scs8hd_decap_12
XFILLER_8_337 vgnd vpwr scs8hd_decap_12
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3246 vgnd vpwr scs8hd_decap_12
XFILLER_4_532 vgnd vpwr scs8hd_decap_12
XFILLER_7_1888 vgnd vpwr scs8hd_decap_3
XFILLER_7_1844 vgnd vpwr scs8hd_decap_12
XFILLER_2_4570 vgnd vpwr scs8hd_decap_8
XFILLER_1_2111 vgnd vpwr scs8hd_decap_12
XFILLER_1_1465 vgnd vpwr scs8hd_decap_12
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_4356 vgnd vpwr scs8hd_decap_12
XFILLER_3_3600 vgnd vpwr scs8hd_decap_12
XFILLER_6_1398 vgnd vpwr scs8hd_decap_12
XFILLER_3_2965 vgnd vpwr scs8hd_decap_12
XFILLER_8_4289 vgnd vpwr scs8hd_decap_12
XFILLER_8_3533 vgnd vpwr scs8hd_decap_12
XFILLER_5_318 vgnd vpwr scs8hd_decap_12
XFILLER_1_513 vgnd vpwr scs8hd_decap_12
XFILLER_2_3143 vgnd vpwr scs8hd_decap_12
XFILLER_9_602 vgnd vpwr scs8hd_decap_12
XFILLER_2_1752 vgnd vpwr scs8hd_decap_12
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
XFILLER_5_830 vgnd vpwr scs8hd_decap_12
XFILLER_9_2629 vgnd vpwr scs8hd_decap_6
XFILLER_7_3087 vgnd vpwr scs8hd_decap_12
XFILLER_7_2375 vgnd vpwr scs8hd_decap_4
XFILLER_4_373 vgnd vpwr scs8hd_decap_12
XFILLER_7_1696 vgnd vpwr scs8hd_decap_12
XFILLER_4_3997 vgnd vpwr scs8hd_decap_12
XFILLER_3_1538 vgnd vpwr scs8hd_decap_12
XFILLER_0_590 vgnd vpwr scs8hd_decap_12
XFILLER_8_2106 vgnd vpwr scs8hd_decap_12
XFILLER_8_690 vgnd vpwr scs8hd_decap_12
XFILLER_5_4429 vgnd vpwr scs8hd_decap_12
XFILLER_3_4197 vgnd vpwr scs8hd_decap_12
XFILLER_3_3441 vgnd vpwr scs8hd_decap_12
XFILLER_6_605 vgnd vpwr scs8hd_decap_12
XFILLER_8_3374 vgnd vpwr scs8hd_decap_12
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
XFILLER_4_3216 vgnd vpwr scs8hd_decap_12
XFILLER_1_354 vgnd vpwr scs8hd_decap_12
XFILLER_2_800 vgnd vpwr scs8hd_decap_12
XFILLER_4_1825 vgnd vpwr scs8hd_decap_12
XFILLER_2_1593 vgnd vpwr scs8hd_decap_12
XFILLER_7_2172 vgnd vpwr scs8hd_decap_12
XFILLER_3_2014 vgnd vpwr scs8hd_decap_12
XFILLER_3_1379 vgnd vpwr scs8hd_decap_12
XFILLER_0_2946 vgnd vpwr scs8hd_decap_12
XFILLER_9_4384 vgnd vpwr scs8hd_decap_12
XFILLER_9_3683 vgnd vpwr scs8hd_decap_6
XFILLER_5_3514 vgnd vpwr scs8hd_decap_12
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XFILLER_5_2868 vgnd vpwr scs8hd_decap_12
XFILLER_3_3282 vgnd vpwr scs8hd_decap_12
XFILLER_7_903 vgnd vpwr scs8hd_decap_12
XFILLER_6_446 vgnd vpwr scs8hd_decap_12
XFILLER_4_3057 vgnd vpwr scs8hd_decap_12
XFILLER_4_2356 vgnd vpwr scs8hd_fill_1
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ top_width_0_height_0__pin_10_ vgnd vpwr scs8hd_diode_2
XFILLER_4_1666 vgnd vpwr scs8hd_decap_12
XFILLER_1_3978 vgnd vpwr scs8hd_decap_12
XFILLER_9_273 vgnd vpwr scs8hd_decap_6
XFILLER_9_2245 vgnd vpwr scs8hd_decap_12
XFILLER_6_4546 vgnd vpwr scs8hd_decap_12
XFILLER_6_3801 vgnd vpwr scs8hd_decap_12
XFILLER_9_1544 vgnd vpwr scs8hd_decap_6
XFILLER_0_2710 vgnd vpwr scs8hd_decap_12
XFILLER_0_3411 vgnd vpwr scs8hd_decap_12
XFILLER_0_3466 vgnd vpwr scs8hd_decap_6
XFILLER_0_4167 vgnd vpwr scs8hd_decap_12
XPHY_529 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_518 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_507 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_1032 vgnd vpwr scs8hd_decap_12
XFILLER_5_1953 vgnd vpwr scs8hd_decap_12
XFILLER_1_1806 vgnd vpwr scs8hd_decap_12
XFILLER_7_733 vgnd vpwr scs8hd_decap_12
XFILLER_6_276 vgnd vpwr scs8hd_decap_12
XFILLER_4_2142 vgnd vpwr scs8hd_decap_12
XFILLER_0_2028 vgnd vpwr scs8hd_decap_12
XFILLER_1_4454 vgnd vpwr scs8hd_decap_12
XFILLER_2_471 vgnd vpwr scs8hd_decap_12
XFILLER_4_1496 vgnd vpwr scs8hd_decap_12
XFILLER_0_1327 vgnd vpwr scs8hd_decap_6
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XFILLER_6_4387 vgnd vpwr scs8hd_decap_12
XFILLER_6_3631 vgnd vpwr scs8hd_decap_12
XFILLER_9_1396 vgnd vpwr scs8hd_decap_12
XFILLER_6_2996 vgnd vpwr scs8hd_decap_12
XFILLER_2_2838 vgnd vpwr scs8hd_decap_12
XPHY_359 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_348 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_337 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_326 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_315 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_1861 vgnd vpwr scs8hd_decap_12
XPHY_304 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3417 vgnd vpwr scs8hd_decap_12
XFILLER_4_703 vgnd vpwr scs8hd_decap_12
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_3185 vgnd vpwr scs8hd_decap_12
XFILLER_0_986 vgnd vpwr scs8hd_decap_6
XFILLER_0_931 vgnd vpwr scs8hd_decap_12
XFILLER_1_2326 vgnd vpwr scs8hd_fill_1
XFILLER_1_3038 vgnd vpwr scs8hd_decap_12
XFILLER_5_1794 vgnd vpwr scs8hd_decap_12
XPHY_893 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_882 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_871 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_860 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_574 vgnd vpwr scs8hd_decap_12
XFILLER_6_2215 vgnd vpwr scs8hd_decap_12
XFILLER_3_4527 vgnd vpwr scs8hd_decap_12
XFILLER_6_1569 vgnd vpwr scs8hd_decap_12
X_07_ _13_/C address[2] _10_/A enable _07_/X vgnd vpwr scs8hd_and4_4
XFILLER_1_4295 vgnd vpwr scs8hd_decap_12
XFILLER_0_1179 vgnd vpwr scs8hd_decap_12
XFILLER_8_3704 vgnd vpwr scs8hd_decap_12
XFILLER_9_1160 vgnd vpwr scs8hd_decap_12
XFILLER_6_3472 vgnd vpwr scs8hd_decap_12
XFILLER_0_249 vgnd vpwr scs8hd_decap_12
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_3082 vgnd vpwr scs8hd_decap_12
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_1923 vgnd vpwr scs8hd_decap_12
XFILLER_2_2679 vgnd vpwr scs8hd_decap_12
XFILLER_8_349 vgnd vpwr scs8hd_decap_12
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3258 vgnd vpwr scs8hd_decap_12
XFILLER_7_2502 vgnd vpwr scs8hd_decap_12
XFILLER_4_544 vgnd vpwr scs8hd_decap_12
XFILLER_7_1856 vgnd vpwr scs8hd_decap_12
XFILLER_3_1709 vgnd vpwr scs8hd_decap_12
XFILLER_1_2123 vgnd vpwr scs8hd_decap_12
XFILLER_1_1477 vgnd vpwr scs8hd_decap_12
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_8_861 vgnd vpwr scs8hd_decap_12
XPHY_690 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XFILLER_7_3770 vgnd vpwr scs8hd_decap_12
XFILLER_6_2045 vgnd vpwr scs8hd_decap_12
XFILLER_6_1300 vgnd vpwr scs8hd_decap_12
XFILLER_3_4368 vgnd vpwr scs8hd_decap_12
XFILLER_3_3612 vgnd vpwr scs8hd_decap_12
XFILLER_3_2977 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ top_width_0_height_0__pin_6_ vgnd vpwr scs8hd_diode_2
XFILLER_1_3380 vgnd vpwr scs8hd_decap_12
XFILLER_8_3545 vgnd vpwr scs8hd_decap_12
XFILLER_1_525 vgnd vpwr scs8hd_decap_12
XFILLER_8_2899 vgnd vpwr scs8hd_decap_12
XFILLER_2_3155 vgnd vpwr scs8hd_decap_12
XFILLER_9_614 vgnd vpwr scs8hd_decap_6
XFILLER_2_1764 vgnd vpwr scs8hd_decap_12
XFILLER_5_842 vgnd vpwr scs8hd_decap_12
XFILLER_7_3099 vgnd vpwr scs8hd_decap_12
XFILLER_4_385 vgnd vpwr scs8hd_decap_12
XFILLER_0_4508 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_3876 vgnd vpwr scs8hd_decap_12
XFILLER_8_2118 vgnd vpwr scs8hd_decap_12
XFILLER_6_1130 vgnd vpwr scs8hd_decap_12
XFILLER_3_3453 vgnd vpwr scs8hd_decap_12
XFILLER_8_4021 vgnd vpwr scs8hd_decap_12
XFILLER_6_617 vgnd vpwr scs8hd_decap_12
XFILLER_8_2630 vgnd vpwr scs8hd_decap_12
XFILLER_4_3228 vgnd vpwr scs8hd_decap_12
XFILLER_2_812 vgnd vpwr scs8hd_decap_12
XFILLER_8_1984 vgnd vpwr scs8hd_decap_12
XFILLER_4_1837 vgnd vpwr scs8hd_decap_12
XFILLER_2_2240 vgnd vpwr scs8hd_decap_12
XFILLER_9_466 vgnd vpwr scs8hd_decap_12
XFILLER_5_672 vgnd vpwr scs8hd_decap_12
XFILLER_9_1737 vgnd vpwr scs8hd_decap_12
XFILLER_7_2184 vgnd vpwr scs8hd_decap_12
XFILLER_4_4485 vgnd vpwr scs8hd_decap_12
XFILLER_4_3740 vgnd vpwr scs8hd_decap_12
XFILLER_3_2026 vgnd vpwr scs8hd_decap_12
XFILLER_0_3659 vgnd vpwr scs8hd_decap_12
XFILLER_0_2958 vgnd vpwr scs8hd_decap_12
XFILLER_9_4341 vgnd vpwr scs8hd_decap_12
XFILLER_9_4396 vgnd vpwr scs8hd_decap_6
XFILLER_9_3640 vgnd vpwr scs8hd_decap_12
XFILLER_8_1203 vgnd vpwr scs8hd_decap_12
XFILLER_5_3526 vgnd vpwr scs8hd_decap_12
XFILLER_3_1892 vgnd vpwr scs8hd_decap_12
XFILLER_2_642 vgnd vpwr scs8hd_decap_12
XFILLER_4_3069 vgnd vpwr scs8hd_decap_12
XFILLER_4_2368 vgnd vpwr scs8hd_decap_12
XFILLER_4_2346 vgnd vpwr scs8hd_decap_3
XFILLER_4_2324 vpwr vgnd scs8hd_fill_2
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XFILLER_2_2081 vgnd vpwr scs8hd_decap_12
XFILLER_9_230 vgnd vpwr scs8hd_decap_12
XFILLER_9_2257 vgnd vpwr scs8hd_decap_6
XFILLER_9_2202 vgnd vpwr scs8hd_decap_12
XFILLER_9_1501 vgnd vpwr scs8hd_decap_12
XFILLER_6_4558 vgnd vpwr scs8hd_decap_12
XFILLER_4_3570 vgnd vpwr scs8hd_decap_12
XFILLER_3_1111 vgnd vpwr scs8hd_decap_12
XFILLER_0_2722 vgnd vpwr scs8hd_decap_6
XFILLER_0_3423 vgnd vpwr scs8hd_decap_12
XFILLER_0_4124 vgnd vpwr scs8hd_decap_12
XFILLER_0_4179 vgnd vpwr scs8hd_decap_6
XPHY_519 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_508 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_4002 vgnd vpwr scs8hd_decap_12
XFILLER_3_428 vgnd vpwr scs8hd_decap_12
XFILLER_9_2791 vgnd vpwr scs8hd_decap_12
XFILLER_8_1044 vgnd vpwr scs8hd_decap_12
XFILLER_5_3356 vgnd vpwr scs8hd_decap_12
XFILLER_5_2611 vgnd vpwr scs8hd_decap_12
XFILLER_1_3209 vgnd vpwr scs8hd_decap_12
XFILLER_5_1965 vgnd vpwr scs8hd_decap_12
XFILLER_1_1818 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ top_width_0_height_0__pin_2_ vgnd vpwr scs8hd_diode_2
XFILLER_7_745 vgnd vpwr scs8hd_decap_12
XFILLER_6_288 vgnd vpwr scs8hd_decap_12
XFILLER_5_4580 vgnd vpwr scs8hd_fill_1
XFILLER_3_940 vgnd vpwr scs8hd_decap_12
XFILLER_2_483 vgnd vpwr scs8hd_decap_12
X_23_ gfpga_pad_GPIO_PAD[4] top_width_0_height_0__pin_9_ vgnd vpwr scs8hd_buf_2
XFILLER_4_2154 vgnd vpwr scs8hd_decap_12
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
XFILLER_1_4466 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _12_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_4399 vgnd vpwr scs8hd_decap_12
XFILLER_6_3643 vgnd vpwr scs8hd_decap_12
XPHY_316 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_1873 vgnd vpwr scs8hd_decap_12
XFILLER_0_2574 vgnd vpwr scs8hd_decap_12
XPHY_305 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_349 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_338 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_327 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3429 vgnd vpwr scs8hd_decap_12
XFILLER_4_715 vgnd vpwr scs8hd_decap_12
XFILLER_3_269 vgnd vpwr scs8hd_decap_12
XFILLER_5_3197 vgnd vpwr scs8hd_decap_12
XFILLER_5_2441 vgnd vpwr scs8hd_decap_12
XFILLER_0_943 vgnd vpwr scs8hd_decap_12
XFILLER_1_2316 vpwr vgnd scs8hd_fill_2
XPHY_872 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_861 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_850 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_1648 vgnd vpwr scs8hd_decap_12
XPHY_894 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_883 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_586 vgnd vpwr scs8hd_decap_12
XFILLER_7_3941 vgnd vpwr scs8hd_decap_12
XFILLER_3_4539 vgnd vpwr scs8hd_decap_12
XFILLER_3_781 vgnd vpwr scs8hd_decap_12
X_06_ address[1] _10_/A vgnd vpwr scs8hd_inv_8
XFILLER_1_3551 vgnd vpwr scs8hd_decap_12
XFILLER_8_3716 vgnd vpwr scs8hd_decap_12
XFILLER_9_1172 vgnd vpwr scs8hd_decap_6
XFILLER_6_3484 vgnd vpwr scs8hd_decap_12
XFILLER_5_1036 vgnd vpwr scs8hd_fill_1
XFILLER_2_1935 vgnd vpwr scs8hd_decap_12
XFILLER_2_3326 vgnd vpwr scs8hd_decap_12
XFILLER_9_807 vgnd vpwr scs8hd_decap_12
XFILLER_0_2382 vgnd vpwr scs8hd_decap_3
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_3094 vgnd vpwr scs8hd_decap_6
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_2514 vgnd vpwr scs8hd_decap_12
XFILLER_4_556 vgnd vpwr scs8hd_decap_12
XFILLER_7_1868 vgnd vpwr scs8hd_decap_12
XPHY_691 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_680 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_1489 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_8_873 vgnd vpwr scs8hd_decap_12
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XFILLER_6_2057 vgnd vpwr scs8hd_decap_12
XFILLER_3_3624 vgnd vpwr scs8hd_decap_12
XFILLER_1_3392 vgnd vpwr scs8hd_decap_12
XFILLER_8_3557 vgnd vpwr scs8hd_decap_12
XFILLER_8_2801 vgnd vpwr scs8hd_decap_12
XFILLER_1_537 vgnd vpwr scs8hd_decap_12
XFILLER_2_1776 vgnd vpwr scs8hd_decap_12
XFILLER_2_2411 vgnd vpwr scs8hd_decap_12
XFILLER_2_3167 vgnd vpwr scs8hd_decap_12
XFILLER_4_3911 vgnd vpwr scs8hd_decap_12
XFILLER_9_4578 vgnd vpwr scs8hd_decap_3
XFILLER_9_3888 vgnd vpwr scs8hd_decap_12
XFILLER_3_4100 vgnd vpwr scs8hd_decap_12
XFILLER_6_1142 vgnd vpwr scs8hd_decap_12
XFILLER_3_3465 vgnd vpwr scs8hd_decap_12
XFILLER_8_4033 vgnd vpwr scs8hd_decap_12
XFILLER_6_629 vgnd vpwr scs8hd_decap_12
XFILLER_8_3387 vgnd vpwr scs8hd_decap_12
XFILLER_8_2642 vgnd vpwr scs8hd_decap_12
XFILLER_8_1996 vgnd vpwr scs8hd_decap_12
XFILLER_1_367 vgnd vpwr scs8hd_decap_12
XFILLER_4_1849 vgnd vpwr scs8hd_decap_12
XFILLER_2_2252 vgnd vpwr scs8hd_decap_12
XFILLER_9_478 vgnd vpwr scs8hd_decap_12
XFILLER_9_1749 vgnd vpwr scs8hd_decap_12
XFILLER_5_684 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_7_1440 vgnd vpwr scs8hd_decap_12
XFILLER_4_4497 vgnd vpwr scs8hd_decap_12
XFILLER_3_2038 vgnd vpwr scs8hd_decap_12
XFILLER_0_2915 vgnd vpwr scs8hd_decap_12
XFILLER_1_1050 vgnd vpwr scs8hd_decap_12
XFILLER_9_4353 vgnd vpwr scs8hd_decap_12
XFILLER_9_3652 vgnd vpwr scs8hd_decap_6
XFILLER_8_1215 vgnd vpwr scs8hd_decap_12
XFILLER_3_3295 vgnd vpwr scs8hd_decap_12
XFILLER_3_2550 vgnd vpwr scs8hd_decap_12
XFILLER_7_949 vpwr vgnd scs8hd_fill_2
XFILLER_7_916 vgnd vpwr scs8hd_decap_12
XFILLER_6_459 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_654 vgnd vpwr scs8hd_decap_12
XFILLER_8_2472 vgnd vpwr scs8hd_decap_12
XFILLER_4_2303 vgnd vpwr scs8hd_decap_8
XFILLER_4_1679 vgnd vpwr scs8hd_decap_12
XFILLER_2_2093 vgnd vpwr scs8hd_decap_12
XFILLER_9_242 vgnd vpwr scs8hd_decap_6
XFILLER_6_971 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _05_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_2214 vgnd vpwr scs8hd_decap_12
XFILLER_9_1513 vgnd vpwr scs8hd_decap_6
XFILLER_6_3814 vgnd vpwr scs8hd_decap_12
XFILLER_0_4136 vgnd vpwr scs8hd_decap_12
XFILLER_4_3582 vgnd vpwr scs8hd_decap_12
XFILLER_3_1123 vgnd vpwr scs8hd_decap_12
XFILLER_0_3435 vgnd vpwr scs8hd_decap_6
XPHY_509 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_4014 vgnd vpwr scs8hd_decap_12
XFILLER_8_1056 vgnd vpwr scs8hd_decap_12
XFILLER_5_3368 vgnd vpwr scs8hd_decap_12
XFILLER_5_1977 vgnd vpwr scs8hd_decap_12
XFILLER_3_2380 vgnd vpwr scs8hd_decap_12
XFILLER_7_757 vgnd vpwr scs8hd_decap_12
XFILLER_5_3880 vgnd vpwr scs8hd_decap_12
XFILLER_3_952 vgnd vpwr scs8hd_decap_12
XFILLER_2_495 vgnd vpwr scs8hd_decap_12
XFILLER_4_1410 vgnd vpwr scs8hd_decap_12
XFILLER_1_3722 vgnd vpwr scs8hd_decap_12
X_22_ gfpga_pad_GPIO_PAD[3] top_width_0_height_0__pin_7_ vgnd vpwr scs8hd_buf_2
XFILLER_1_4478 vgnd vpwr scs8hd_decap_12
XFILLER_9_1365 vgnd vpwr scs8hd_decap_12
XFILLER_6_3655 vgnd vpwr scs8hd_decap_12
XPHY_339 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_328 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_317 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_1830 vgnd vpwr scs8hd_decap_12
XFILLER_0_1885 vgnd vpwr scs8hd_decap_6
XFILLER_0_2586 vgnd vpwr scs8hd_decap_12
XFILLER_0_3287 vgnd vpwr scs8hd_decap_12
XPHY_306 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_2420 vgnd vpwr scs8hd_fill_1
XFILLER_4_727 vgnd vpwr scs8hd_decap_12
XFILLER_0_955 vgnd vpwr scs8hd_decap_6
XFILLER_0_900 vgnd vpwr scs8hd_decap_12
XFILLER_5_2453 vgnd vpwr scs8hd_decap_12
XFILLER_5_2431 vgnd vpwr scs8hd_decap_8
XPHY_895 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_884 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_873 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_862 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_851 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_840 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_598 vgnd vpwr scs8hd_decap_12
XFILLER_7_3953 vgnd vpwr scs8hd_decap_12
XFILLER_6_2228 vgnd vpwr scs8hd_decap_12
XFILLER_0_1148 vgnd vpwr scs8hd_decap_12
XFILLER_1_3563 vgnd vpwr scs8hd_decap_12
X_05_ _13_/C address[2] address[1] enable _05_/X vgnd vpwr scs8hd_and4_4
XFILLER_8_3728 vgnd vpwr scs8hd_decap_12
XFILLER_6_4131 vgnd vpwr scs8hd_decap_12
XFILLER_1_708 vgnd vpwr scs8hd_decap_12
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XFILLER_6_3496 vgnd vpwr scs8hd_decap_12
XFILLER_6_2740 vgnd vpwr scs8hd_decap_12
XFILLER_5_1004 vpwr vgnd scs8hd_fill_2
XFILLER_0_3051 vgnd vpwr scs8hd_decap_12
XFILLER_2_1947 vgnd vpwr scs8hd_decap_12
XFILLER_2_3338 vgnd vpwr scs8hd_decap_12
XFILLER_9_819 vgnd vpwr scs8hd_decap_12
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_568 vgnd vpwr scs8hd_decap_12
XFILLER_7_2526 vgnd vpwr scs8hd_decap_12
XFILLER_2_3850 vgnd vpwr scs8hd_decap_12
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_1_2136 vgnd vpwr scs8hd_decap_12
XPHY_692 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_681 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_670 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
XFILLER_7_3783 vgnd vpwr scs8hd_decap_12
XFILLER_6_2069 vgnd vpwr scs8hd_decap_12
XFILLER_6_1313 vgnd vpwr scs8hd_decap_12
XFILLER_3_3636 vgnd vpwr scs8hd_decap_12
XFILLER_4_1081 vgnd vpwr scs8hd_decap_12
XFILLER_8_4204 vgnd vpwr scs8hd_decap_12
XFILLER_8_2813 vgnd vpwr scs8hd_decap_12
XFILLER_6_2581 vgnd vpwr scs8hd_decap_12
XFILLER_2_1788 vgnd vpwr scs8hd_decap_12
XFILLER_2_2423 vgnd vpwr scs8hd_decap_12
XFILLER_2_3179 vgnd vpwr scs8hd_decap_12
XFILLER_7_3002 vgnd vpwr scs8hd_decap_12
XFILLER_5_855 vgnd vpwr scs8hd_decap_12
XFILLER_4_398 vgnd vpwr scs8hd_decap_12
XFILLER_7_1611 vgnd vpwr scs8hd_decap_12
XFILLER_4_3923 vgnd vpwr scs8hd_decap_12
XFILLER_3_2209 vgnd vpwr scs8hd_decap_12
XFILLER_0_571 vgnd vpwr scs8hd_decap_12
XFILLER_0_3809 vgnd vpwr scs8hd_decap_4
XFILLER_1_1221 vgnd vpwr scs8hd_decap_12
XFILLER_9_3845 vgnd vpwr scs8hd_decap_12
XFILLER_5_3709 vgnd vpwr scs8hd_decap_12
XFILLER_3_4112 vgnd vpwr scs8hd_decap_12
XFILLER_6_1154 vgnd vpwr scs8hd_decap_12
XFILLER_3_2721 vgnd vpwr scs8hd_decap_12
XFILLER_8_4045 vgnd vpwr scs8hd_decap_12
XFILLER_2_825 vgnd vpwr scs8hd_decap_12
XFILLER_8_3399 vgnd vpwr scs8hd_decap_12
XFILLER_1_379 vgnd vpwr scs8hd_decap_12
XFILLER_2_2264 vgnd vpwr scs8hd_decap_12
XFILLER_9_435 vgnd vpwr scs8hd_decap_12
XFILLER_9_1706 vgnd vpwr scs8hd_decap_12
XFILLER_5_696 vgnd vpwr scs8hd_decap_12
XFILLER_4_3753 vgnd vpwr scs8hd_decap_12
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XFILLER_7_2197 vgnd vpwr scs8hd_decap_12
XFILLER_7_1452 vgnd vpwr scs8hd_decap_12
XFILLER_1_891 vgnd vpwr scs8hd_decap_12
XFILLER_0_2927 vgnd vpwr scs8hd_decap_12
XFILLER_0_3628 vgnd vpwr scs8hd_decap_12
XFILLER_1_1062 vgnd vpwr scs8hd_decap_12
XFILLER_9_4365 vgnd vpwr scs8hd_decap_6
XFILLER_9_4310 vgnd vpwr scs8hd_decap_12
XFILLER_8_1227 vgnd vpwr scs8hd_decap_12
XFILLER_5_3539 vgnd vpwr scs8hd_decap_12
XFILLER_7_928 vgnd vpwr scs8hd_decap_12
XFILLER_8_3130 vgnd vpwr scs8hd_decap_12
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XFILLER_2_666 vgnd vpwr scs8hd_decap_12
XFILLER_8_2484 vgnd vpwr scs8hd_decap_12
XFILLER_9_2226 vgnd vpwr scs8hd_decap_6
XFILLER_6_983 vgnd vpwr scs8hd_decap_12
XFILLER_6_3826 vgnd vpwr scs8hd_decap_12
XFILLER_4_3594 vgnd vpwr scs8hd_decap_12
XFILLER_0_4148 vgnd vpwr scs8hd_decap_6
XFILLER_7_1282 vgnd vpwr scs8hd_decap_12
XFILLER_3_1135 vgnd vpwr scs8hd_decap_12
XFILLER_9_2760 vgnd vpwr scs8hd_decap_12
XFILLER_5_2624 vgnd vpwr scs8hd_decap_12
XFILLER_5_1989 vgnd vpwr scs8hd_decap_12
XFILLER_3_2392 vgnd vpwr scs8hd_decap_12
XFILLER_0_3981 vgnd vpwr scs8hd_decap_12
XFILLER_7_769 vgnd vpwr scs8hd_decap_12
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
XFILLER_5_3892 vgnd vpwr scs8hd_decap_12
XFILLER_3_964 vgnd vpwr scs8hd_decap_12
X_21_ gfpga_pad_GPIO_PAD[2] top_width_0_height_0__pin_5_ vgnd vpwr scs8hd_buf_2
XFILLER_1_3734 vgnd vpwr scs8hd_decap_12
XFILLER_4_2167 vgnd vpwr scs8hd_decap_12
XFILLER_4_1422 vgnd vpwr scs8hd_decap_12
XFILLER_0_2009 vgnd vpwr scs8hd_decap_6
XFILLER_6_4302 vgnd vpwr scs8hd_decap_12
XFILLER_6_2911 vgnd vpwr scs8hd_decap_12
XFILLER_9_2078 vgnd vpwr scs8hd_decap_12
XFILLER_9_1377 vgnd vpwr scs8hd_decap_12
XFILLER_6_3667 vgnd vpwr scs8hd_decap_12
XFILLER_5_1208 vgnd vpwr scs8hd_decap_12
XFILLER_4_4070 vgnd vpwr scs8hd_decap_12
XFILLER_0_2543 vgnd vpwr scs8hd_decap_12
XFILLER_2_3509 vgnd vpwr scs8hd_decap_12
XPHY_329 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_318 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_1842 vgnd vpwr scs8hd_decap_12
XFILLER_0_2598 vgnd vpwr scs8hd_decap_6
XFILLER_0_3299 vgnd vpwr scs8hd_decap_12
XPHY_307 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_739 vgnd vpwr scs8hd_decap_12
XFILLER_9_3280 vgnd vpwr scs8hd_decap_6
XFILLER_0_912 vgnd vpwr scs8hd_decap_12
XFILLER_5_2465 vgnd vpwr scs8hd_decap_12
XFILLER_1_2329 vpwr vgnd scs8hd_fill_2
XPHY_896 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_885 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_874 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_863 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_852 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_841 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_830 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xlogical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _13_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_1252 vgnd vpwr scs8hd_decap_12
XFILLER_3_3807 vgnd vpwr scs8hd_decap_12
XFILLER_3_794 vgnd vpwr scs8hd_decap_12
X_04_ address[3] _13_/C vgnd vpwr scs8hd_buf_1
XFILLER_1_3575 vgnd vpwr scs8hd_decap_12
XFILLER_1_4210 vgnd vpwr scs8hd_decap_12
XFILLER_9_1141 vgnd vpwr scs8hd_decap_6
XFILLER_6_4143 vgnd vpwr scs8hd_decap_12
XFILLER_6_2752 vgnd vpwr scs8hd_decap_12
XFILLER_5_1038 vgnd vpwr scs8hd_decap_12
XFILLER_0_3063 vgnd vpwr scs8hd_decap_6
XFILLER_2_1959 vgnd vpwr scs8hd_decap_12
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_2538 vgnd vpwr scs8hd_decap_12
XFILLER_5_1550 vgnd vpwr scs8hd_decap_12
XFILLER_2_3862 vgnd vpwr scs8hd_decap_12
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_1_2148 vgnd vpwr scs8hd_decap_12
XFILLER_8_886 vgnd vpwr scs8hd_decap_12
XPHY_693 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_682 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_671 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_660 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_330 vgnd vpwr scs8hd_decap_12
XFILLER_7_4441 vgnd vpwr scs8hd_decap_12
XFILLER_7_3795 vgnd vpwr scs8hd_decap_12
XFILLER_6_1325 vgnd vpwr scs8hd_decap_12
XFILLER_4_1093 vgnd vpwr scs8hd_decap_12
XFILLER_3_3648 vgnd vpwr scs8hd_decap_12
XFILLER_1_2660 vgnd vpwr scs8hd_decap_12
XFILLER_1_4051 vgnd vpwr scs8hd_decap_12
XFILLER_8_4216 vgnd vpwr scs8hd_decap_12
XFILLER_8_2825 vgnd vpwr scs8hd_decap_12
XFILLER_2_2435 vgnd vpwr scs8hd_decap_12
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_4_300 vgnd vpwr scs8hd_decap_12
XFILLER_7_3014 vgnd vpwr scs8hd_decap_12
XFILLER_5_867 vgnd vpwr scs8hd_decap_12
XFILLER_7_1623 vgnd vpwr scs8hd_decap_12
XFILLER_5_1391 vgnd vpwr scs8hd_decap_12
XFILLER_1_1233 vgnd vpwr scs8hd_decap_12
XFILLER_0_583 vgnd vpwr scs8hd_decap_6
XFILLER_2_3692 vgnd vpwr scs8hd_decap_12
XFILLER_9_4558 vgnd vpwr scs8hd_decap_12
XFILLER_9_3857 vgnd vpwr scs8hd_decap_12
XFILLER_7_171 vgnd vpwr scs8hd_decap_12
XPHY_490 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4271 vgnd vpwr scs8hd_decap_12
XFILLER_7_2880 vgnd vpwr scs8hd_decap_12
XFILLER_3_4124 vgnd vpwr scs8hd_decap_12
XFILLER_3_3478 vgnd vpwr scs8hd_decap_12
XFILLER_3_2733 vgnd vpwr scs8hd_decap_12
XFILLER_6_1166 vgnd vpwr scs8hd_decap_12
XFILLER_2_1008 vgnd vpwr scs8hd_decap_12
XFILLER_8_3301 vgnd vpwr scs8hd_decap_12
XFILLER_8_2655 vgnd vpwr scs8hd_decap_12
XFILLER_8_1910 vgnd vpwr scs8hd_decap_12
XFILLER_2_837 vgnd vpwr scs8hd_decap_12
XFILLER_4_2508 vgnd vpwr scs8hd_decap_12
XFILLER_3_3990 vgnd vpwr scs8hd_decap_12
XFILLER_2_1520 vgnd vpwr scs8hd_decap_12
XFILLER_2_2276 vgnd vpwr scs8hd_decap_12
XFILLER_9_447 vgnd vpwr scs8hd_decap_12
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XFILLER_9_2419 vgnd vpwr scs8hd_decap_12
XFILLER_9_1718 vgnd vpwr scs8hd_decap_12
XFILLER_4_4411 vgnd vpwr scs8hd_decap_12
XFILLER_4_3765 vgnd vpwr scs8hd_decap_12
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ top_width_0_height_0__pin_12_ logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[6] vgnd vpwr scs8hd_ebufn_1
XFILLER_3_1306 vgnd vpwr scs8hd_decap_12
XFILLER_1_1074 vgnd vpwr scs8hd_decap_12
XFILLER_0_2939 vgnd vpwr scs8hd_decap_6
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_4322 vgnd vpwr scs8hd_decap_12
XFILLER_9_3621 vgnd vpwr scs8hd_decap_6
XFILLER_8_1239 vgnd vpwr scs8hd_decap_12
XFILLER_3_2563 vgnd vpwr scs8hd_decap_12
XFILLER_8_2496 vgnd vpwr scs8hd_decap_12
XFILLER_8_1740 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_3905 vgnd vpwr scs8hd_decap_12
XFILLER_2_678 vgnd vpwr scs8hd_decap_12
XFILLER_2_1361 vgnd vpwr scs8hd_decap_12
XFILLER_9_211 vgnd vpwr scs8hd_decap_6
XFILLER_6_3838 vgnd vpwr scs8hd_decap_12
XFILLER_6_995 vgnd vpwr scs8hd_decap_12
XFILLER_7_1294 vgnd vpwr scs8hd_decap_12
XFILLER_4_4241 vgnd vpwr scs8hd_decap_12
XFILLER_4_2850 vgnd vpwr scs8hd_decap_12
XFILLER_0_3404 vgnd vpwr scs8hd_decap_6
XFILLER_0_4105 vgnd vpwr scs8hd_decap_12
XFILLER_3_1147 vgnd vpwr scs8hd_decap_12
XFILLER_9_3473 vgnd vpwr scs8hd_decap_12
XFILLER_9_2772 vgnd vpwr scs8hd_decap_12
XFILLER_8_1003 vgnd vpwr scs8hd_decap_4
XFILLER_5_4027 vgnd vpwr scs8hd_decap_12
XFILLER_5_2636 vgnd vpwr scs8hd_decap_12
XFILLER_8_1069 vgnd vpwr scs8hd_decap_12
XFILLER_0_3993 vgnd vpwr scs8hd_decap_6
X_20_ gfpga_pad_GPIO_PAD[1] top_width_0_height_0__pin_3_ vgnd vpwr scs8hd_buf_2
XFILLER_8_1581 vgnd vpwr scs8hd_decap_12
XFILLER_4_2179 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_3746 vgnd vpwr scs8hd_decap_12
XFILLER_2_1191 vgnd vpwr scs8hd_decap_12
XFILLER_9_1334 vgnd vpwr scs8hd_decap_12
XFILLER_6_4314 vgnd vpwr scs8hd_decap_12
XFILLER_6_3679 vgnd vpwr scs8hd_decap_12
XFILLER_6_2923 vgnd vpwr scs8hd_decap_12
XFILLER_4_4082 vgnd vpwr scs8hd_decap_12
XFILLER_9_1389 vgnd vpwr scs8hd_decap_6
XFILLER_4_2691 vgnd vpwr scs8hd_decap_12
XFILLER_0_2555 vgnd vpwr scs8hd_decap_12
XFILLER_0_3256 vgnd vpwr scs8hd_decap_12
XPHY_319 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_1854 vgnd vpwr scs8hd_decap_6
XPHY_308 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_2709 vgnd vpwr scs8hd_decap_12
XFILLER_5_3112 vgnd vpwr scs8hd_decap_12
XFILLER_5_2477 vgnd vpwr scs8hd_decap_12
XFILLER_5_1721 vgnd vpwr scs8hd_decap_12
XFILLER_0_924 vgnd vpwr scs8hd_decap_6
XFILLER_1_2308 vpwr vgnd scs8hd_fill_2
XPHY_820 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_897 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_886 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_875 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_864 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_853 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_842 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_831 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_501 vgnd vpwr scs8hd_decap_12
XFILLER_7_3966 vgnd vpwr scs8hd_decap_12
XFILLER_5_4380 vgnd vpwr scs8hd_decap_12
XFILLER_3_3819 vgnd vpwr scs8hd_decap_12
XFILLER_4_1264 vgnd vpwr scs8hd_decap_12
XFILLER_0_1117 vgnd vpwr scs8hd_decap_12
XFILLER_1_2831 vgnd vpwr scs8hd_decap_12
XFILLER_1_3587 vgnd vpwr scs8hd_decap_12
XFILLER_1_4222 vgnd vpwr scs8hd_decap_12
XFILLER_6_4155 vgnd vpwr scs8hd_decap_12
XFILLER_6_2764 vgnd vpwr scs8hd_decap_12
XFILLER_0_3020 vgnd vpwr scs8hd_decap_12
XFILLER_2_2606 vgnd vpwr scs8hd_decap_12
XFILLER_0_2352 vpwr vgnd scs8hd_fill_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_1562 vgnd vpwr scs8hd_decap_12
XFILLER_1_1404 vgnd vpwr scs8hd_decap_12
XFILLER_0_776 vgnd vpwr scs8hd_decap_12
XPHY_661 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_650 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_8_898 vgnd vpwr scs8hd_decap_12
XPHY_694 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_683 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_672 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_342 vgnd vpwr scs8hd_decap_12
XFILLER_6_1337 vgnd vpwr scs8hd_decap_12
XFILLER_3_2904 vgnd vpwr scs8hd_decap_12
XFILLER_1_4063 vgnd vpwr scs8hd_decap_12
XFILLER_1_2672 vgnd vpwr scs8hd_decap_12
XFILLER_8_4228 vgnd vpwr scs8hd_decap_12
XFILLER_6_3240 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _05_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_2594 vgnd vpwr scs8hd_decap_12
XFILLER_2_2447 vgnd vpwr scs8hd_decap_12
XFILLER_0_1470 vgnd vpwr scs8hd_decap_12
XFILLER_0_2171 vgnd vpwr scs8hd_decap_12
XFILLER_8_117 vgnd vpwr scs8hd_decap_12
XFILLER_4_312 vgnd vpwr scs8hd_decap_12
XFILLER_7_3026 vgnd vpwr scs8hd_decap_12
XFILLER_7_1635 vgnd vpwr scs8hd_decap_12
XFILLER_5_879 vgnd vpwr scs8hd_decap_12
XFILLER_4_3936 vgnd vpwr scs8hd_decap_12
XFILLER_2_4350 vgnd vpwr scs8hd_decap_12
XFILLER_0_540 vgnd vpwr scs8hd_decap_12
XFILLER_1_1245 vgnd vpwr scs8hd_decap_12
XPHY_491 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_480 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3869 vgnd vpwr scs8hd_decap_6
XFILLER_9_3814 vgnd vpwr scs8hd_decap_12
XFILLER_7_4283 vgnd vpwr scs8hd_decap_12
XFILLER_7_2892 vgnd vpwr scs8hd_decap_12
XFILLER_6_1178 vgnd vpwr scs8hd_decap_12
XFILLER_3_4136 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_4058 vgnd vpwr scs8hd_decap_12
XFILLER_8_3313 vgnd vpwr scs8hd_decap_12
XFILLER_8_2667 vgnd vpwr scs8hd_decap_12
XFILLER_2_849 vgnd vpwr scs8hd_decap_12
XFILLER_2_1532 vgnd vpwr scs8hd_decap_12
XFILLER_2_2299 vpwr vgnd scs8hd_fill_2
XFILLER_9_459 vgnd vpwr scs8hd_decap_6
XFILLER_9_404 vgnd vpwr scs8hd_decap_12
XFILLER_8_4570 vgnd vpwr scs8hd_decap_8
XFILLER_7_2111 vgnd vpwr scs8hd_decap_12
XFILLER_7_1465 vgnd vpwr scs8hd_decap_12
XFILLER_4_3777 vgnd vpwr scs8hd_decap_12
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XFILLER_3_1318 vgnd vpwr scs8hd_decap_12
XFILLER_2_4180 vgnd vpwr scs8hd_decap_12
XFILLER_1_1086 vgnd vpwr scs8hd_decap_12
XFILLER_9_4334 vgnd vpwr scs8hd_decap_6
XFILLER_9_993 vgnd vpwr scs8hd_decap_3
XFILLER_5_2807 vgnd vpwr scs8hd_decap_12
XFILLER_3_3221 vgnd vpwr scs8hd_decap_12
XFILLER_3_2575 vgnd vpwr scs8hd_decap_12
XFILLER_8_3143 vgnd vpwr scs8hd_decap_12
XFILLER_8_1752 vgnd vpwr scs8hd_decap_12
XFILLER_4_2339 vgnd vpwr scs8hd_decap_4
XFILLER_4_1605 vgnd vpwr scs8hd_decap_12
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_3917 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_440 vgnd vpwr scs8hd_decap_12
XFILLER_4_4253 vgnd vpwr scs8hd_decap_12
XFILLER_4_2862 vgnd vpwr scs8hd_decap_12
XFILLER_0_4117 vgnd vpwr scs8hd_decap_6
XFILLER_9_4186 vgnd vpwr scs8hd_decap_12
XFILLER_9_3485 vgnd vpwr scs8hd_decap_12
XFILLER_9_2784 vgnd vpwr scs8hd_decap_6
XFILLER_5_4039 vgnd vpwr scs8hd_decap_12
XFILLER_5_2648 vgnd vpwr scs8hd_decap_12
XFILLER_3_3051 vgnd vpwr scs8hd_decap_12
XFILLER_3_1660 vgnd vpwr scs8hd_decap_12
XFILLER_0_3950 vgnd vpwr scs8hd_decap_12
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_4551 vgnd vpwr scs8hd_decap_12
XFILLER_3_977 vgnd vpwr scs8hd_decap_12
XFILLER_2_410 vgnd vpwr scs8hd_decap_12
XFILLER_8_1593 vgnd vpwr scs8hd_decap_12
XFILLER_4_1435 vgnd vpwr scs8hd_decap_12
XFILLER_1_3758 vgnd vpwr scs8hd_decap_12
XFILLER_9_2047 vgnd vpwr scs8hd_decap_12
XFILLER_9_1346 vgnd vpwr scs8hd_decap_12
XFILLER_6_4326 vgnd vpwr scs8hd_decap_12
XFILLER_6_2935 vgnd vpwr scs8hd_decap_12
XFILLER_5_281 vgnd vpwr scs8hd_decap_12
XFILLER_4_4094 vgnd vpwr scs8hd_decap_12
XFILLER_0_1811 vgnd vpwr scs8hd_decap_12
XFILLER_0_2512 vgnd vpwr scs8hd_decap_12
XFILLER_0_2567 vgnd vpwr scs8hd_decap_6
XFILLER_0_3268 vgnd vpwr scs8hd_decap_12
XPHY_309 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_3124 vgnd vpwr scs8hd_decap_12
XFILLER_5_2489 vgnd vpwr scs8hd_decap_12
XFILLER_5_1733 vgnd vpwr scs8hd_decap_12
XPHY_854 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_843 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_832 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_821 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_810 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_898 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_887 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_876 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_865 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_513 vgnd vpwr scs8hd_decap_12
XFILLER_7_3978 vgnd vpwr scs8hd_decap_12
XFILLER_6_1508 vgnd vpwr scs8hd_decap_12
XFILLER_1_4234 vgnd vpwr scs8hd_decap_12
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_2990 vgnd vpwr scs8hd_decap_12
XFILLER_4_1276 vgnd vpwr scs8hd_decap_12
XFILLER_0_1129 vgnd vpwr scs8hd_decap_12
XFILLER_1_2843 vgnd vpwr scs8hd_decap_12
XFILLER_6_4167 vgnd vpwr scs8hd_decap_12
XFILLER_6_3411 vgnd vpwr scs8hd_decap_12
XFILLER_9_1110 vgnd vpwr scs8hd_decap_6
XFILLER_0_3032 vgnd vpwr scs8hd_decap_6
XFILLER_2_2618 vgnd vpwr scs8hd_decap_12
XFILLER_2_4009 vgnd vpwr scs8hd_decap_12
XFILLER_0_2375 vgnd vpwr scs8hd_fill_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_1806 vgnd vpwr scs8hd_decap_12
XFILLER_2_4521 vgnd vpwr scs8hd_decap_12
XFILLER_7_1839 vgnd vpwr scs8hd_decap_3
XFILLER_5_2253 vpwr vgnd scs8hd_fill_2
XFILLER_5_1574 vgnd vpwr scs8hd_decap_12
XFILLER_1_1416 vgnd vpwr scs8hd_decap_12
XFILLER_0_788 vgnd vpwr scs8hd_decap_12
XFILLER_2_3875 vgnd vpwr scs8hd_decap_12
XFILLER_8_800 vgnd vpwr scs8hd_decap_12
XPHY_695 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_684 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_673 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_662 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_651 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_640 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_7_4454 vgnd vpwr scs8hd_decap_12
XFILLER_7_354 vgnd vpwr scs8hd_decap_12
XFILLER_6_1349 vgnd vpwr scs8hd_decap_12
XFILLER_3_4307 vgnd vpwr scs8hd_decap_12
XFILLER_3_2916 vgnd vpwr scs8hd_decap_12
XFILLER_1_4075 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_2838 vgnd vpwr scs8hd_decap_12
XFILLER_6_3252 vgnd vpwr scs8hd_decap_12
XFILLER_2_1703 vgnd vpwr scs8hd_decap_12
XFILLER_2_2459 vgnd vpwr scs8hd_decap_12
XFILLER_0_1482 vgnd vpwr scs8hd_decap_6
XFILLER_0_2183 vgnd vpwr scs8hd_decap_12
XFILLER_8_129 vgnd vpwr scs8hd_decap_12
XFILLER_4_324 vgnd vpwr scs8hd_decap_12
XFILLER_7_3038 vgnd vpwr scs8hd_decap_12
XFILLER_5_2050 vgnd vpwr scs8hd_decap_12
XFILLER_4_3948 vgnd vpwr scs8hd_decap_12
XFILLER_0_552 vgnd vpwr scs8hd_decap_6
XFILLER_1_1257 vgnd vpwr scs8hd_decap_12
XFILLER_2_2960 vgnd vpwr scs8hd_decap_12
XPHY_492 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_481 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_470 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_4527 vgnd vpwr scs8hd_decap_12
XFILLER_9_3826 vgnd vpwr scs8hd_decap_12
XFILLER_7_4295 vgnd vpwr scs8hd_decap_12
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_2746 vgnd vpwr scs8hd_decap_12
XFILLER_1_3160 vgnd vpwr scs8hd_decap_12
XFILLER_8_2679 vgnd vpwr scs8hd_decap_12
XFILLER_8_1923 vgnd vpwr scs8hd_decap_12
XFILLER_6_3082 vgnd vpwr scs8hd_decap_12
XFILLER_6_2370 vgnd vpwr scs8hd_decap_12
XFILLER_6_1691 vgnd vpwr scs8hd_decap_12
XFILLER_2_1544 vgnd vpwr scs8hd_decap_12
XFILLER_2_2289 vgnd vpwr scs8hd_decap_8
XFILLER_9_416 vgnd vpwr scs8hd_decap_12
XFILLER_7_2123 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_611 vgnd vpwr scs8hd_decap_12
XFILLER_4_4424 vgnd vpwr scs8hd_decap_12
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_7_1477 vgnd vpwr scs8hd_decap_12
XFILLER_4_3789 vgnd vpwr scs8hd_decap_12
XFILLER_0_2908 vgnd vpwr scs8hd_decap_6
XFILLER_0_3609 vgnd vpwr scs8hd_decap_12
XFILLER_2_4192 vgnd vpwr scs8hd_decap_12
XFILLER_8_471 vgnd vpwr scs8hd_decap_12
XFILLER_9_2977 vgnd vpwr scs8hd_decap_12
XFILLER_7_3380 vgnd vpwr scs8hd_decap_12
XFILLER_5_2819 vgnd vpwr scs8hd_decap_12
XFILLER_3_2587 vgnd vpwr scs8hd_decap_12
XFILLER_3_1831 vgnd vpwr scs8hd_decap_12
XFILLER_8_3155 vgnd vpwr scs8hd_decap_12
XFILLER_8_1764 vgnd vpwr scs8hd_decap_12
XFILLER_4_3008 vgnd vpwr scs8hd_decap_12
XFILLER_3_4490 vgnd vpwr scs8hd_decap_12
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_1_3929 vgnd vpwr scs8hd_decap_12
XFILLER_2_2020 vgnd vpwr scs8hd_decap_12
XFILLER_2_1374 vgnd vpwr scs8hd_decap_12
XFILLER_5_452 vgnd vpwr scs8hd_decap_12
XFILLER_4_4265 vgnd vpwr scs8hd_decap_12
XFILLER_4_2874 vgnd vpwr scs8hd_decap_12
XFILLER_9_4198 vgnd vpwr scs8hd_decap_12
XFILLER_9_3442 vgnd vpwr scs8hd_decap_12
XFILLER_9_3497 vgnd vpwr scs8hd_decap_6
XFILLER_9_2741 vgnd vpwr scs8hd_decap_12
XFILLER_5_1904 vgnd vpwr scs8hd_decap_12
XFILLER_3_3063 vgnd vpwr scs8hd_decap_12
XFILLER_3_1672 vgnd vpwr scs8hd_decap_12
XFILLER_0_3962 vgnd vpwr scs8hd_decap_6
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
XFILLER_8_2240 vgnd vpwr scs8hd_decap_12
XFILLER_5_4563 vgnd vpwr scs8hd_decap_12
XFILLER_3_989 vgnd vpwr scs8hd_decap_12
XFILLER_1_4405 vgnd vpwr scs8hd_decap_12
XFILLER_2_422 vgnd vpwr scs8hd_decap_12
XFILLER_4_1447 vgnd vpwr scs8hd_decap_12
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XFILLER_6_4338 vgnd vpwr scs8hd_decap_12
XFILLER_9_2059 vgnd vpwr scs8hd_decap_12
XFILLER_9_1358 vgnd vpwr scs8hd_decap_6
XFILLER_9_1303 vgnd vpwr scs8hd_decap_12
XFILLER_6_2947 vgnd vpwr scs8hd_decap_12
XFILLER_5_293 vgnd vpwr scs8hd_decap_12
XFILLER_4_3350 vgnd vpwr scs8hd_decap_12
XFILLER_0_3225 vgnd vpwr scs8hd_decap_12
XFILLER_0_1823 vgnd vpwr scs8hd_decap_6
XFILLER_0_2524 vgnd vpwr scs8hd_decap_12
XFILLER_5_3136 vgnd vpwr scs8hd_decap_12
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_9_1892 vgnd vpwr scs8hd_decap_12
XFILLER_5_1745 vgnd vpwr scs8hd_decap_12
XPHY_888 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_877 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_866 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_855 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_844 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_833 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_822 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_811 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_800 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_899 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_525 vgnd vpwr scs8hd_decap_12
XFILLER_3_720 vgnd vpwr scs8hd_decap_12
XFILLER_8_2081 vgnd vpwr scs8hd_decap_12
XFILLER_5_4393 vgnd vpwr scs8hd_decap_12
XFILLER_1_4246 vgnd vpwr scs8hd_decap_12
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XFILLER_4_1288 vgnd vpwr scs8hd_decap_12
XFILLER_1_2855 vgnd vpwr scs8hd_decap_12
XFILLER_6_3423 vgnd vpwr scs8hd_decap_12
XFILLER_6_2777 vgnd vpwr scs8hd_decap_12
XFILLER_5_1008 vgnd vpwr scs8hd_decap_12
XFILLER_4_3191 vgnd vpwr scs8hd_decap_12
XFILLER_0_2321 vpwr vgnd scs8hd_fill_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XFILLER_0_1675 vgnd vpwr scs8hd_decap_12
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3209 vgnd vpwr scs8hd_decap_12
XANTENNA__10__A _10_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_1818 vgnd vpwr scs8hd_decap_12
XFILLER_5_2221 vgnd vpwr scs8hd_decap_12
XFILLER_2_4533 vgnd vpwr scs8hd_decap_12
XFILLER_0_745 vgnd vpwr scs8hd_decap_12
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_1_1428 vgnd vpwr scs8hd_decap_12
XFILLER_2_3887 vgnd vpwr scs8hd_decap_12
XFILLER_8_812 vgnd vpwr scs8hd_decap_12
XPHY_696 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_685 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_674 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_663 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_652 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_641 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_630 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4466 vgnd vpwr scs8hd_decap_12
XFILLER_3_4319 vgnd vpwr scs8hd_decap_12
XFILLER_3_550 vgnd vpwr scs8hd_decap_12
XFILLER_1_3331 vgnd vpwr scs8hd_decap_12
XFILLER_1_1940 vgnd vpwr scs8hd_decap_12
XFILLER_1_2685 vgnd vpwr scs8hd_decap_12
XFILLER_2_3106 vgnd vpwr scs8hd_decap_12
XFILLER_6_1862 vgnd vpwr scs8hd_decap_12
XFILLER_0_2140 vgnd vpwr scs8hd_decap_12
XFILLER_2_1715 vgnd vpwr scs8hd_decap_12
XFILLER_0_2195 vgnd vpwr scs8hd_decap_6
XANTENNA__05__A _13_/C vgnd vpwr scs8hd_diode_2
XFILLER_7_2327 vpwr vgnd scs8hd_fill_2
XFILLER_7_1648 vgnd vpwr scs8hd_decap_12
XFILLER_5_2062 vgnd vpwr scs8hd_decap_12
XFILLER_2_4363 vgnd vpwr scs8hd_decap_12
XFILLER_1_1269 vgnd vpwr scs8hd_decap_12
XFILLER_2_2972 vgnd vpwr scs8hd_decap_12
XFILLER_9_4539 vgnd vpwr scs8hd_decap_12
XFILLER_8_642 vgnd vpwr scs8hd_decap_12
XPHY_493 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_482 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_471 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_460 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3838 vgnd vpwr scs8hd_decap_6
XFILLER_7_3551 vgnd vpwr scs8hd_decap_12
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_4149 vgnd vpwr scs8hd_decap_12
XFILLER_3_3404 vgnd vpwr scs8hd_decap_12
XFILLER_3_391 vgnd vpwr scs8hd_decap_12
XFILLER_3_2758 vgnd vpwr scs8hd_decap_12
XFILLER_1_1770 vgnd vpwr scs8hd_decap_12
XFILLER_8_3326 vgnd vpwr scs8hd_decap_12
XFILLER_1_306 vgnd vpwr scs8hd_decap_12
XFILLER_8_1935 vgnd vpwr scs8hd_decap_12
XFILLER_6_3094 vgnd vpwr scs8hd_decap_12
XFILLER_6_2382 vgnd vpwr scs8hd_decap_12
XFILLER_9_428 vgnd vpwr scs8hd_decap_6
XFILLER_5_623 vgnd vpwr scs8hd_decap_12
XFILLER_4_4436 vgnd vpwr scs8hd_decap_12
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_1489 vgnd vpwr scs8hd_decap_12
XFILLER_1_1099 vgnd vpwr scs8hd_decap_12
XFILLER_9_4303 vgnd vpwr scs8hd_decap_6
XFILLER_9_962 vgnd vpwr scs8hd_decap_12
XFILLER_8_483 vgnd vpwr scs8hd_decap_12
XPHY_290 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_2989 vgnd vpwr scs8hd_decap_12
XFILLER_7_3392 vgnd vpwr scs8hd_decap_12
XFILLER_3_3234 vgnd vpwr scs8hd_decap_12
XFILLER_3_2599 vgnd vpwr scs8hd_decap_12
XFILLER_3_1843 vgnd vpwr scs8hd_decap_12
XFILLER_8_3167 vgnd vpwr scs8hd_decap_12
XFILLER_8_2411 vgnd vpwr scs8hd_decap_12
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_8_1776 vgnd vpwr scs8hd_decap_12
XFILLER_4_1618 vgnd vpwr scs8hd_decap_12
XFILLER_2_2032 vgnd vpwr scs8hd_decap_12
XFILLER_2_1386 vgnd vpwr scs8hd_decap_12
XFILLER_6_4509 vgnd vpwr scs8hd_decap_12
XFILLER_6_910 vgnd vpwr scs8hd_decap_12
XFILLER_5_464 vgnd vpwr scs8hd_decap_12
XFILLER_4_4277 vgnd vpwr scs8hd_decap_12
XFILLER_4_3521 vgnd vpwr scs8hd_decap_12
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_4_2886 vgnd vpwr scs8hd_decap_12
XFILLER_9_4155 vgnd vpwr scs8hd_decap_12
XFILLER_9_3454 vgnd vpwr scs8hd_decap_12
XFILLER_9_2753 vgnd vpwr scs8hd_decap_6
XFILLER_5_3307 vgnd vpwr scs8hd_decap_12
XFILLER_5_1916 vgnd vpwr scs8hd_decap_12
XFILLER_3_3075 vgnd vpwr scs8hd_decap_12
XFILLER_3_2363 vgnd vpwr scs8hd_decap_12
XFILLER_3_2352 vgnd vpwr scs8hd_decap_4
XFILLER_3_1684 vgnd vpwr scs8hd_decap_12
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
XANTENNA__13__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_2252 vgnd vpwr scs8hd_decap_12
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_4417 vgnd vpwr scs8hd_decap_12
XFILLER_2_434 vgnd vpwr scs8hd_decap_12
XFILLER_4_1459 vgnd vpwr scs8hd_decap_12
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XFILLER_9_2016 vgnd vpwr scs8hd_decap_12
XFILLER_6_751 vgnd vpwr scs8hd_decap_12
XFILLER_9_1315 vgnd vpwr scs8hd_decap_12
XFILLER_7_1050 vgnd vpwr scs8hd_decap_12
XFILLER_4_3362 vgnd vpwr scs8hd_decap_12
XFILLER_0_3237 vgnd vpwr scs8hd_decap_12
XFILLER_4_1971 vgnd vpwr scs8hd_decap_12
XFILLER_0_2536 vgnd vpwr scs8hd_decap_6
XFILLER_5_3148 vgnd vpwr scs8hd_decap_12
XFILLER_5_1757 vgnd vpwr scs8hd_decap_12
XFILLER_3_2160 vgnd vpwr scs8hd_decap_12
XANTENNA__08__A address[2] vgnd vpwr scs8hd_diode_2
XPHY_889 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_878 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_867 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_856 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_845 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_834 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_823 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_812 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_801 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_537 vgnd vpwr scs8hd_decap_12
XFILLER_8_2093 vgnd vpwr scs8hd_decap_12
XFILLER_1_3502 vgnd vpwr scs8hd_decap_12
XFILLER_1_4258 vgnd vpwr scs8hd_decap_12
XFILLER_6_3435 vgnd vpwr scs8hd_decap_12
XFILLER_6_581 vgnd vpwr scs8hd_decap_12
XFILLER_6_2789 vgnd vpwr scs8hd_decap_12
XFILLER_0_2344 vpwr vgnd scs8hd_fill_2
XFILLER_0_3001 vgnd vpwr scs8hd_decap_6
XFILLER_0_1687 vgnd vpwr scs8hd_decap_12
XFILLER_0_2388 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_507 vgnd vpwr scs8hd_decap_12
XFILLER_9_3070 vgnd vpwr scs8hd_decap_12
XFILLER_5_2266 vgnd vpwr scs8hd_decap_12
XFILLER_5_2233 vgnd vpwr scs8hd_decap_12
XANTENNA__10__B enable vgnd vpwr scs8hd_diode_2
XFILLER_2_4578 vgnd vpwr scs8hd_decap_3
XFILLER_0_757 vgnd vpwr scs8hd_decap_12
XPHY_620 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_1587 vgnd vpwr scs8hd_decap_12
XFILLER_0_3590 vgnd vpwr scs8hd_decap_6
XFILLER_0_4291 vgnd vpwr scs8hd_decap_12
XFILLER_2_3899 vgnd vpwr scs8hd_decap_12
XPHY_697 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_686 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_675 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_664 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_653 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_642 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_631 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_4478 vgnd vpwr scs8hd_decap_12
XFILLER_7_3722 vgnd vpwr scs8hd_decap_12
XFILLER_6_2008 vgnd vpwr scs8hd_decap_12
XFILLER_7_367 vgnd vpwr scs8hd_decap_12
XFILLER_3_562 vgnd vpwr scs8hd_decap_12
XFILLER_5_3490 vgnd vpwr scs8hd_decap_12
XFILLER_4_1020 vgnd vpwr scs8hd_decap_12
XFILLER_3_2929 vgnd vpwr scs8hd_decap_12
XFILLER_1_3343 vgnd vpwr scs8hd_decap_12
XFILLER_1_4088 vgnd vpwr scs8hd_decap_12
XFILLER_1_2697 vgnd vpwr scs8hd_decap_12
XFILLER_6_3265 vgnd vpwr scs8hd_decap_12
XFILLER_6_2520 vgnd vpwr scs8hd_decap_12
XFILLER_2_3118 vgnd vpwr scs8hd_decap_12
XFILLER_6_1874 vgnd vpwr scs8hd_decap_12
XFILLER_0_1451 vgnd vpwr scs8hd_decap_6
XFILLER_0_2152 vgnd vpwr scs8hd_decap_12
XFILLER_2_1727 vgnd vpwr scs8hd_decap_12
XANTENNA__05__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_2339 vgnd vpwr scs8hd_decap_12
XFILLER_7_2306 vgnd vpwr scs8hd_decap_12
XFILLER_4_337 vgnd vpwr scs8hd_decap_12
XFILLER_0_521 vgnd vpwr scs8hd_decap_6
XANTENNA__21__A gfpga_pad_GPIO_PAD[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_4375 vgnd vpwr scs8hd_decap_12
XPHY_461 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_450 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_2984 vgnd vpwr scs8hd_decap_12
XFILLER_8_654 vgnd vpwr scs8hd_decap_12
XPHY_494 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_483 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_472 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3563 vgnd vpwr scs8hd_decap_12
XFILLER_1_3173 vgnd vpwr scs8hd_decap_12
XFILLER_1_1782 vgnd vpwr scs8hd_decap_12
XFILLER_8_3338 vgnd vpwr scs8hd_decap_12
XFILLER_8_80 vgnd vpwr scs8hd_decap_12
XFILLER_1_318 vgnd vpwr scs8hd_decap_12
XFILLER_8_1947 vgnd vpwr scs8hd_decap_12
XFILLER_6_2394 vgnd vpwr scs8hd_decap_12
XFILLER_2_2203 vgnd vpwr scs8hd_decap_12
XANTENNA__16__A gfpga_pad_GPIO_PAD[5] vgnd vpwr scs8hd_diode_2
XFILLER_2_1557 vgnd vpwr scs8hd_decap_12
XFILLER_5_635 vgnd vpwr scs8hd_decap_12
XFILLER_8_3850 vgnd vpwr scs8hd_decap_12
XFILLER_7_2136 vgnd vpwr scs8hd_decap_12
XFILLER_4_4448 vgnd vpwr scs8hd_decap_12
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_830 vgnd vpwr scs8hd_decap_12
XFILLER_0_373 vgnd vpwr scs8hd_decap_12
XFILLER_1_1001 vgnd vpwr scs8hd_decap_12
XFILLER_2_3460 vgnd vpwr scs8hd_decap_12
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_291 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_2946 vgnd vpwr scs8hd_decap_12
XFILLER_9_974 vgnd vpwr scs8hd_decap_12
XFILLER_8_495 vgnd vpwr scs8hd_decap_12
XFILLER_4_690 vgnd vpwr scs8hd_decap_12
XFILLER_3_3246 vgnd vpwr scs8hd_decap_12
XFILLER_3_1855 vgnd vpwr scs8hd_decap_12
XFILLER_8_3179 vgnd vpwr scs8hd_decap_12
XFILLER_8_2445 vgnd vpwr scs8hd_decap_12
XFILLER_8_2423 vgnd vpwr scs8hd_decap_12
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XFILLER_2_605 vgnd vpwr scs8hd_decap_12
XFILLER_8_1788 vgnd vpwr scs8hd_decap_12
XFILLER_6_2191 vgnd vpwr scs8hd_decap_12
XFILLER_2_1398 vgnd vpwr scs8hd_decap_12
XFILLER_6_922 vgnd vpwr scs8hd_decap_12
XFILLER_5_476 vgnd vpwr scs8hd_decap_12
XFILLER_7_1221 vgnd vpwr scs8hd_decap_12
XFILLER_4_4289 vgnd vpwr scs8hd_decap_12
XFILLER_4_3533 vgnd vpwr scs8hd_decap_12
XFILLER_0_2729 vgnd vpwr scs8hd_decap_12
XFILLER_9_4167 vgnd vpwr scs8hd_decap_12
XFILLER_9_3466 vgnd vpwr scs8hd_decap_6
XFILLER_9_3411 vgnd vpwr scs8hd_decap_12
XFILLER_9_2710 vgnd vpwr scs8hd_decap_12
XFILLER_5_3319 vgnd vpwr scs8hd_decap_12
XFILLER_5_1928 vgnd vpwr scs8hd_decap_12
XFILLER_3_3087 vgnd vpwr scs8hd_decap_12
XFILLER_3_2375 vgnd vpwr scs8hd_decap_4
XFILLER_0_3931 vgnd vpwr scs8hd_decap_6
XFILLER_3_1696 vgnd vpwr scs8hd_decap_12
XFILLER_7_708 vgnd vpwr scs8hd_decap_12
XANTENNA__13__B _11_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_903 vgnd vpwr scs8hd_decap_12
XFILLER_8_2264 vgnd vpwr scs8hd_decap_12
XFILLER_5_4576 vgnd vpwr scs8hd_decap_4
XFILLER_5_3831 vgnd vpwr scs8hd_decap_12
XFILLER_4_2106 vgnd vpwr scs8hd_decap_12
XFILLER_1_4429 vgnd vpwr scs8hd_decap_12
XFILLER_2_446 vgnd vpwr scs8hd_decap_12
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
XFILLER_9_2028 vgnd vpwr scs8hd_decap_12
XFILLER_9_1327 vgnd vpwr scs8hd_decap_6
XFILLER_6_3606 vgnd vpwr scs8hd_decap_12
XFILLER_7_1062 vgnd vpwr scs8hd_decap_12
XFILLER_4_3374 vgnd vpwr scs8hd_decap_12
XFILLER_0_3249 vgnd vpwr scs8hd_decap_6
XFILLER_9_590 vgnd vpwr scs8hd_decap_12
XFILLER_9_1861 vgnd vpwr scs8hd_decap_12
XPHY_802 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_2172 vgnd vpwr scs8hd_decap_12
XFILLER_0_3783 vgnd vpwr scs8hd_decap_12
XPHY_879 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_868 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_857 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_846 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_835 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_824 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_813 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_733 vgnd vpwr scs8hd_decap_12
XFILLER_5_3661 vgnd vpwr scs8hd_decap_12
XFILLER_1_3514 vgnd vpwr scs8hd_decap_12
XFILLER_2_276 vgnd vpwr scs8hd_decap_12
XFILLER_1_2868 vgnd vpwr scs8hd_decap_12
XFILLER_9_1179 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ top_width_0_height_0__pin_14_ logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[7] vgnd vpwr scs8hd_ebufn_1
XFILLER_6_593 vgnd vpwr scs8hd_decap_12
XFILLER_0_1644 vgnd vpwr scs8hd_decap_12
XFILLER_0_2378 vpwr vgnd scs8hd_fill_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XFILLER_0_1699 vgnd vpwr scs8hd_decap_6
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3082 vgnd vpwr scs8hd_decap_12
XANTENNA__10__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_0_714 vgnd vpwr scs8hd_decap_12
XFILLER_9_2381 vgnd vpwr scs8hd_decap_6
XANTENNA__19__A gfpga_pad_GPIO_PAD[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_2278 vgnd vpwr scs8hd_decap_12
XFILLER_5_2245 vgnd vpwr scs8hd_decap_8
XFILLER_2_4546 vgnd vpwr scs8hd_decap_12
XFILLER_0_769 vgnd vpwr scs8hd_decap_6
XFILLER_2_3801 vgnd vpwr scs8hd_decap_12
XPHY_610 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_643 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_632 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_621 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_1599 vgnd vpwr scs8hd_decap_12
XFILLER_8_825 vgnd vpwr scs8hd_decap_12
XPHY_698 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_687 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_676 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_665 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_654 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_379 vgnd vpwr scs8hd_decap_12
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XFILLER_7_3734 vgnd vpwr scs8hd_decap_12
XFILLER_3_574 vgnd vpwr scs8hd_decap_12
XFILLER_4_1032 vgnd vpwr scs8hd_decap_12
XFILLER_1_1953 vgnd vpwr scs8hd_decap_12
XFILLER_8_3509 vgnd vpwr scs8hd_decap_12
XFILLER_7_891 vgnd vpwr scs8hd_decap_12
XFILLER_6_3277 vgnd vpwr scs8hd_decap_12
XFILLER_2_2407 vgnd vpwr scs8hd_decap_3
XFILLER_6_1886 vgnd vpwr scs8hd_decap_12
XFILLER_0_2164 vgnd vpwr scs8hd_decap_6
XFILLER_5_806 vgnd vpwr scs8hd_decap_12
XANTENNA__05__C address[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_349 vgnd vpwr scs8hd_decap_12
XFILLER_5_2075 vgnd vpwr scs8hd_decap_12
XFILLER_5_1330 vgnd vpwr scs8hd_decap_12
XFILLER_2_4387 vgnd vpwr scs8hd_decap_12
XFILLER_2_2996 vgnd vpwr scs8hd_decap_12
XFILLER_2_3631 vgnd vpwr scs8hd_decap_12
XPHY_495 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_484 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_473 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_462 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_451 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_440 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_4508 vgnd vpwr scs8hd_decap_12
XFILLER_9_3807 vgnd vpwr scs8hd_decap_6
XFILLER_8_666 vgnd vpwr scs8hd_decap_12
XFILLER_7_4210 vgnd vpwr scs8hd_decap_12
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
XFILLER_4_861 vgnd vpwr scs8hd_decap_12
XFILLER_7_3575 vgnd vpwr scs8hd_decap_12
XFILLER_6_1105 vgnd vpwr scs8hd_decap_12
XFILLER_3_3417 vgnd vpwr scs8hd_decap_12
XFILLER_1_1794 vgnd vpwr scs8hd_decap_12
XFILLER_1_3185 vgnd vpwr scs8hd_decap_12
XFILLER_8_1959 vgnd vpwr scs8hd_decap_12
XFILLER_2_2215 vgnd vpwr scs8hd_decap_12
XFILLER_2_1569 vgnd vpwr scs8hd_decap_12
XFILLER_5_647 vgnd vpwr scs8hd_decap_12
XFILLER_8_3862 vgnd vpwr scs8hd_decap_12
XFILLER_7_2148 vgnd vpwr scs8hd_decap_12
XFILLER_4_3704 vgnd vpwr scs8hd_decap_12
XFILLER_1_842 vgnd vpwr scs8hd_decap_12
XFILLER_0_385 vgnd vpwr scs8hd_decap_12
XFILLER_5_1160 vgnd vpwr scs8hd_decap_12
XFILLER_1_1013 vgnd vpwr scs8hd_decap_12
XFILLER_2_3472 vgnd vpwr scs8hd_decap_12
XFILLER_9_986 vgnd vpwr scs8hd_decap_6
XFILLER_9_931 vgnd vpwr scs8hd_decap_12
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_292 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3659 vgnd vpwr scs8hd_decap_12
XFILLER_9_2958 vgnd vpwr scs8hd_decap_12
XFILLER_7_4051 vgnd vpwr scs8hd_decap_12
XFILLER_7_2660 vgnd vpwr scs8hd_decap_12
XFILLER_3_3258 vgnd vpwr scs8hd_decap_12
XFILLER_3_2502 vgnd vpwr scs8hd_decap_12
XFILLER_3_1867 vgnd vpwr scs8hd_decap_12
XFILLER_1_2270 vgnd vpwr scs8hd_decap_12
XFILLER_8_2457 vgnd vpwr scs8hd_decap_12
XFILLER_8_2435 vpwr vgnd scs8hd_fill_2
XFILLER_2_617 vgnd vpwr scs8hd_decap_12
XFILLER_3_3770 vgnd vpwr scs8hd_decap_12
XFILLER_2_1300 vgnd vpwr scs8hd_decap_12
XFILLER_2_2045 vgnd vpwr scs8hd_decap_12
XFILLER_9_249 vgnd vpwr scs8hd_decap_12
XFILLER_6_934 vgnd vpwr scs8hd_decap_12
XFILLER_8_3692 vgnd vpwr scs8hd_decap_12
XFILLER_7_1233 vgnd vpwr scs8hd_decap_12
XFILLER_4_3545 vgnd vpwr scs8hd_decap_12
XFILLER_4_2899 vgnd vpwr scs8hd_decap_12
XFILLER_1_672 vgnd vpwr scs8hd_decap_12
XFILLER_9_4124 vgnd vpwr scs8hd_decap_12
XFILLER_9_3423 vgnd vpwr scs8hd_decap_12
XFILLER_9_4179 vgnd vpwr scs8hd_decap_6
XFILLER_9_2722 vgnd vpwr scs8hd_decap_6
XFILLER_8_1008 vgnd vpwr scs8hd_decap_12
XFILLER_3_3099 vgnd vpwr scs8hd_decap_12
XFILLER_3_2310 vpwr vgnd scs8hd_fill_2
XANTENNA__13__C _13_/C vgnd vpwr scs8hd_diode_2
XFILLER_8_2276 vgnd vpwr scs8hd_decap_12
XFILLER_8_1520 vgnd vpwr scs8hd_decap_12
XFILLER_4_2118 vgnd vpwr scs8hd_decap_12
XFILLER_2_1130 vgnd vpwr scs8hd_decap_12
XFILLER_6_764 vgnd vpwr scs8hd_decap_12
XFILLER_6_3618 vgnd vpwr scs8hd_decap_12
XFILLER_4_4021 vgnd vpwr scs8hd_decap_12
XFILLER_7_1074 vgnd vpwr scs8hd_decap_12
XFILLER_4_2630 vgnd vpwr scs8hd_decap_12
XFILLER_4_1984 vgnd vpwr scs8hd_decap_12
XFILLER_0_2505 vgnd vpwr scs8hd_decap_6
XFILLER_0_3206 vgnd vpwr scs8hd_decap_12
XFILLER_9_2574 vgnd vpwr scs8hd_decap_12
XFILLER_9_1873 vgnd vpwr scs8hd_decap_12
XPHY_836 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_825 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_814 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_803 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_2184 vgnd vpwr scs8hd_decap_12
XFILLER_0_3795 vgnd vpwr scs8hd_decap_6
XFILLER_0_4496 vgnd vpwr scs8hd_decap_12
XPHY_869 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_858 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_847 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3905 vgnd vpwr scs8hd_decap_12
XFILLER_3_745 vgnd vpwr scs8hd_decap_12
XFILLER_2_288 vgnd vpwr scs8hd_decap_12
XFILLER_8_1361 vgnd vpwr scs8hd_decap_12
XFILLER_5_3673 vgnd vpwr scs8hd_decap_12
XFILLER_4_1203 vgnd vpwr scs8hd_decap_12
XFILLER_1_3526 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _13_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_3448 vgnd vpwr scs8hd_decap_12
XFILLER_6_2703 vgnd vpwr scs8hd_decap_12
XFILLER_0_1656 vgnd vpwr scs8hd_decap_12
XFILLER_0_2357 vgnd vpwr scs8hd_decap_12
XFILLER_9_3094 vgnd vpwr scs8hd_decap_6
XFILLER_6_3960 vgnd vpwr scs8hd_decap_12
XANTENNA__10__D _10_/D vgnd vpwr scs8hd_diode_2
XFILLER_0_726 vgnd vpwr scs8hd_decap_12
XFILLER_5_1501 vgnd vpwr scs8hd_decap_12
XFILLER_2_4558 vgnd vpwr scs8hd_decap_12
XFILLER_0_4260 vgnd vpwr scs8hd_decap_12
XPHY_611 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_677 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_600 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_666 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_655 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_644 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_633 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_622 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xlogical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _07_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_837 vgnd vpwr scs8hd_decap_12
XPHY_699 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_688 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XFILLER_7_3746 vgnd vpwr scs8hd_decap_12
XFILLER_3_586 vgnd vpwr scs8hd_decap_12
XFILLER_1_4002 vgnd vpwr scs8hd_decap_12
XFILLER_8_1191 vgnd vpwr scs8hd_decap_12
XFILLER_4_1044 vgnd vpwr scs8hd_decap_12
XFILLER_1_1965 vgnd vpwr scs8hd_decap_12
XFILLER_1_2611 vgnd vpwr scs8hd_decap_12
XFILLER_1_3356 vgnd vpwr scs8hd_decap_12
XFILLER_6_3289 vgnd vpwr scs8hd_decap_12
XFILLER_6_2533 vgnd vpwr scs8hd_decap_12
XFILLER_6_1898 vgnd vpwr scs8hd_decap_12
XFILLER_0_2121 vgnd vpwr scs8hd_decap_12
XFILLER_1_4580 vgnd vpwr scs8hd_fill_1
XFILLER_0_1420 vgnd vpwr scs8hd_decap_6
XANTENNA__05__D enable vgnd vpwr scs8hd_diode_2
XFILLER_5_818 vgnd vpwr scs8hd_decap_12
XFILLER_7_2319 vgnd vpwr scs8hd_decap_8
XFILLER_5_2087 vgnd vpwr scs8hd_decap_12
XFILLER_2_4399 vgnd vpwr scs8hd_decap_12
XFILLER_2_3643 vgnd vpwr scs8hd_decap_12
XPHY_496 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_485 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_474 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_463 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_452 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_441 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_430 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_678 vgnd vpwr scs8hd_decap_12
XFILLER_7_4222 vgnd vpwr scs8hd_decap_12
XFILLER_4_873 vgnd vpwr scs8hd_decap_12
XFILLER_7_3587 vgnd vpwr scs8hd_decap_12
XFILLER_7_2831 vgnd vpwr scs8hd_decap_12
XFILLER_6_1117 vgnd vpwr scs8hd_decap_12
XFILLER_3_3429 vgnd vpwr scs8hd_decap_12
XFILLER_1_2441 vgnd vpwr scs8hd_decap_12
XFILLER_1_3197 vgnd vpwr scs8hd_decap_12
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_2606 vgnd vpwr scs8hd_decap_12
XFILLER_3_3941 vgnd vpwr scs8hd_decap_12
XFILLER_0_1272 vgnd vpwr scs8hd_decap_12
XFILLER_5_659 vgnd vpwr scs8hd_decap_12
XFILLER_7_1404 vgnd vpwr scs8hd_decap_12
XFILLER_4_3716 vgnd vpwr scs8hd_decap_12
XFILLER_0_342 vgnd vpwr scs8hd_decap_12
XFILLER_0_397 vgnd vpwr scs8hd_decap_6
XFILLER_2_3484 vgnd vpwr scs8hd_decap_12
XFILLER_5_1172 vgnd vpwr scs8hd_decap_12
XFILLER_1_1025 vgnd vpwr scs8hd_decap_12
XFILLER_9_943 vgnd vpwr scs8hd_decap_12
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_293 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_2915 vgnd vpwr scs8hd_decap_12
XFILLER_7_4063 vgnd vpwr scs8hd_decap_12
XFILLER_7_2672 vgnd vpwr scs8hd_decap_12
XFILLER_3_2514 vgnd vpwr scs8hd_decap_12
XFILLER_3_1879 vgnd vpwr scs8hd_decap_12
XFILLER_1_2282 vgnd vpwr scs8hd_decap_4
XFILLER_1_2293 vpwr vgnd scs8hd_fill_2
XFILLER_2_629 vgnd vpwr scs8hd_decap_12
XFILLER_8_2469 vpwr vgnd scs8hd_fill_2
XFILLER_2_2057 vgnd vpwr scs8hd_decap_12
XFILLER_8_4350 vgnd vpwr scs8hd_decap_12
XFILLER_5_489 vgnd vpwr scs8hd_decap_12
XFILLER_7_1245 vgnd vpwr scs8hd_decap_12
XFILLER_4_3557 vgnd vpwr scs8hd_decap_12
XFILLER_4_2801 vgnd vpwr scs8hd_decap_12
XFILLER_1_684 vgnd vpwr scs8hd_decap_12
XFILLER_9_4136 vgnd vpwr scs8hd_decap_12
XFILLER_9_3435 vgnd vpwr scs8hd_decap_6
XFILLER_0_3900 vgnd vpwr scs8hd_decap_6
XANTENNA__13__D _10_/D vgnd vpwr scs8hd_diode_2
XFILLER_3_916 vgnd vpwr scs8hd_decap_12
XFILLER_2_459 vgnd vpwr scs8hd_decap_12
XFILLER_8_1532 vgnd vpwr scs8hd_decap_12
XFILLER_5_3844 vgnd vpwr scs8hd_decap_12
XFILLER_2_1142 vgnd vpwr scs8hd_decap_12
XFILLER_6_776 vgnd vpwr scs8hd_decap_12
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_4180 vgnd vpwr scs8hd_decap_12
XFILLER_4_4033 vgnd vpwr scs8hd_decap_12
XFILLER_4_2642 vgnd vpwr scs8hd_decap_12
XFILLER_0_3218 vgnd vpwr scs8hd_decap_6
XFILLER_2_971 vgnd vpwr scs8hd_decap_12
XFILLER_7_1086 vgnd vpwr scs8hd_decap_12
XFILLER_4_3387 vgnd vpwr scs8hd_decap_12
XFILLER_4_1996 vgnd vpwr scs8hd_decap_12
XFILLER_9_3287 vgnd vpwr scs8hd_decap_12
XFILLER_9_2586 vgnd vpwr scs8hd_decap_12
XFILLER_9_1885 vgnd vpwr scs8hd_decap_6
XFILLER_9_1830 vgnd vpwr scs8hd_decap_12
XFILLER_5_2439 vgnd vpwr scs8hd_fill_1
XFILLER_3_1440 vgnd vpwr scs8hd_decap_12
XFILLER_0_3752 vgnd vpwr scs8hd_decap_12
XPHY_859 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_848 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_837 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_826 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_815 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_804 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3917 vgnd vpwr scs8hd_decap_12
XFILLER_5_3685 vgnd vpwr scs8hd_decap_12
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_757 vgnd vpwr scs8hd_decap_12
XFILLER_4_1215 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_4106 vgnd vpwr scs8hd_decap_12
XFILLER_9_1148 vgnd vpwr scs8hd_decap_12
XFILLER_4_2472 vgnd vpwr scs8hd_decap_12
XFILLER_4_2461 vgnd vpwr scs8hd_decap_8
XFILLER_0_1668 vgnd vpwr scs8hd_decap_6
XFILLER_0_1613 vgnd vpwr scs8hd_decap_12
XFILLER_0_2369 vgnd vpwr scs8hd_decap_6
XFILLER_9_3051 vgnd vpwr scs8hd_decap_12
XFILLER_9_2350 vgnd vpwr scs8hd_decap_6
XFILLER_6_3972 vgnd vpwr scs8hd_decap_12
XFILLER_0_738 vgnd vpwr scs8hd_decap_6
XFILLER_2_3814 vgnd vpwr scs8hd_decap_12
XFILLER_5_1513 vgnd vpwr scs8hd_decap_12
XFILLER_0_4272 vgnd vpwr scs8hd_decap_6
XPHY_689 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_612 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_678 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_601 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_667 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_656 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_645 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_634 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_623 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_849 vgnd vpwr scs8hd_decap_12
XFILLER_7_3758 vgnd vpwr scs8hd_decap_12
XFILLER_5_4161 vgnd vpwr scs8hd_decap_12
XFILLER_5_2770 vgnd vpwr scs8hd_decap_12
XFILLER_3_598 vgnd vpwr scs8hd_decap_12
XFILLER_1_3368 vgnd vpwr scs8hd_decap_12
XFILLER_1_4014 vgnd vpwr scs8hd_decap_12
XFILLER_4_1056 vgnd vpwr scs8hd_decap_12
XFILLER_1_1977 vgnd vpwr scs8hd_decap_12
XFILLER_6_2545 vgnd vpwr scs8hd_decap_12
XFILLER_0_2133 vgnd vpwr scs8hd_decap_6
XFILLER_1_3880 vgnd vpwr scs8hd_decap_12
XFILLER_2_3655 vgnd vpwr scs8hd_decap_12
XFILLER_5_2099 vgnd vpwr scs8hd_decap_12
XFILLER_5_1343 vgnd vpwr scs8hd_decap_12
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XPHY_497 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_486 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_475 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_464 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_453 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_442 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_431 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_420 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4234 vgnd vpwr scs8hd_decap_12
XFILLER_7_2843 vgnd vpwr scs8hd_decap_12
XFILLER_1_2453 vgnd vpwr scs8hd_decap_12
XFILLER_8_4009 vgnd vpwr scs8hd_decap_12
XFILLER_8_2618 vgnd vpwr scs8hd_decap_12
XFILLER_6_3021 vgnd vpwr scs8hd_decap_12
XFILLER_6_1630 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _14_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_3953 vgnd vpwr scs8hd_decap_12
XFILLER_2_2228 vgnd vpwr scs8hd_decap_12
XFILLER_0_1284 vgnd vpwr scs8hd_decap_12
XFILLER_8_4521 vgnd vpwr scs8hd_decap_12
XFILLER_8_3875 vgnd vpwr scs8hd_decap_12
XFILLER_7_1416 vgnd vpwr scs8hd_decap_12
XFILLER_5_1184 vgnd vpwr scs8hd_decap_12
XFILLER_4_3728 vgnd vpwr scs8hd_decap_12
XFILLER_1_855 vgnd vpwr scs8hd_decap_12
XFILLER_0_354 vgnd vpwr scs8hd_decap_12
XFILLER_2_2740 vgnd vpwr scs8hd_decap_12
XFILLER_2_3496 vgnd vpwr scs8hd_decap_12
XFILLER_2_4131 vgnd vpwr scs8hd_decap_12
XFILLER_9_900 vgnd vpwr scs8hd_decap_12
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3628 vgnd vpwr scs8hd_decap_12
XFILLER_9_955 vgnd vpwr scs8hd_decap_6
XFILLER_8_410 vgnd vpwr scs8hd_decap_12
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_294 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_2927 vgnd vpwr scs8hd_decap_12
XFILLER_7_4075 vgnd vpwr scs8hd_decap_12
XFILLER_3_2526 vgnd vpwr scs8hd_decap_12
XFILLER_8_1703 vgnd vpwr scs8hd_decap_12
XFILLER_6_1471 vgnd vpwr scs8hd_decap_12
XFILLER_3_3783 vgnd vpwr scs8hd_decap_12
XFILLER_2_1313 vgnd vpwr scs8hd_decap_12
XFILLER_2_2069 vgnd vpwr scs8hd_decap_12
XFILLER_9_218 vgnd vpwr scs8hd_decap_12
XFILLER_6_947 vgnd vpwr scs8hd_decap_12
XFILLER_8_2960 vgnd vpwr scs8hd_decap_12
XFILLER_4_4204 vgnd vpwr scs8hd_decap_12
XFILLER_4_2813 vgnd vpwr scs8hd_decap_12
XFILLER_1_696 vgnd vpwr scs8hd_decap_12
XFILLER_7_1257 vgnd vpwr scs8hd_decap_12
XFILLER_2_2581 vgnd vpwr scs8hd_decap_12
XFILLER_9_4148 vgnd vpwr scs8hd_decap_6
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_3160 vgnd vpwr scs8hd_decap_12
XFILLER_7_2481 vgnd vpwr scs8hd_decap_12
XFILLER_3_3002 vgnd vpwr scs8hd_decap_12
XFILLER_3_2356 vgnd vpwr scs8hd_fill_1
XFILLER_3_2323 vpwr vgnd scs8hd_fill_2
XFILLER_3_1611 vgnd vpwr scs8hd_decap_12
XFILLER_9_3981 vgnd vpwr scs8hd_decap_12
XFILLER_8_1544 vgnd vpwr scs8hd_decap_12
XFILLER_5_4502 vgnd vpwr scs8hd_decap_12
XFILLER_5_3856 vgnd vpwr scs8hd_decap_12
XFILLER_3_928 vgnd vpwr scs8hd_decap_12
XFILLER_8_2289 vgnd vpwr scs8hd_decap_12
XFILLER_1_3709 vgnd vpwr scs8hd_decap_12
XFILLER_2_1154 vgnd vpwr scs8hd_decap_12
XFILLER_9_2009 vgnd vpwr scs8hd_decap_6
XFILLER_6_788 vgnd vpwr scs8hd_decap_12
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_4192 vgnd vpwr scs8hd_decap_12
XFILLER_4_4045 vgnd vpwr scs8hd_decap_12
XFILLER_4_3399 vgnd vpwr scs8hd_decap_12
XFILLER_2_983 vgnd vpwr scs8hd_decap_12
XFILLER_9_571 vgnd vpwr scs8hd_decap_12
XFILLER_9_3299 vgnd vpwr scs8hd_decap_12
XFILLER_9_2543 vgnd vpwr scs8hd_decap_12
XFILLER_9_1842 vgnd vpwr scs8hd_decap_12
XFILLER_9_2598 vgnd vpwr scs8hd_decap_6
XFILLER_3_2197 vgnd vpwr scs8hd_decap_12
XFILLER_3_1452 vgnd vpwr scs8hd_decap_12
XFILLER_0_3764 vgnd vpwr scs8hd_decap_12
XFILLER_0_4465 vgnd vpwr scs8hd_decap_12
XPHY_849 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_838 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_827 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_816 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_805 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XFILLER_8_2020 vgnd vpwr scs8hd_decap_12
XFILLER_8_1374 vgnd vpwr scs8hd_decap_12
XFILLER_7_3929 vgnd vpwr scs8hd_decap_12
XFILLER_5_4332 vgnd vpwr scs8hd_decap_12
XFILLER_5_3697 vgnd vpwr scs8hd_decap_12
XFILLER_5_2941 vgnd vpwr scs8hd_decap_12
XFILLER_3_769 vgnd vpwr scs8hd_decap_12
XFILLER_1_3539 vgnd vpwr scs8hd_decap_12
XFILLER_4_1227 vgnd vpwr scs8hd_decap_12
XPHY_70 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_2716 vgnd vpwr scs8hd_decap_12
XFILLER_4_3130 vgnd vpwr scs8hd_decap_12
XFILLER_4_2484 vgnd vpwr scs8hd_decap_12
XFILLER_0_2304 vpwr vgnd scs8hd_fill_2
XFILLER_0_2326 vgnd vpwr scs8hd_fill_1
XFILLER_0_2348 vpwr vgnd scs8hd_fill_2
XFILLER_0_1625 vgnd vpwr scs8hd_decap_12
XFILLER_9_3063 vgnd vpwr scs8hd_decap_6
XFILLER_6_3984 vgnd vpwr scs8hd_decap_12
XFILLER_2_3826 vgnd vpwr scs8hd_decap_12
XPHY_602 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1282 vgnd vpwr scs8hd_decap_12
XPHY_613 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_679 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_668 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_657 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_646 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_635 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_624 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4405 vgnd vpwr scs8hd_decap_12
XFILLER_5_4173 vgnd vpwr scs8hd_decap_12
XFILLER_5_2782 vgnd vpwr scs8hd_decap_12
XFILLER_1_2624 vgnd vpwr scs8hd_decap_12
XFILLER_1_1989 vgnd vpwr scs8hd_decap_12
XFILLER_6_2557 vgnd vpwr scs8hd_decap_12
XFILLER_6_1801 vgnd vpwr scs8hd_decap_12
XFILLER_1_3892 vgnd vpwr scs8hd_decap_12
XFILLER_6_4460 vgnd vpwr scs8hd_decap_12
XFILLER_2_4302 vgnd vpwr scs8hd_decap_12
XFILLER_5_2001 vgnd vpwr scs8hd_decap_12
XFILLER_5_1355 vgnd vpwr scs8hd_decap_12
XFILLER_2_2911 vgnd vpwr scs8hd_decap_12
XFILLER_2_3667 vgnd vpwr scs8hd_decap_12
XPHY_443 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_432 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_421 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_410 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_1208 vgnd vpwr scs8hd_decap_12
XFILLER_0_3380 vgnd vpwr scs8hd_decap_12
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
XPHY_498 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_487 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_476 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_465 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_454 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4246 vgnd vpwr scs8hd_decap_12
XFILLER_7_2855 vgnd vpwr scs8hd_decap_12
XFILLER_4_886 vgnd vpwr scs8hd_decap_12
XFILLER_3_330 vgnd vpwr scs8hd_decap_12
XFILLER_1_2465 vgnd vpwr scs8hd_decap_12
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_6_3033 vgnd vpwr scs8hd_decap_12
XFILLER_6_2343 vgnd vpwr scs8hd_fill_1
XFILLER_6_1642 vgnd vpwr scs8hd_decap_12
XFILLER_0_1296 vgnd vpwr scs8hd_decap_6
XFILLER_0_1241 vgnd vpwr scs8hd_decap_12
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XFILLER_8_4533 vgnd vpwr scs8hd_decap_12
XFILLER_8_3887 vgnd vpwr scs8hd_decap_12
XFILLER_1_867 vgnd vpwr scs8hd_decap_12
XFILLER_0_311 vgnd vpwr scs8hd_decap_12
XFILLER_2_4143 vgnd vpwr scs8hd_decap_12
XFILLER_7_1428 vgnd vpwr scs8hd_decap_12
XFILLER_5_1196 vgnd vpwr scs8hd_decap_12
XFILLER_1_1038 vgnd vpwr scs8hd_decap_12
XFILLER_0_366 vgnd vpwr scs8hd_decap_6
XFILLER_2_2752 vgnd vpwr scs8hd_decap_12
XFILLER_9_912 vgnd vpwr scs8hd_decap_12
XFILLER_8_422 vgnd vpwr scs8hd_decap_12
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_295 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_2939 vgnd vpwr scs8hd_decap_6
XFILLER_7_3331 vgnd vpwr scs8hd_decap_12
XFILLER_7_2685 vgnd vpwr scs8hd_decap_12
XFILLER_7_1940 vgnd vpwr scs8hd_decap_12
XFILLER_3_2538 vgnd vpwr scs8hd_decap_12
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XFILLER_1_1550 vgnd vpwr scs8hd_decap_12
XFILLER_8_3106 vgnd vpwr scs8hd_decap_12
XFILLER_8_1715 vgnd vpwr scs8hd_decap_12
XFILLER_3_4441 vgnd vpwr scs8hd_decap_12
XFILLER_6_1483 vgnd vpwr scs8hd_decap_12
XFILLER_3_3795 vgnd vpwr scs8hd_decap_12
XFILLER_2_1325 vgnd vpwr scs8hd_decap_12
XFILLER_8_4363 vgnd vpwr scs8hd_decap_12
XFILLER_6_959 vgnd vpwr scs8hd_decap_12
XFILLER_5_403 vgnd vpwr scs8hd_decap_12
XFILLER_8_2972 vgnd vpwr scs8hd_decap_12
XFILLER_7_1269 vgnd vpwr scs8hd_decap_12
XFILLER_4_4216 vgnd vpwr scs8hd_decap_12
XFILLER_4_2825 vgnd vpwr scs8hd_decap_12
XFILLER_9_4105 vgnd vpwr scs8hd_decap_12
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XFILLER_9_3404 vgnd vpwr scs8hd_decap_6
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_7_2493 vgnd vpwr scs8hd_decap_8
XFILLER_7_1770 vgnd vpwr scs8hd_decap_12
XFILLER_3_3014 vgnd vpwr scs8hd_decap_12
XFILLER_3_1623 vgnd vpwr scs8hd_decap_12
XFILLER_1_1391 vgnd vpwr scs8hd_decap_12
XFILLER_9_3993 vgnd vpwr scs8hd_decap_6
XFILLER_5_3868 vgnd vpwr scs8hd_decap_12
XFILLER_3_4271 vgnd vpwr scs8hd_decap_12
XFILLER_3_2880 vgnd vpwr scs8hd_decap_12
XFILLER_2_1166 vgnd vpwr scs8hd_decap_12
XFILLER_4_3301 vgnd vpwr scs8hd_decap_12
XFILLER_7_1099 vgnd vpwr scs8hd_decap_12
XFILLER_4_2655 vgnd vpwr scs8hd_decap_12
XFILLER_4_1910 vgnd vpwr scs8hd_decap_12
XFILLER_2_995 vgnd vpwr scs8hd_decap_12
XFILLER_9_583 vgnd vpwr scs8hd_decap_6
XFILLER_9_3256 vgnd vpwr scs8hd_decap_12
XFILLER_9_2555 vgnd vpwr scs8hd_decap_12
XFILLER_9_1854 vgnd vpwr scs8hd_decap_6
XFILLER_5_2408 vgnd vpwr scs8hd_decap_12
XFILLER_0_3721 vgnd vpwr scs8hd_decap_12
XFILLER_0_3776 vgnd vpwr scs8hd_decap_6
XFILLER_0_4477 vgnd vpwr scs8hd_decap_12
XPHY_839 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_828 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_817 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_806 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_4344 vgnd vpwr scs8hd_decap_12
XFILLER_8_2032 vgnd vpwr scs8hd_decap_12
XFILLER_8_1386 vgnd vpwr scs8hd_decap_12
XFILLER_5_2953 vgnd vpwr scs8hd_decap_12
XFILLER_4_1239 vgnd vpwr scs8hd_decap_12
XPHY_71 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_60 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_520 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_1117 vgnd vpwr scs8hd_decap_12
XFILLER_6_4119 vgnd vpwr scs8hd_decap_12
XFILLER_6_2728 vgnd vpwr scs8hd_decap_12
XFILLER_4_2496 vgnd vpwr scs8hd_decap_12
XFILLER_4_1740 vgnd vpwr scs8hd_decap_12
XFILLER_0_1637 vgnd vpwr scs8hd_decap_6
XFILLER_0_3039 vgnd vpwr scs8hd_decap_12
XFILLER_9_3020 vgnd vpwr scs8hd_decap_12
XFILLER_5_1526 vgnd vpwr scs8hd_decap_12
XFILLER_0_707 vgnd vpwr scs8hd_decap_6
XFILLER_0_4241 vgnd vpwr scs8hd_decap_6
XFILLER_2_3838 vgnd vpwr scs8hd_decap_12
XPHY_614 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_603 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_625 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1294 vgnd vpwr scs8hd_decap_12
XPHY_669 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_658 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_647 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_636 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_306 vgnd vpwr scs8hd_decap_12
XFILLER_7_4417 vgnd vpwr scs8hd_decap_12
XFILLER_5_4185 vgnd vpwr scs8hd_decap_12
XFILLER_3_501 vgnd vpwr scs8hd_decap_12
XFILLER_1_4027 vgnd vpwr scs8hd_decap_12
XFILLER_5_2794 vgnd vpwr scs8hd_decap_12
XFILLER_4_1069 vgnd vpwr scs8hd_decap_12
XFILLER_1_2636 vgnd vpwr scs8hd_decap_12
XFILLER_6_3204 vgnd vpwr scs8hd_decap_12
XFILLER_6_361 vgnd vpwr scs8hd_decap_12
XFILLER_6_2569 vgnd vpwr scs8hd_decap_12
XFILLER_6_1813 vgnd vpwr scs8hd_decap_12
XFILLER_4_2260 vgnd vpwr scs8hd_decap_12
XFILLER_4_1581 vgnd vpwr scs8hd_decap_12
XFILLER_0_1489 vgnd vpwr scs8hd_decap_12
XFILLER_0_2102 vgnd vpwr scs8hd_decap_6
XFILLER_9_2171 vgnd vpwr scs8hd_decap_12
XFILLER_6_4472 vgnd vpwr scs8hd_decap_12
XFILLER_2_4314 vgnd vpwr scs8hd_decap_12
XFILLER_9_1470 vgnd vpwr scs8hd_decap_12
XFILLER_5_1367 vgnd vpwr scs8hd_decap_12
XFILLER_0_559 vgnd vpwr scs8hd_decap_12
XFILLER_0_4093 vgnd vpwr scs8hd_decap_12
XFILLER_2_2923 vgnd vpwr scs8hd_decap_12
XFILLER_2_3679 vgnd vpwr scs8hd_decap_12
XPHY_477 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_466 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_455 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_444 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_433 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_422 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_411 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_400 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_2691 vgnd vpwr scs8hd_decap_6
XFILLER_0_3392 vgnd vpwr scs8hd_decap_12
XFILLER_7_3502 vgnd vpwr scs8hd_decap_12
XFILLER_7_147 vgnd vpwr scs8hd_decap_12
XPHY_499 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_488 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4258 vgnd vpwr scs8hd_decap_12
XFILLER_5_3270 vgnd vpwr scs8hd_decap_12
XFILLER_4_898 vgnd vpwr scs8hd_decap_12
XFILLER_3_2709 vgnd vpwr scs8hd_decap_12
XFILLER_3_342 vgnd vpwr scs8hd_decap_12
XFILLER_1_3112 vgnd vpwr scs8hd_decap_12
XFILLER_1_1721 vgnd vpwr scs8hd_decap_12
XFILLER_1_2477 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ top_width_0_height_0__pin_0_ logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[0] vgnd vpwr scs8hd_ebufn_1
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _07_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_3045 vgnd vpwr scs8hd_decap_12
XFILLER_6_1654 vgnd vpwr scs8hd_decap_12
XFILLER_3_3966 vgnd vpwr scs8hd_decap_12
XFILLER_1_4380 vgnd vpwr scs8hd_decap_12
XFILLER_0_1253 vgnd vpwr scs8hd_decap_12
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XFILLER_8_4578 vgnd vpwr scs8hd_decap_3
XFILLER_8_3899 vgnd vpwr scs8hd_decap_12
XFILLER_1_879 vgnd vpwr scs8hd_decap_12
XFILLER_0_323 vgnd vpwr scs8hd_decap_12
XFILLER_2_4155 vgnd vpwr scs8hd_decap_12
XFILLER_2_2764 vgnd vpwr scs8hd_decap_12
XFILLER_9_924 vgnd vpwr scs8hd_decap_6
XFILLER_8_434 vgnd vpwr scs8hd_decap_12
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_296 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4088 vgnd vpwr scs8hd_decap_12
XFILLER_7_3343 vgnd vpwr scs8hd_decap_12
XFILLER_7_2697 vgnd vpwr scs8hd_decap_12
XFILLER_1_1562 vgnd vpwr scs8hd_decap_12
XFILLER_8_3118 vgnd vpwr scs8hd_decap_12
XFILLER_8_1727 vgnd vpwr scs8hd_decap_12
XFILLER_6_2130 vgnd vpwr scs8hd_decap_12
XFILLER_2_1337 vgnd vpwr scs8hd_decap_12
XFILLER_8_4375 vgnd vpwr scs8hd_decap_12
XFILLER_5_415 vgnd vpwr scs8hd_decap_12
XFILLER_4_4228 vgnd vpwr scs8hd_decap_12
XFILLER_8_2984 vgnd vpwr scs8hd_decap_12
XFILLER_2_3240 vgnd vpwr scs8hd_decap_12
XFILLER_2_2594 vgnd vpwr scs8hd_decap_12
XFILLER_9_4117 vgnd vpwr scs8hd_decap_6
XFILLER_9_776 vgnd vpwr scs8hd_decap_12
XFILLER_7_3173 vgnd vpwr scs8hd_decap_12
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_3_3026 vgnd vpwr scs8hd_decap_12
XFILLER_7_1782 vgnd vpwr scs8hd_decap_12
XFILLER_3_2314 vpwr vgnd scs8hd_fill_2
XFILLER_3_1635 vgnd vpwr scs8hd_decap_12
XFILLER_0_3969 vgnd vpwr scs8hd_decap_12
XFILLER_9_3950 vgnd vpwr scs8hd_decap_12
XFILLER_8_2203 vgnd vpwr scs8hd_decap_12
XFILLER_5_4515 vgnd vpwr scs8hd_decap_12
XFILLER_8_1557 vgnd vpwr scs8hd_decap_12
XFILLER_3_4283 vgnd vpwr scs8hd_decap_12
XFILLER_3_2892 vgnd vpwr scs8hd_decap_12
XFILLER_2_1178 vgnd vpwr scs8hd_decap_12
XFILLER_8_3460 vgnd vpwr scs8hd_decap_12
XFILLER_7_1001 vgnd vpwr scs8hd_decap_12
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_4_4058 vgnd vpwr scs8hd_decap_12
XFILLER_4_3313 vgnd vpwr scs8hd_decap_12
XFILLER_1_440 vgnd vpwr scs8hd_decap_12
XFILLER_4_2667 vgnd vpwr scs8hd_decap_12
XFILLER_9_2501 vgnd vpwr scs8hd_decap_8
XFILLER_9_540 vgnd vpwr scs8hd_decap_12
XFILLER_9_3268 vgnd vpwr scs8hd_decap_12
XFILLER_9_2567 vgnd vpwr scs8hd_decap_6
XFILLER_9_2512 vgnd vpwr scs8hd_decap_12
XFILLER_9_1811 vgnd vpwr scs8hd_decap_12
XFILLER_4_4570 vgnd vpwr scs8hd_decap_8
XFILLER_3_2111 vgnd vpwr scs8hd_decap_12
XFILLER_0_4434 vgnd vpwr scs8hd_decap_12
XPHY_818 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_807 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1465 vgnd vpwr scs8hd_decap_12
XFILLER_0_3733 vgnd vpwr scs8hd_decap_12
XFILLER_0_4489 vgnd vpwr scs8hd_decap_6
XPHY_829 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_4356 vgnd vpwr scs8hd_decap_12
XFILLER_5_3600 vgnd vpwr scs8hd_decap_12
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_1398 vgnd vpwr scs8hd_decap_12
XFILLER_5_2965 vgnd vpwr scs8hd_decap_12
XFILLER_1_2807 vgnd vpwr scs8hd_decap_12
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_61 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_532 vgnd vpwr scs8hd_decap_12
XFILLER_9_1129 vgnd vpwr scs8hd_decap_12
XFILLER_4_3143 vgnd vpwr scs8hd_decap_12
XFILLER_1_281 vgnd vpwr scs8hd_decap_12
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_1752 vgnd vpwr scs8hd_decap_12
XFILLER_0_2317 vpwr vgnd scs8hd_fill_2
XFILLER_9_3032 vgnd vpwr scs8hd_decap_6
XFILLER_6_3997 vgnd vpwr scs8hd_decap_12
XFILLER_5_1538 vgnd vpwr scs8hd_decap_12
XPHY_615 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_604 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_659 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_648 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_637 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_626 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_2884 vgnd vpwr scs8hd_decap_12
XFILLER_7_4429 vgnd vpwr scs8hd_decap_12
XFILLER_7_318 vgnd vpwr scs8hd_decap_12
XFILLER_5_4197 vgnd vpwr scs8hd_decap_12
XFILLER_5_3441 vgnd vpwr scs8hd_decap_12
XFILLER_3_513 vgnd vpwr scs8hd_decap_12
XFILLER_1_4039 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_2648 vgnd vpwr scs8hd_decap_12
XFILLER_6_3216 vgnd vpwr scs8hd_decap_12
XFILLER_7_830 vgnd vpwr scs8hd_decap_12
XFILLER_6_373 vgnd vpwr scs8hd_decap_12
XFILLER_6_1825 vgnd vpwr scs8hd_decap_12
XFILLER_4_2272 vgnd vpwr scs8hd_decap_12
XFILLER_1_4551 vgnd vpwr scs8hd_decap_12
XFILLER_4_1593 vgnd vpwr scs8hd_decap_12
XFILLER_9_2183 vgnd vpwr scs8hd_decap_12
XFILLER_5_2014 vgnd vpwr scs8hd_decap_12
XFILLER_2_4326 vgnd vpwr scs8hd_decap_12
XFILLER_9_1482 vgnd vpwr scs8hd_decap_6
XFILLER_5_1379 vgnd vpwr scs8hd_decap_12
XFILLER_2_2935 vgnd vpwr scs8hd_decap_12
XFILLER_8_605 vgnd vpwr scs8hd_decap_12
XPHY_489 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_478 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_467 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_456 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_445 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_434 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_423 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_412 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_401 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3514 vgnd vpwr scs8hd_decap_12
XFILLER_7_159 vgnd vpwr scs8hd_decap_12
XFILLER_4_800 vgnd vpwr scs8hd_decap_12
XFILLER_3_354 vgnd vpwr scs8hd_decap_12
XFILLER_7_2868 vgnd vpwr scs8hd_decap_12
XFILLER_5_3282 vgnd vpwr scs8hd_decap_12
XFILLER_1_3124 vgnd vpwr scs8hd_decap_12
XFILLER_1_1733 vgnd vpwr scs8hd_decap_12
XFILLER_1_2489 vgnd vpwr scs8hd_decap_12
XFILLER_6_3057 vgnd vpwr scs8hd_decap_12
XFILLER_6_2301 vgnd vpwr scs8hd_decap_12
XFILLER_6_1666 vgnd vpwr scs8hd_decap_12
XFILLER_3_3978 vgnd vpwr scs8hd_decap_12
XFILLER_0_1210 vgnd vpwr scs8hd_decap_12
XFILLER_2_1508 vgnd vpwr scs8hd_decap_12
XFILLER_0_1265 vgnd vpwr scs8hd_decap_6
XFILLER_1_2990 vgnd vpwr scs8hd_decap_12
XFILLER_8_4546 vgnd vpwr scs8hd_decap_12
XFILLER_8_3801 vgnd vpwr scs8hd_decap_12
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_0_335 vgnd vpwr scs8hd_decap_6
XFILLER_2_3411 vgnd vpwr scs8hd_decap_12
XFILLER_2_4167 vgnd vpwr scs8hd_decap_12
XFILLER_8_446 vgnd vpwr scs8hd_decap_12
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_286 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_297 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3609 vgnd vpwr scs8hd_decap_12
XFILLER_9_2908 vgnd vpwr scs8hd_decap_6
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XFILLER_7_1953 vgnd vpwr scs8hd_decap_12
XFILLER_3_1806 vgnd vpwr scs8hd_decap_12
XFILLER_1_1574 vgnd vpwr scs8hd_decap_12
XFILLER_1_2286 vgnd vpwr scs8hd_fill_1
XFILLER_8_991 vgnd vpwr scs8hd_decap_12
XFILLER_6_2142 vgnd vpwr scs8hd_decap_12
XFILLER_3_4454 vgnd vpwr scs8hd_decap_12
XFILLER_6_1496 vgnd vpwr scs8hd_decap_12
XFILLER_2_1349 vgnd vpwr scs8hd_decap_12
XFILLER_8_4387 vgnd vpwr scs8hd_decap_12
XFILLER_8_3631 vgnd vpwr scs8hd_decap_12
XFILLER_1_611 vgnd vpwr scs8hd_decap_12
XFILLER_8_2996 vgnd vpwr scs8hd_decap_12
XFILLER_4_2838 vgnd vpwr scs8hd_decap_12
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_2_3252 vgnd vpwr scs8hd_decap_12
XFILLER_9_788 vgnd vpwr scs8hd_decap_12
XFILLER_8_276 vgnd vpwr scs8hd_decap_12
XFILLER_7_3185 vgnd vpwr scs8hd_decap_12
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_4_471 vgnd vpwr scs8hd_decap_12
XFILLER_3_3038 vgnd vpwr scs8hd_decap_12
XFILLER_7_1794 vgnd vpwr scs8hd_decap_12
XFILLER_3_2359 vpwr vgnd scs8hd_fill_2
XFILLER_3_2348 vpwr vgnd scs8hd_fill_2
XFILLER_1_2050 vgnd vpwr scs8hd_decap_12
XFILLER_9_3962 vgnd vpwr scs8hd_decap_6
XFILLER_8_2215 vgnd vpwr scs8hd_decap_12
XFILLER_5_4527 vgnd vpwr scs8hd_decap_12
XFILLER_8_1569 vgnd vpwr scs8hd_decap_12
XFILLER_3_4295 vgnd vpwr scs8hd_decap_12
XFILLER_6_703 vgnd vpwr scs8hd_decap_12
XFILLER_8_3472 vgnd vpwr scs8hd_decap_12
XFILLER_7_1013 vgnd vpwr scs8hd_decap_12
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_1_452 vgnd vpwr scs8hd_decap_12
XFILLER_4_2679 vgnd vpwr scs8hd_decap_12
XFILLER_4_1923 vgnd vpwr scs8hd_decap_12
XFILLER_2_3082 vgnd vpwr scs8hd_decap_12
XFILLER_9_552 vgnd vpwr scs8hd_decap_6
XFILLER_2_1691 vgnd vpwr scs8hd_decap_12
XFILLER_9_3225 vgnd vpwr scs8hd_decap_12
XFILLER_9_2524 vgnd vpwr scs8hd_decap_12
XFILLER_9_1823 vgnd vpwr scs8hd_decap_6
XFILLER_7_2270 vgnd vpwr scs8hd_decap_12
XFILLER_5_1709 vgnd vpwr scs8hd_decap_12
XFILLER_3_2123 vgnd vpwr scs8hd_decap_12
XFILLER_0_3745 vgnd vpwr scs8hd_decap_6
XFILLER_0_4446 vgnd vpwr scs8hd_decap_12
XPHY_819 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_808 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1477 vgnd vpwr scs8hd_decap_12
XFILLER_8_2045 vgnd vpwr scs8hd_decap_12
XFILLER_8_1300 vgnd vpwr scs8hd_decap_12
XFILLER_5_4368 vgnd vpwr scs8hd_decap_12
XFILLER_5_3612 vgnd vpwr scs8hd_decap_12
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_2977 vgnd vpwr scs8hd_decap_12
XFILLER_3_3380 vgnd vpwr scs8hd_decap_12
XFILLER_1_2819 vgnd vpwr scs8hd_decap_12
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_62 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_51 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_544 vgnd vpwr scs8hd_decap_12
XFILLER_4_3155 vgnd vpwr scs8hd_decap_12
XFILLER_1_293 vgnd vpwr scs8hd_decap_12
XFILLER_0_3008 vgnd vpwr scs8hd_decap_12
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_4_1764 vgnd vpwr scs8hd_decap_12
XFILLER_0_1606 vgnd vpwr scs8hd_decap_6
XFILLER_9_1675 vgnd vpwr scs8hd_decap_12
XFILLER_0_3597 vgnd vpwr scs8hd_decap_12
XFILLER_0_4210 vgnd vpwr scs8hd_decap_6
XPHY_616 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_605 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_649 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_638 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_627 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_2896 vgnd vpwr scs8hd_decap_12
XFILLER_3_525 vgnd vpwr scs8hd_decap_12
XFILLER_8_1130 vgnd vpwr scs8hd_decap_12
XFILLER_5_3453 vgnd vpwr scs8hd_decap_12
XFILLER_1_1904 vgnd vpwr scs8hd_decap_12
XFILLER_7_842 vgnd vpwr scs8hd_decap_12
XFILLER_6_3228 vgnd vpwr scs8hd_decap_12
XFILLER_6_385 vgnd vpwr scs8hd_decap_12
XFILLER_6_1837 vgnd vpwr scs8hd_decap_12
XFILLER_4_2284 vgnd vpwr scs8hd_decap_4
XFILLER_4_2240 vgnd vpwr scs8hd_decap_12
XFILLER_1_4563 vgnd vpwr scs8hd_decap_12
XFILLER_0_1458 vgnd vpwr scs8hd_decap_12
XFILLER_9_2195 vgnd vpwr scs8hd_decap_6
XFILLER_9_2140 vgnd vpwr scs8hd_decap_12
XFILLER_6_4485 vgnd vpwr scs8hd_decap_12
XFILLER_6_3740 vgnd vpwr scs8hd_decap_12
XFILLER_5_2026 vgnd vpwr scs8hd_decap_12
XFILLER_2_4338 vgnd vpwr scs8hd_decap_12
XFILLER_0_528 vgnd vpwr scs8hd_decap_12
XFILLER_0_2660 vgnd vpwr scs8hd_decap_6
XFILLER_0_4062 vgnd vpwr scs8hd_decap_12
XFILLER_2_2947 vgnd vpwr scs8hd_decap_12
XFILLER_8_617 vgnd vpwr scs8hd_decap_12
XPHY_479 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_468 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_457 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_446 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_435 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_424 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_413 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_402 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3526 vgnd vpwr scs8hd_decap_12
XFILLER_4_812 vgnd vpwr scs8hd_decap_12
XFILLER_1_3136 vgnd vpwr scs8hd_decap_12
XFILLER_5_1892 vgnd vpwr scs8hd_decap_12
XFILLER_1_1745 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XFILLER_7_672 vgnd vpwr scs8hd_decap_12
XFILLER_6_3069 vgnd vpwr scs8hd_decap_12
XFILLER_6_2346 vgnd vpwr scs8hd_decap_3
XFILLER_6_2335 vgnd vpwr scs8hd_decap_8
XFILLER_6_2313 vgnd vpwr scs8hd_decap_12
X_19_ gfpga_pad_GPIO_PAD[0] top_width_0_height_0__pin_1_ vgnd vpwr scs8hd_buf_2
XFILLER_4_2081 vgnd vpwr scs8hd_decap_12
XFILLER_0_1222 vgnd vpwr scs8hd_decap_12
XFILLER_1_4393 vgnd vpwr scs8hd_decap_12
XFILLER_8_4558 vgnd vpwr scs8hd_decap_12
XFILLER_6_3570 vgnd vpwr scs8hd_decap_12
XFILLER_5_1111 vgnd vpwr scs8hd_decap_12
XFILLER_2_3423 vgnd vpwr scs8hd_decap_12
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_2777 vgnd vpwr scs8hd_decap_12
XFILLER_7_4002 vgnd vpwr scs8hd_decap_12
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_287 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_298 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3356 vgnd vpwr scs8hd_decap_12
XFILLER_7_2611 vgnd vpwr scs8hd_decap_12
XFILLER_4_642 vgnd vpwr scs8hd_decap_12
XFILLER_3_3209 vgnd vpwr scs8hd_decap_12
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XFILLER_7_1965 vgnd vpwr scs8hd_decap_12
XFILLER_3_1818 vgnd vpwr scs8hd_decap_12
XFILLER_0_881 vgnd vpwr scs8hd_decap_12
XFILLER_1_2221 vgnd vpwr scs8hd_decap_12
XFILLER_7_4580 vgnd vpwr scs8hd_fill_1
XFILLER_6_2154 vgnd vpwr scs8hd_decap_12
XFILLER_3_4466 vgnd vpwr scs8hd_decap_12
XFILLER_5_428 vgnd vpwr scs8hd_decap_12
XFILLER_8_4399 vgnd vpwr scs8hd_decap_12
XFILLER_8_3643 vgnd vpwr scs8hd_decap_12
XFILLER_1_623 vgnd vpwr scs8hd_decap_12
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_9_745 vgnd vpwr scs8hd_decap_12
XFILLER_2_1862 vgnd vpwr scs8hd_decap_12
XFILLER_8_288 vgnd vpwr scs8hd_decap_12
XFILLER_5_940 vgnd vpwr scs8hd_decap_12
XFILLER_7_3197 vgnd vpwr scs8hd_decap_12
XFILLER_7_2441 vpwr vgnd scs8hd_fill_2
XFILLER_4_483 vgnd vpwr scs8hd_decap_12
XFILLER_3_2327 vpwr vgnd scs8hd_fill_2
XFILLER_0_3938 vgnd vpwr scs8hd_decap_12
XFILLER_3_1648 vgnd vpwr scs8hd_decap_12
XFILLER_1_2062 vgnd vpwr scs8hd_decap_12
XFILLER_5_4539 vgnd vpwr scs8hd_decap_12
XFILLER_3_3551 vgnd vpwr scs8hd_decap_12
XFILLER_6_715 vgnd vpwr scs8hd_decap_12
XFILLER_5_269 vgnd vpwr scs8hd_decap_12
XFILLER_8_3484 vgnd vpwr scs8hd_decap_12
XFILLER_7_1025 vgnd vpwr scs8hd_decap_12
XFILLER_4_3326 vgnd vpwr scs8hd_decap_12
XFILLER_1_464 vgnd vpwr scs8hd_decap_12
XFILLER_2_910 vgnd vpwr scs8hd_decap_12
XFILLER_4_1935 vgnd vpwr scs8hd_decap_12
XFILLER_2_2371 vgnd vpwr scs8hd_decap_4
XFILLER_2_3094 vgnd vpwr scs8hd_decap_12
XFILLER_9_3237 vgnd vpwr scs8hd_decap_12
XFILLER_9_2536 vgnd vpwr scs8hd_decap_6
XFILLER_5_781 vgnd vpwr scs8hd_decap_12
XFILLER_7_2282 vgnd vpwr scs8hd_decap_12
XFILLER_0_3702 vgnd vpwr scs8hd_decap_12
XFILLER_0_4403 vgnd vpwr scs8hd_decap_12
XFILLER_0_4458 vgnd vpwr scs8hd_decap_6
XPHY_809 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1489 vgnd vpwr scs8hd_decap_12
XFILLER_8_2057 vgnd vpwr scs8hd_decap_12
XFILLER_5_3624 vgnd vpwr scs8hd_decap_12
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XFILLER_3_3392 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_63 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_52 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_556 vgnd vpwr scs8hd_decap_12
XFILLER_2_751 vgnd vpwr scs8hd_decap_12
XFILLER_4_3167 vgnd vpwr scs8hd_decap_12
XFILLER_4_2411 vgnd vpwr scs8hd_decap_12
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_4_1776 vgnd vpwr scs8hd_decap_12
XFILLER_9_3001 vgnd vpwr scs8hd_decap_6
XFILLER_9_2388 vgnd vpwr scs8hd_decap_12
XFILLER_6_3911 vgnd vpwr scs8hd_decap_12
XFILLER_2_4509 vgnd vpwr scs8hd_decap_12
XFILLER_9_1687 vgnd vpwr scs8hd_decap_12
XFILLER_0_2853 vgnd vpwr scs8hd_decap_12
XPHY_606 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_639 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_628 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_617 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_4291 vgnd vpwr scs8hd_decap_12
XFILLER_5_4100 vgnd vpwr scs8hd_decap_12
XFILLER_3_537 vgnd vpwr scs8hd_decap_12
XFILLER_9_3590 vgnd vpwr scs8hd_decap_6
XFILLER_8_1142 vgnd vpwr scs8hd_decap_12
XFILLER_5_3465 vgnd vpwr scs8hd_decap_12
XFILLER_1_3307 vgnd vpwr scs8hd_decap_12
XFILLER_1_1916 vgnd vpwr scs8hd_decap_12
XFILLER_2_581 vgnd vpwr scs8hd_decap_12
XFILLER_6_1849 vgnd vpwr scs8hd_decap_12
XFILLER_4_2252 vgnd vpwr scs8hd_decap_6
XFILLER_9_180 vgnd vpwr scs8hd_decap_6
XFILLER_9_2152 vgnd vpwr scs8hd_decap_12
XFILLER_9_1451 vgnd vpwr scs8hd_decap_6
XFILLER_6_4497 vgnd vpwr scs8hd_decap_12
XFILLER_5_2038 vgnd vpwr scs8hd_decap_12
XFILLER_0_4074 vgnd vpwr scs8hd_decap_12
XPHY_425 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_414 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_403 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1050 vgnd vpwr scs8hd_decap_12
XFILLER_8_629 vgnd vpwr scs8hd_decap_12
XPHY_469 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_458 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_447 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_436 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_367 vgnd vpwr scs8hd_decap_12
XFILLER_5_3295 vgnd vpwr scs8hd_decap_12
XFILLER_5_2550 vgnd vpwr scs8hd_decap_12
XFILLER_1_2403 vgnd vpwr scs8hd_decap_12
XFILLER_1_3148 vgnd vpwr scs8hd_decap_12
XFILLER_1_1757 vgnd vpwr scs8hd_decap_12
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_7_684 vgnd vpwr scs8hd_decap_12
XFILLER_6_2358 vgnd vpwr scs8hd_decap_12
XFILLER_6_2325 vgnd vpwr scs8hd_fill_1
X_18_ gfpga_pad_GPIO_PAD[7] top_width_0_height_0__pin_15_ vgnd vpwr scs8hd_buf_2
XFILLER_6_1679 vgnd vpwr scs8hd_decap_12
XFILLER_4_2093 vgnd vpwr scs8hd_decap_12
XFILLER_0_1234 vgnd vpwr scs8hd_decap_6
XFILLER_8_3814 vgnd vpwr scs8hd_decap_12
XFILLER_0_304 vgnd vpwr scs8hd_decap_6
XFILLER_6_3582 vgnd vpwr scs8hd_decap_12
XFILLER_5_1123 vgnd vpwr scs8hd_decap_12
XFILLER_2_2789 vgnd vpwr scs8hd_decap_12
XFILLER_2_3435 vgnd vpwr scs8hd_decap_12
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_459 vgnd vpwr scs8hd_decap_12
XFILLER_7_4014 vgnd vpwr scs8hd_decap_12
XPHY_288 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_299 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3368 vgnd vpwr scs8hd_decap_12
XFILLER_4_654 vgnd vpwr scs8hd_decap_12
XFILLER_0_893 vgnd vpwr scs8hd_decap_6
XFILLER_7_1977 vgnd vpwr scs8hd_decap_12
XFILLER_5_2380 vgnd vpwr scs8hd_decap_3
XFILLER_1_1587 vgnd vpwr scs8hd_decap_12
XFILLER_1_2233 vgnd vpwr scs8hd_decap_12
XFILLER_7_3880 vgnd vpwr scs8hd_decap_12
XFILLER_6_1410 vgnd vpwr scs8hd_decap_12
XFILLER_3_4478 vgnd vpwr scs8hd_decap_12
XFILLER_3_3722 vgnd vpwr scs8hd_decap_12
XFILLER_2_2008 vgnd vpwr scs8hd_decap_12
XFILLER_0_1086 vgnd vpwr scs8hd_decap_12
XFILLER_1_3490 vgnd vpwr scs8hd_decap_12
XFILLER_8_3655 vgnd vpwr scs8hd_decap_12
XFILLER_1_635 vgnd vpwr scs8hd_decap_12
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_2_1874 vgnd vpwr scs8hd_decap_12
XFILLER_2_2520 vgnd vpwr scs8hd_decap_12
XFILLER_2_3265 vgnd vpwr scs8hd_decap_12
XFILLER_9_757 vgnd vpwr scs8hd_decap_12
XFILLER_9_2729 vgnd vpwr scs8hd_decap_12
XFILLER_5_952 vgnd vpwr scs8hd_decap_12
XFILLER_4_495 vgnd vpwr scs8hd_decap_12
XFILLER_9_3931 vgnd vpwr scs8hd_decap_6
XFILLER_8_2228 vgnd vpwr scs8hd_decap_12
XFILLER_3_3563 vgnd vpwr scs8hd_decap_12
XFILLER_8_4131 vgnd vpwr scs8hd_decap_12
XFILLER_6_727 vgnd vpwr scs8hd_decap_12
XFILLER_2_922 vgnd vpwr scs8hd_decap_12
XFILLER_8_3496 vgnd vpwr scs8hd_decap_12
XFILLER_8_2740 vgnd vpwr scs8hd_decap_12
XFILLER_4_3338 vgnd vpwr scs8hd_decap_12
XFILLER_1_476 vgnd vpwr scs8hd_decap_12
XFILLER_4_1947 vgnd vpwr scs8hd_decap_12
XFILLER_9_521 vgnd vpwr scs8hd_decap_6
XFILLER_9_3249 vgnd vpwr scs8hd_decap_6
XFILLER_0_4415 vgnd vpwr scs8hd_decap_12
XFILLER_7_2294 vgnd vpwr scs8hd_decap_12
XFILLER_4_3850 vgnd vpwr scs8hd_decap_12
XFILLER_3_2136 vgnd vpwr scs8hd_decap_12
XFILLER_0_3714 vgnd vpwr scs8hd_decap_6
XFILLER_3_708 vgnd vpwr scs8hd_decap_12
XFILLER_9_3783 vgnd vpwr scs8hd_decap_12
XFILLER_8_2069 vgnd vpwr scs8hd_decap_12
XFILLER_8_1313 vgnd vpwr scs8hd_decap_12
XFILLER_5_3636 vgnd vpwr scs8hd_decap_12
XFILLER_6_1081 vgnd vpwr scs8hd_decap_12
XPHY_64 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_53 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_42 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_20 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_31 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_568 vgnd vpwr scs8hd_decap_12
XFILLER_8_2581 vgnd vpwr scs8hd_decap_12
XFILLER_4_3179 vgnd vpwr scs8hd_decap_12
XFILLER_4_1788 vgnd vpwr scs8hd_decap_12
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_2_2191 vgnd vpwr scs8hd_decap_12
XFILLER_9_373 vgnd vpwr scs8hd_decap_12
XFILLER_9_1699 vgnd vpwr scs8hd_decap_6
XFILLER_9_1644 vgnd vpwr scs8hd_decap_12
XFILLER_6_3923 vgnd vpwr scs8hd_decap_12
XFILLER_5_2209 vgnd vpwr scs8hd_decap_12
XPHY_607 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1221 vgnd vpwr scs8hd_decap_12
XFILLER_0_2865 vgnd vpwr scs8hd_decap_12
XFILLER_0_3566 vgnd vpwr scs8hd_decap_12
XPHY_629 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_618 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3709 vgnd vpwr scs8hd_decap_12
XFILLER_5_4112 vgnd vpwr scs8hd_decap_12
XFILLER_8_1154 vgnd vpwr scs8hd_decap_12
XFILLER_5_2721 vgnd vpwr scs8hd_decap_12
XFILLER_1_3319 vgnd vpwr scs8hd_decap_12
XFILLER_1_1928 vgnd vpwr scs8hd_decap_12
XFILLER_7_855 vgnd vpwr scs8hd_decap_12
XFILLER_6_398 vgnd vpwr scs8hd_decap_12
XFILLER_2_593 vgnd vpwr scs8hd_decap_12
XFILLER_4_2297 vgnd vpwr scs8hd_decap_4
XFILLER_0_1427 vgnd vpwr scs8hd_decap_12
XFILLER_1_3831 vgnd vpwr scs8hd_decap_12
XFILLER_1_4576 vgnd vpwr scs8hd_decap_4
XFILLER_9_2164 vgnd vpwr scs8hd_decap_6
XFILLER_6_3753 vgnd vpwr scs8hd_decap_12
XFILLER_0_3330 vgnd vpwr scs8hd_decap_12
XFILLER_0_4031 vgnd vpwr scs8hd_decap_12
XFILLER_0_4086 vgnd vpwr scs8hd_decap_6
XFILLER_2_3606 vgnd vpwr scs8hd_decap_12
XPHY_459 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_448 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_437 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_426 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_415 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_404 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1062 vgnd vpwr scs8hd_decap_12
XFILLER_4_825 vgnd vpwr scs8hd_decap_12
XFILLER_7_3539 vgnd vpwr scs8hd_decap_12
XFILLER_3_379 vgnd vpwr scs8hd_decap_12
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_2415 vgnd vpwr scs8hd_decap_12
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
XFILLER_7_696 vgnd vpwr scs8hd_decap_12
XFILLER_3_891 vgnd vpwr scs8hd_decap_12
XFILLER_1_3661 vgnd vpwr scs8hd_decap_12
X_17_ gfpga_pad_GPIO_PAD[6] top_width_0_height_0__pin_13_ vgnd vpwr scs8hd_buf_2
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_3826 vgnd vpwr scs8hd_decap_12
XFILLER_1_806 vgnd vpwr scs8hd_decap_12
XFILLER_6_3594 vgnd vpwr scs8hd_decap_12
XFILLER_5_1135 vgnd vpwr scs8hd_decap_12
XFILLER_0_1780 vgnd vpwr scs8hd_decap_12
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_2481 vgnd vpwr scs8hd_decap_12
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_289 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_666 vgnd vpwr scs8hd_decap_12
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
XFILLER_7_2624 vgnd vpwr scs8hd_decap_12
XFILLER_7_1989 vgnd vpwr scs8hd_decap_12
XFILLER_0_850 vgnd vpwr scs8hd_decap_12
XFILLER_1_1599 vgnd vpwr scs8hd_decap_12
XFILLER_1_2245 vgnd vpwr scs8hd_decap_12
XFILLER_1_2289 vpwr vgnd scs8hd_fill_2
XPHY_790 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xlogical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _09_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_3892 vgnd vpwr scs8hd_decap_12
XFILLER_6_2167 vgnd vpwr scs8hd_decap_12
XFILLER_6_1422 vgnd vpwr scs8hd_decap_12
XFILLER_3_3734 vgnd vpwr scs8hd_decap_12
XFILLER_0_1098 vgnd vpwr scs8hd_decap_12
XFILLER_8_4302 vgnd vpwr scs8hd_decap_12
XFILLER_8_3667 vgnd vpwr scs8hd_decap_12
XFILLER_8_2911 vgnd vpwr scs8hd_decap_12
XFILLER_6_4070 vgnd vpwr scs8hd_decap_12
XFILLER_7_1208 vgnd vpwr scs8hd_decap_12
XFILLER_4_3509 vgnd vpwr scs8hd_decap_12
XFILLER_1_647 vgnd vpwr scs8hd_decap_12
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XFILLER_2_1886 vgnd vpwr scs8hd_decap_12
XFILLER_2_3277 vgnd vpwr scs8hd_decap_12
XFILLER_9_769 vgnd vpwr scs8hd_decap_6
XFILLER_9_714 vgnd vpwr scs8hd_decap_12
XFILLER_8_202 vgnd vpwr scs8hd_decap_12
XFILLER_5_997 vgnd vpwr scs8hd_decap_3
XFILLER_5_964 vgnd vpwr scs8hd_decap_12
XFILLER_0_3907 vgnd vpwr scs8hd_decap_12
XFILLER_1_1330 vgnd vpwr scs8hd_decap_12
XFILLER_1_2075 vgnd vpwr scs8hd_decap_12
XFILLER_5_3807 vgnd vpwr scs8hd_decap_12
XFILLER_3_4210 vgnd vpwr scs8hd_decap_12
XFILLER_6_1252 vgnd vpwr scs8hd_decap_12
XFILLER_3_3575 vgnd vpwr scs8hd_decap_12
XFILLER_2_1105 vgnd vpwr scs8hd_decap_12
XFILLER_8_4143 vgnd vpwr scs8hd_decap_12
XFILLER_6_739 vgnd vpwr scs8hd_decap_12
XFILLER_2_934 vgnd vpwr scs8hd_decap_12
XFILLER_8_2752 vgnd vpwr scs8hd_decap_12
XFILLER_7_1038 vgnd vpwr scs8hd_decap_12
XFILLER_4_1959 vgnd vpwr scs8hd_decap_12
XFILLER_2_2340 vpwr vgnd scs8hd_fill_2
XFILLER_9_3206 vgnd vpwr scs8hd_decap_12
XFILLER_5_794 vgnd vpwr scs8hd_decap_12
XFILLER_4_3862 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ top_width_0_height_0__pin_2_ logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[1] vgnd vpwr scs8hd_ebufn_1
XFILLER_0_4427 vgnd vpwr scs8hd_decap_6
XFILLER_7_1550 vgnd vpwr scs8hd_decap_12
XFILLER_3_2148 vgnd vpwr scs8hd_decap_12
XFILLER_1_1160 vgnd vpwr scs8hd_decap_12
XFILLER_9_4496 vgnd vpwr scs8hd_decap_12
XFILLER_9_3795 vgnd vpwr scs8hd_decap_12
XFILLER_8_1325 vgnd vpwr scs8hd_decap_12
XFILLER_5_3648 vgnd vpwr scs8hd_decap_12
XFILLER_3_4051 vgnd vpwr scs8hd_decap_12
XFILLER_3_2660 vgnd vpwr scs8hd_decap_12
XFILLER_6_1093 vgnd vpwr scs8hd_decap_12
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_54 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_43 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_32 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_764 vgnd vpwr scs8hd_decap_12
XFILLER_9_385 vgnd vpwr scs8hd_decap_12
XFILLER_9_2357 vgnd vpwr scs8hd_decap_12
XFILLER_9_1656 vgnd vpwr scs8hd_decap_12
XFILLER_4_3692 vgnd vpwr scs8hd_decap_12
XFILLER_0_4279 vgnd vpwr scs8hd_decap_12
XPHY_608 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_1391 vgnd vpwr scs8hd_decap_12
XPHY_619 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1233 vgnd vpwr scs8hd_decap_12
XFILLER_0_2822 vgnd vpwr scs8hd_decap_12
XFILLER_0_2877 vgnd vpwr scs8hd_decap_6
XFILLER_0_3578 vgnd vpwr scs8hd_decap_12
XFILLER_9_4260 vgnd vpwr scs8hd_decap_12
XFILLER_5_4124 vgnd vpwr scs8hd_decap_12
XFILLER_8_1166 vgnd vpwr scs8hd_decap_12
XFILLER_5_3478 vgnd vpwr scs8hd_decap_12
XFILLER_5_2733 vgnd vpwr scs8hd_decap_12
XFILLER_4_1008 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _14_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_867 vgnd vpwr scs8hd_decap_12
XFILLER_6_300 vgnd vpwr scs8hd_decap_12
XFILLER_6_2508 vgnd vpwr scs8hd_decap_12
XFILLER_5_3990 vgnd vpwr scs8hd_decap_12
XFILLER_4_1520 vgnd vpwr scs8hd_decap_12
XFILLER_0_1439 vgnd vpwr scs8hd_decap_12
XFILLER_9_2121 vgnd vpwr scs8hd_decap_12
XFILLER_9_1420 vgnd vpwr scs8hd_decap_6
XFILLER_6_4411 vgnd vpwr scs8hd_decap_12
XFILLER_6_3765 vgnd vpwr scs8hd_decap_12
XFILLER_0_509 vgnd vpwr scs8hd_decap_12
XFILLER_5_1306 vgnd vpwr scs8hd_decap_12
XFILLER_0_4043 vgnd vpwr scs8hd_decap_12
XFILLER_2_3618 vgnd vpwr scs8hd_decap_12
XPHY_449 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_438 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_427 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_416 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_405 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1074 vgnd vpwr scs8hd_decap_12
XFILLER_4_837 vgnd vpwr scs8hd_decap_12
XFILLER_5_2563 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ top_width_0_height_0__pin_12_ vgnd vpwr scs8hd_diode_2
XFILLER_1_2427 vgnd vpwr scs8hd_decap_12
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
XFILLER_3_3905 vgnd vpwr scs8hd_decap_12
X_16_ gfpga_pad_GPIO_PAD[5] top_width_0_height_0__pin_11_ vgnd vpwr scs8hd_buf_2
XFILLER_4_1361 vgnd vpwr scs8hd_decap_12
XFILLER_0_1203 vgnd vpwr scs8hd_decap_6
XFILLER_1_3673 vgnd vpwr scs8hd_decap_12
XFILLER_9_1272 vgnd vpwr scs8hd_decap_12
XFILLER_8_3838 vgnd vpwr scs8hd_decap_12
XFILLER_6_4241 vgnd vpwr scs8hd_decap_12
XFILLER_6_2850 vgnd vpwr scs8hd_decap_12
XFILLER_1_818 vgnd vpwr scs8hd_decap_12
XFILLER_2_2703 vgnd vpwr scs8hd_decap_12
XFILLER_2_3448 vgnd vpwr scs8hd_decap_12
XFILLER_5_1147 vgnd vpwr scs8hd_decap_12
XFILLER_0_2493 vgnd vpwr scs8hd_decap_12
XFILLER_0_3194 vgnd vpwr scs8hd_decap_12
XFILLER_0_1792 vgnd vpwr scs8hd_decap_6
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4027 vgnd vpwr scs8hd_decap_12
XFILLER_4_678 vgnd vpwr scs8hd_decap_12
XFILLER_7_2636 vgnd vpwr scs8hd_decap_12
XFILLER_1_1501 vgnd vpwr scs8hd_decap_12
XFILLER_0_862 vgnd vpwr scs8hd_decap_6
XFILLER_2_3960 vgnd vpwr scs8hd_decap_12
XPHY_791 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_780 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_3746 vgnd vpwr scs8hd_decap_12
XFILLER_6_2179 vgnd vpwr scs8hd_decap_12
XFILLER_4_1191 vgnd vpwr scs8hd_decap_12
XFILLER_0_1055 vgnd vpwr scs8hd_decap_12
XFILLER_8_4314 vgnd vpwr scs8hd_decap_12
XFILLER_8_2923 vgnd vpwr scs8hd_decap_12
XFILLER_8_3679 vgnd vpwr scs8hd_decap_12
XFILLER_6_4082 vgnd vpwr scs8hd_decap_12
XFILLER_6_2691 vgnd vpwr scs8hd_decap_12
XFILLER_1_659 vgnd vpwr scs8hd_decap_12
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_2_2533 vgnd vpwr scs8hd_decap_12
XFILLER_2_3289 vgnd vpwr scs8hd_decap_12
XFILLER_0_2290 vpwr vgnd scs8hd_fill_2
XFILLER_2_1898 vgnd vpwr scs8hd_decap_12
XFILLER_9_726 vgnd vpwr scs8hd_decap_12
XFILLER_7_3112 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_1721 vgnd vpwr scs8hd_decap_12
XFILLER_3_2319 vpwr vgnd scs8hd_fill_2
XFILLER_1_2087 vgnd vpwr scs8hd_decap_12
XFILLER_0_3919 vgnd vpwr scs8hd_decap_12
XFILLER_9_3900 vgnd vpwr scs8hd_decap_6
XFILLER_7_4380 vgnd vpwr scs8hd_decap_12
XFILLER_6_1264 vgnd vpwr scs8hd_decap_12
XFILLER_5_3819 vgnd vpwr scs8hd_decap_12
XFILLER_3_4222 vgnd vpwr scs8hd_decap_12
XFILLER_3_3587 vgnd vpwr scs8hd_decap_12
XFILLER_3_2831 vgnd vpwr scs8hd_decap_12
XFILLER_2_1117 vgnd vpwr scs8hd_decap_12
XFILLER_8_4155 vgnd vpwr scs8hd_decap_12
XFILLER_8_2764 vgnd vpwr scs8hd_decap_12
XFILLER_4_2606 vgnd vpwr scs8hd_decap_12
XFILLER_1_489 vgnd vpwr scs8hd_decap_12
XFILLER_9_3218 vgnd vpwr scs8hd_decap_6
Xlogical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _15_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_1562 vgnd vpwr scs8hd_decap_12
XFILLER_3_1404 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ top_width_0_height_0__pin_8_ vgnd vpwr scs8hd_diode_2
XFILLER_1_1172 vgnd vpwr scs8hd_decap_12
XFILLER_9_3752 vgnd vpwr scs8hd_decap_12
XFILLER_5_2904 vgnd vpwr scs8hd_decap_12
XFILLER_8_1337 vgnd vpwr scs8hd_decap_12
XFILLER_3_4063 vgnd vpwr scs8hd_decap_12
XFILLER_3_2672 vgnd vpwr scs8hd_decap_12
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_55 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_44 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_33 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_3240 vgnd vpwr scs8hd_decap_12
XFILLER_8_2594 vgnd vpwr scs8hd_decap_12
XFILLER_4_2425 vgnd vpwr scs8hd_decap_12
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_776 vgnd vpwr scs8hd_decap_12
XFILLER_4_2469 vpwr vgnd scs8hd_fill_2
XFILLER_9_342 vgnd vpwr scs8hd_decap_12
XFILLER_9_2369 vgnd vpwr scs8hd_decap_12
XFILLER_9_1613 vgnd vpwr scs8hd_decap_12
XFILLER_9_397 vgnd vpwr scs8hd_decap_6
XFILLER_6_3936 vgnd vpwr scs8hd_decap_12
XFILLER_9_1668 vgnd vpwr scs8hd_decap_6
XFILLER_4_4350 vgnd vpwr scs8hd_decap_12
XFILLER_3_1245 vgnd vpwr scs8hd_decap_12
XFILLER_0_2834 vgnd vpwr scs8hd_decap_12
XFILLER_0_3535 vgnd vpwr scs8hd_decap_12
XPHY_609 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_4272 vgnd vpwr scs8hd_decap_6
XFILLER_5_4136 vgnd vpwr scs8hd_decap_12
XFILLER_8_1178 vgnd vpwr scs8hd_decap_12
XFILLER_7_879 vgnd vpwr scs8hd_decap_12
XFILLER_6_312 vgnd vpwr scs8hd_decap_12
XFILLER_4_1532 vgnd vpwr scs8hd_decap_12
XFILLER_1_3844 vgnd vpwr scs8hd_decap_12
XFILLER_9_2133 vgnd vpwr scs8hd_decap_6
XFILLER_6_3777 vgnd vpwr scs8hd_decap_12
XFILLER_4_4180 vgnd vpwr scs8hd_decap_12
XFILLER_0_4000 vgnd vpwr scs8hd_decap_12
XFILLER_5_1318 vgnd vpwr scs8hd_decap_12
XFILLER_3_1086 vgnd vpwr scs8hd_decap_12
XFILLER_0_4055 vgnd vpwr scs8hd_decap_6
XPHY_439 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_428 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_417 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_406 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_1985 vgnd vpwr scs8hd_decap_12
XFILLER_7_2807 vgnd vpwr scs8hd_decap_12
XANTENNA__11__A enable vgnd vpwr scs8hd_diode_2
XFILLER_4_849 vgnd vpwr scs8hd_decap_12
XFILLER_5_3221 vgnd vpwr scs8hd_decap_12
XFILLER_5_2575 vgnd vpwr scs8hd_decap_12
XFILLER_1_2439 vgnd vpwr scs8hd_fill_1
XFILLER_6_1605 vgnd vpwr scs8hd_decap_12
XFILLER_3_3917 vgnd vpwr scs8hd_decap_12
XFILLER_1_3685 vgnd vpwr scs8hd_decap_12
X_15_ address[1] _11_/Y _13_/C address[2] _15_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_9_1284 vgnd vpwr scs8hd_decap_12
XFILLER_6_4253 vgnd vpwr scs8hd_decap_12
XFILLER_6_2862 vgnd vpwr scs8hd_decap_12
XFILLER_2_4106 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ top_width_0_height_0__pin_4_ vgnd vpwr scs8hd_diode_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_2450 vgnd vpwr scs8hd_decap_12
XFILLER_0_2472 vpwr vgnd scs8hd_fill_2
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__06__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4039 vgnd vpwr scs8hd_decap_12
XFILLER_7_2648 vgnd vpwr scs8hd_decap_12
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XFILLER_5_3051 vgnd vpwr scs8hd_decap_12
XFILLER_5_2361 vgnd vpwr scs8hd_decap_12
XFILLER_5_1660 vgnd vpwr scs8hd_decap_12
XFILLER_1_1513 vgnd vpwr scs8hd_decap_12
XFILLER_1_2258 vgnd vpwr scs8hd_decap_12
XFILLER_2_3972 vgnd vpwr scs8hd_decap_12
XPHY_781 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_770 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_792 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4551 vgnd vpwr scs8hd_decap_12
XFILLER_7_440 vgnd vpwr scs8hd_decap_12
XFILLER_6_1435 vgnd vpwr scs8hd_decap_12
XFILLER_3_3758 vgnd vpwr scs8hd_decap_12
XFILLER_1_4161 vgnd vpwr scs8hd_decap_12
XFILLER_0_1067 vgnd vpwr scs8hd_decap_12
XFILLER_1_2770 vgnd vpwr scs8hd_decap_12
XFILLER_8_4326 vgnd vpwr scs8hd_decap_12
XFILLER_8_2935 vgnd vpwr scs8hd_decap_12
XFILLER_6_4094 vgnd vpwr scs8hd_decap_12
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XFILLER_2_2545 vgnd vpwr scs8hd_decap_12
XFILLER_9_738 vgnd vpwr scs8hd_decap_6
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_410 vgnd vpwr scs8hd_decap_12
XFILLER_7_3124 vgnd vpwr scs8hd_decap_12
XFILLER_7_2445 vgnd vpwr scs8hd_decap_12
XFILLER_7_1733 vgnd vpwr scs8hd_decap_12
XFILLER_5_977 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XFILLER_1_1343 vgnd vpwr scs8hd_decap_12
XFILLER_1_2099 vgnd vpwr scs8hd_decap_12
XFILLER_8_1508 vgnd vpwr scs8hd_decap_12
XFILLER_7_281 vgnd vpwr scs8hd_decap_12
XFILLER_7_2990 vgnd vpwr scs8hd_decap_12
XFILLER_6_1276 vgnd vpwr scs8hd_decap_12
XFILLER_3_4234 vgnd vpwr scs8hd_decap_12
XFILLER_3_2843 vgnd vpwr scs8hd_decap_12
XFILLER_8_4167 vgnd vpwr scs8hd_decap_12
XFILLER_8_3411 vgnd vpwr scs8hd_decap_12
XFILLER_4_4009 vgnd vpwr scs8hd_decap_12
XFILLER_4_2618 vgnd vpwr scs8hd_decap_12
XFILLER_2_947 vgnd vpwr scs8hd_decap_12
XFILLER_2_3021 vgnd vpwr scs8hd_decap_12
XFILLER_2_1630 vgnd vpwr scs8hd_decap_12
XFILLER_2_2375 vgnd vpwr scs8hd_fill_1
XFILLER_4_4521 vgnd vpwr scs8hd_decap_12
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
XFILLER_7_1574 vgnd vpwr scs8hd_decap_12
XFILLER_4_3875 vgnd vpwr scs8hd_decap_12
XFILLER_3_1416 vgnd vpwr scs8hd_decap_12
XFILLER_0_490 vgnd vpwr scs8hd_decap_6
XFILLER_1_1184 vgnd vpwr scs8hd_decap_12
XFILLER_9_4465 vgnd vpwr scs8hd_decap_12
XFILLER_9_3764 vgnd vpwr scs8hd_decap_12
XFILLER_8_1349 vgnd vpwr scs8hd_decap_12
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XFILLER_5_4307 vgnd vpwr scs8hd_decap_12
XFILLER_5_2916 vgnd vpwr scs8hd_decap_12
XFILLER_3_4075 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XPHY_67 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_56 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_45 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_34 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__14__A _10_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_3252 vgnd vpwr scs8hd_decap_12
XFILLER_4_2437 vgnd vpwr scs8hd_decap_12
XFILLER_4_1703 vgnd vpwr scs8hd_decap_12
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_2_788 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ top_width_0_height_0__pin_0_ vgnd vpwr scs8hd_diode_2
XFILLER_2_1471 vgnd vpwr scs8hd_decap_12
XFILLER_9_354 vgnd vpwr scs8hd_decap_12
XFILLER_9_2326 vgnd vpwr scs8hd_decap_12
XFILLER_9_1625 vgnd vpwr scs8hd_decap_12
XFILLER_6_3948 vgnd vpwr scs8hd_decap_12
XFILLER_7_2050 vgnd vpwr scs8hd_decap_12
XFILLER_4_2960 vgnd vpwr scs8hd_decap_12
XFILLER_3_1257 vgnd vpwr scs8hd_decap_12
XFILLER_0_2846 vgnd vpwr scs8hd_decap_6
XFILLER_0_3547 vgnd vpwr scs8hd_decap_12
XFILLER_0_4248 vgnd vpwr scs8hd_decap_12
XFILLER_5_2746 vgnd vpwr scs8hd_decap_12
XFILLER_3_3160 vgnd vpwr scs8hd_decap_12
XANTENNA__09__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_6_324 vgnd vpwr scs8hd_decap_12
XFILLER_8_3082 vgnd vpwr scs8hd_decap_12
XFILLER_1_4502 vgnd vpwr scs8hd_decap_12
XFILLER_8_1691 vgnd vpwr scs8hd_decap_12
XFILLER_4_2289 vgnd vpwr scs8hd_decap_6
XFILLER_4_1544 vgnd vpwr scs8hd_decap_12
XFILLER_0_1408 vgnd vpwr scs8hd_decap_12
XFILLER_0_2109 vgnd vpwr scs8hd_decap_12
XFILLER_1_3856 vgnd vpwr scs8hd_decap_12
XFILLER_6_4424 vgnd vpwr scs8hd_decap_12
XFILLER_6_3789 vgnd vpwr scs8hd_decap_12
XFILLER_4_4192 vgnd vpwr scs8hd_decap_12
XFILLER_0_3311 vgnd vpwr scs8hd_decap_6
XFILLER_0_4012 vgnd vpwr scs8hd_decap_12
XPHY_407 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_2698 vgnd vpwr scs8hd_decap_12
XFILLER_0_3344 vpwr vgnd scs8hd_fill_2
XFILLER_0_3377 vpwr vgnd scs8hd_fill_2
XPHY_429 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_418 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_1997 vgnd vpwr scs8hd_decap_12
XFILLER_9_3380 vgnd vpwr scs8hd_decap_12
XFILLER_7_2819 vgnd vpwr scs8hd_decap_12
XFILLER_5_2587 vgnd vpwr scs8hd_decap_12
XFILLER_5_1831 vgnd vpwr scs8hd_decap_12
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_611 vgnd vpwr scs8hd_decap_12
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XFILLER_6_3008 vgnd vpwr scs8hd_decap_12
XFILLER_5_4490 vgnd vpwr scs8hd_decap_12
XFILLER_4_2020 vgnd vpwr scs8hd_decap_12
XFILLER_3_3929 vgnd vpwr scs8hd_decap_12
XFILLER_1_4332 vgnd vpwr scs8hd_decap_12
XFILLER_4_1374 vgnd vpwr scs8hd_decap_12
X_14_ _10_/A _11_/Y _13_/C address[2] _14_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_1_2941 vgnd vpwr scs8hd_decap_12
XFILLER_1_3697 vgnd vpwr scs8hd_decap_12
XFILLER_6_4265 vgnd vpwr scs8hd_decap_12
XFILLER_9_1296 vgnd vpwr scs8hd_decap_6
XFILLER_9_1241 vgnd vpwr scs8hd_decap_12
XFILLER_6_2874 vgnd vpwr scs8hd_decap_12
XFILLER_0_3163 vgnd vpwr scs8hd_decap_12
XFILLER_2_2716 vgnd vpwr scs8hd_decap_12
XFILLER_0_1761 vgnd vpwr scs8hd_decap_6
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_2462 vgnd vpwr scs8hd_decap_6
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__22__A gfpga_pad_GPIO_PAD[3] vgnd vpwr scs8hd_diode_2
XFILLER_7_1904 vgnd vpwr scs8hd_decap_12
XFILLER_5_3063 vgnd vpwr scs8hd_decap_12
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XFILLER_0_831 vgnd vpwr scs8hd_decap_6
XFILLER_5_2373 vgnd vpwr scs8hd_decap_6
XFILLER_5_2340 vpwr vgnd scs8hd_fill_2
XFILLER_5_1672 vgnd vpwr scs8hd_decap_12
XFILLER_2_3984 vgnd vpwr scs8hd_decap_12
XPHY_793 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_782 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_771 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_760 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4563 vgnd vpwr scs8hd_decap_12
XFILLER_7_452 vgnd vpwr scs8hd_decap_12
XFILLER_3_4405 vgnd vpwr scs8hd_decap_12
XFILLER_6_1447 vgnd vpwr scs8hd_decap_12
XFILLER_1_4173 vgnd vpwr scs8hd_decap_12
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XFILLER_0_1079 vgnd vpwr scs8hd_decap_6
XFILLER_0_1024 vgnd vpwr scs8hd_decap_12
XFILLER_1_2782 vgnd vpwr scs8hd_decap_12
XFILLER_8_4338 vgnd vpwr scs8hd_decap_12
XFILLER_8_2947 vgnd vpwr scs8hd_decap_12
XFILLER_6_3350 vgnd vpwr scs8hd_decap_12
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XANTENNA__17__A gfpga_pad_GPIO_PAD[6] vgnd vpwr scs8hd_diode_2
XFILLER_2_1801 vgnd vpwr scs8hd_decap_12
XFILLER_2_2557 vgnd vpwr scs8hd_decap_12
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_989 vgnd vpwr scs8hd_decap_8
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XFILLER_4_422 vgnd vpwr scs8hd_decap_12
XFILLER_7_3136 vgnd vpwr scs8hd_decap_12
XFILLER_7_2457 vgnd vpwr scs8hd_decap_12
XFILLER_7_1745 vgnd vpwr scs8hd_decap_12
XFILLER_2_4460 vgnd vpwr scs8hd_decap_12
XFILLER_0_683 vgnd vpwr scs8hd_decap_12
XFILLER_1_2001 vgnd vpwr scs8hd_decap_12
XFILLER_1_1355 vgnd vpwr scs8hd_decap_12
XPHY_590 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4393 vgnd vpwr scs8hd_decap_12
XFILLER_7_293 vgnd vpwr scs8hd_decap_12
XFILLER_3_4246 vgnd vpwr scs8hd_decap_12
XFILLER_6_1288 vgnd vpwr scs8hd_decap_12
XFILLER_3_2855 vgnd vpwr scs8hd_decap_12
XFILLER_8_3423 vgnd vpwr scs8hd_decap_12
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XFILLER_8_2777 vgnd vpwr scs8hd_decap_12
XFILLER_6_3191 vgnd vpwr scs8hd_decap_12
XFILLER_1_403 vgnd vpwr scs8hd_decap_12
XFILLER_2_959 vgnd vpwr scs8hd_decap_12
XFILLER_2_3033 vgnd vpwr scs8hd_decap_12
XFILLER_2_1642 vgnd vpwr scs8hd_decap_12
XFILLER_2_2387 vgnd vpwr scs8hd_decap_12
XFILLER_7_2221 vgnd vpwr scs8hd_decap_12
XFILLER_5_720 vgnd vpwr scs8hd_decap_12
XFILLER_4_4533 vgnd vpwr scs8hd_decap_12
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XFILLER_4_3887 vgnd vpwr scs8hd_decap_12
XFILLER_3_1428 vgnd vpwr scs8hd_decap_12
XFILLER_1_1196 vgnd vpwr scs8hd_decap_12
XFILLER_9_4477 vgnd vpwr scs8hd_decap_12
XFILLER_9_3721 vgnd vpwr scs8hd_decap_12
XFILLER_9_3776 vgnd vpwr scs8hd_decap_6
XFILLER_5_4319 vgnd vpwr scs8hd_decap_12
XFILLER_3_3331 vgnd vpwr scs8hd_decap_12
XPHY_13 vgnd vpwr scs8hd_decap_3
XFILLER_3_2685 vgnd vpwr scs8hd_decap_12
XFILLER_3_1940 vgnd vpwr scs8hd_decap_12
XPHY_46 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_35 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_24 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_68 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_57 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__14__B _11_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_4_3106 vgnd vpwr scs8hd_decap_12
XFILLER_8_1862 vgnd vpwr scs8hd_decap_12
XFILLER_4_2449 vgnd vpwr scs8hd_decap_12
XFILLER_4_1715 vgnd vpwr scs8hd_decap_12
XFILLER_2_1483 vgnd vpwr scs8hd_decap_12
XFILLER_9_366 vgnd vpwr scs8hd_decap_6
XFILLER_9_311 vgnd vpwr scs8hd_decap_12
XFILLER_5_550 vgnd vpwr scs8hd_decap_12
XFILLER_9_3039 vgnd vpwr scs8hd_decap_12
XFILLER_9_2338 vgnd vpwr scs8hd_decap_12
XFILLER_9_1637 vgnd vpwr scs8hd_decap_6
XFILLER_7_2062 vgnd vpwr scs8hd_decap_12
XFILLER_4_4363 vgnd vpwr scs8hd_decap_12
XFILLER_4_2972 vgnd vpwr scs8hd_decap_12
XFILLER_3_1269 vgnd vpwr scs8hd_decap_12
XFILLER_0_2803 vgnd vpwr scs8hd_decap_12
XFILLER_0_3504 vgnd vpwr scs8hd_decap_12
XFILLER_0_3559 vgnd vpwr scs8hd_decap_6
XFILLER_9_4241 vgnd vpwr scs8hd_decap_6
XFILLER_5_4149 vgnd vpwr scs8hd_decap_12
XFILLER_5_3404 vgnd vpwr scs8hd_decap_12
XFILLER_5_2758 vgnd vpwr scs8hd_decap_12
XANTENNA__09__B enable vgnd vpwr scs8hd_diode_2
XFILLER_3_1770 vgnd vpwr scs8hd_decap_12
XFILLER_8_3094 vgnd vpwr scs8hd_decap_12
XFILLER_2_520 vgnd vpwr scs8hd_decap_12
XFILLER_1_3868 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_2102 vgnd vpwr scs8hd_decap_6
XFILLER_6_4436 vgnd vpwr scs8hd_decap_12
XFILLER_5_391 vgnd vpwr scs8hd_decap_12
XFILLER_9_1489 vgnd vpwr scs8hd_decap_12
XFILLER_0_4024 vgnd vpwr scs8hd_decap_6
XPHY_419 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_408 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1099 vgnd vpwr scs8hd_decap_12
XFILLER_0_1954 vgnd vpwr scs8hd_decap_12
XFILLER_9_4093 vgnd vpwr scs8hd_decap_12
XFILLER_9_3392 vgnd vpwr scs8hd_decap_12
XFILLER_5_3234 vgnd vpwr scs8hd_decap_12
XFILLER_3_306 vgnd vpwr scs8hd_decap_12
XFILLER_9_2691 vgnd vpwr scs8hd_decap_6
XFILLER_5_2599 vgnd vpwr scs8hd_decap_12
XFILLER_5_1843 vgnd vpwr scs8hd_decap_12
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XFILLER_7_623 vgnd vpwr scs8hd_decap_12
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_6_1618 vgnd vpwr scs8hd_decap_12
XFILLER_4_2032 vgnd vpwr scs8hd_decap_12
XFILLER_1_4344 vgnd vpwr scs8hd_decap_12
XFILLER_2_361 vgnd vpwr scs8hd_decap_12
XFILLER_4_1386 vgnd vpwr scs8hd_decap_12
X_13_ address[1] _11_/Y _13_/C _10_/D _13_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_1_2953 vgnd vpwr scs8hd_decap_12
XFILLER_8_4509 vgnd vpwr scs8hd_decap_12
XFILLER_6_4277 vgnd vpwr scs8hd_decap_12
XFILLER_6_3521 vgnd vpwr scs8hd_decap_12
XFILLER_2_4119 vgnd vpwr scs8hd_decap_12
XFILLER_9_1253 vgnd vpwr scs8hd_decap_12
XFILLER_6_2886 vgnd vpwr scs8hd_decap_12
XFILLER_0_3175 vgnd vpwr scs8hd_decap_12
XFILLER_2_2728 vgnd vpwr scs8hd_decap_12
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3307 vgnd vpwr scs8hd_decap_12
XFILLER_7_1916 vgnd vpwr scs8hd_decap_12
XFILLER_5_3075 vgnd vpwr scs8hd_decap_12
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
XFILLER_5_2396 vgnd vpwr scs8hd_decap_12
XFILLER_5_1684 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _09_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_1526 vgnd vpwr scs8hd_decap_12
XPHY_794 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_783 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_772 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_761 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_750 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_910 vgnd vpwr scs8hd_decap_12
XFILLER_7_464 vgnd vpwr scs8hd_decap_12
XFILLER_3_4417 vgnd vpwr scs8hd_decap_12
XFILLER_6_1459 vgnd vpwr scs8hd_decap_12
XFILLER_1_4185 vgnd vpwr scs8hd_decap_12
XFILLER_0_1036 vgnd vpwr scs8hd_decap_12
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_1_2794 vgnd vpwr scs8hd_decap_12
XFILLER_6_3362 vgnd vpwr scs8hd_decap_12
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XFILLER_2_3204 vgnd vpwr scs8hd_decap_12
XFILLER_6_1971 vgnd vpwr scs8hd_decap_12
XFILLER_2_1813 vgnd vpwr scs8hd_decap_12
XFILLER_2_2569 vgnd vpwr scs8hd_decap_12
XFILLER_9_707 vgnd vpwr scs8hd_decap_6
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XFILLER_7_3148 vgnd vpwr scs8hd_decap_12
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XFILLER_4_434 vgnd vpwr scs8hd_decap_12
XFILLER_7_2469 vgnd vpwr scs8hd_decap_12
XFILLER_7_2436 vgnd vpwr scs8hd_fill_1
XFILLER_7_1757 vgnd vpwr scs8hd_decap_12
XFILLER_5_2160 vgnd vpwr scs8hd_decap_12
XFILLER_2_4472 vgnd vpwr scs8hd_decap_12
XFILLER_0_695 vgnd vpwr scs8hd_decap_12
XFILLER_1_1367 vgnd vpwr scs8hd_decap_12
XFILLER_8_751 vgnd vpwr scs8hd_decap_12
XPHY_591 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_580 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3969 vgnd vpwr scs8hd_decap_12
XFILLER_3_4258 vgnd vpwr scs8hd_decap_12
XFILLER_3_3502 vgnd vpwr scs8hd_decap_12
XFILLER_1_3270 vgnd vpwr scs8hd_decap_12
XFILLER_8_3435 vgnd vpwr scs8hd_decap_12
XFILLER_1_415 vgnd vpwr scs8hd_decap_12
XFILLER_8_2789 vgnd vpwr scs8hd_decap_12
XFILLER_2_2344 vpwr vgnd scs8hd_fill_2
XFILLER_2_3045 vgnd vpwr scs8hd_decap_12
XFILLER_0_2090 vgnd vpwr scs8hd_decap_12
XFILLER_2_1654 vgnd vpwr scs8hd_decap_12
XFILLER_2_2399 vgnd vpwr scs8hd_decap_8
XFILLER_9_559 vgnd vpwr scs8hd_decap_12
XFILLER_9_2509 vpwr vgnd scs8hd_fill_2
XFILLER_7_2233 vgnd vpwr scs8hd_decap_12
XFILLER_4_4578 vgnd vpwr scs8hd_decap_3
XFILLER_7_1587 vgnd vpwr scs8hd_decap_12
XFILLER_4_3899 vgnd vpwr scs8hd_decap_12
XFILLER_9_4489 vgnd vpwr scs8hd_decap_6
XFILLER_9_4434 vgnd vpwr scs8hd_decap_12
XFILLER_9_3733 vgnd vpwr scs8hd_decap_12
XFILLER_8_2008 vgnd vpwr scs8hd_decap_12
XFILLER_8_581 vgnd vpwr scs8hd_decap_12
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_3490 vgnd vpwr scs8hd_decap_12
XFILLER_6_1020 vgnd vpwr scs8hd_decap_12
XFILLER_5_2929 vgnd vpwr scs8hd_decap_12
XFILLER_3_4088 vgnd vpwr scs8hd_decap_12
XFILLER_3_3343 vgnd vpwr scs8hd_decap_12
XPHY_14 vgnd vpwr scs8hd_decap_3
XFILLER_3_2697 vgnd vpwr scs8hd_decap_12
XPHY_69 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_58 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_47 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_36 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_25 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_507 vgnd vpwr scs8hd_decap_12
XANTENNA__14__C _13_/C vgnd vpwr scs8hd_diode_2
XFILLER_8_3265 vgnd vpwr scs8hd_decap_12
XFILLER_8_2520 vgnd vpwr scs8hd_decap_12
XFILLER_4_3118 vgnd vpwr scs8hd_decap_12
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_8_1874 vgnd vpwr scs8hd_decap_12
XFILLER_8_1841 vgnd vpwr scs8hd_fill_1
XFILLER_4_1727 vgnd vpwr scs8hd_decap_12
XFILLER_2_2130 vgnd vpwr scs8hd_decap_12
XFILLER_9_323 vgnd vpwr scs8hd_decap_12
XFILLER_5_562 vgnd vpwr scs8hd_decap_12
XFILLER_4_4375 vgnd vpwr scs8hd_decap_12
XFILLER_0_3516 vgnd vpwr scs8hd_decap_12
XFILLER_0_4217 vgnd vpwr scs8hd_decap_12
XFILLER_4_2984 vgnd vpwr scs8hd_decap_12
XFILLER_0_2815 vgnd vpwr scs8hd_decap_6
XFILLER_9_2884 vgnd vpwr scs8hd_decap_12
XFILLER_3_3173 vgnd vpwr scs8hd_decap_12
XANTENNA__09__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_3_1782 vgnd vpwr scs8hd_decap_12
XFILLER_6_337 vgnd vpwr scs8hd_decap_12
XFILLER_8_2350 vgnd vpwr scs8hd_decap_12
XFILLER_4_2203 vgnd vpwr scs8hd_decap_12
XFILLER_1_4515 vgnd vpwr scs8hd_decap_12
XFILLER_2_532 vgnd vpwr scs8hd_decap_12
XFILLER_4_1557 vgnd vpwr scs8hd_decap_12
XFILLER_6_4448 vgnd vpwr scs8hd_decap_12
XFILLER_4_3460 vgnd vpwr scs8hd_decap_12
XFILLER_3_1001 vgnd vpwr scs8hd_decap_12
XFILLER_0_3357 vgnd vpwr scs8hd_decap_12
XPHY_409 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_1966 vgnd vpwr scs8hd_decap_12
XFILLER_0_2667 vgnd vpwr scs8hd_decap_12
XFILLER_3_318 vgnd vpwr scs8hd_decap_12
XFILLER_5_3246 vgnd vpwr scs8hd_decap_12
XFILLER_5_1855 vgnd vpwr scs8hd_decap_12
XFILLER_0_4570 vgnd vpwr scs8hd_decap_8
XPHY_910 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_635 vgnd vpwr scs8hd_decap_12
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
XFILLER_3_830 vgnd vpwr scs8hd_decap_12
XFILLER_8_2191 vgnd vpwr scs8hd_decap_12
X_12_ _10_/A _11_/Y _13_/C _10_/D _12_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_1_3600 vgnd vpwr scs8hd_decap_12
XFILLER_1_4356 vgnd vpwr scs8hd_decap_12
XFILLER_2_373 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ top_width_0_height_0__pin_4_ logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[2] vgnd vpwr scs8hd_ebufn_1
XFILLER_4_1398 vgnd vpwr scs8hd_decap_12
XFILLER_1_2965 vgnd vpwr scs8hd_decap_12
XFILLER_9_1265 vgnd vpwr scs8hd_decap_6
XFILLER_9_1210 vgnd vpwr scs8hd_decap_12
XFILLER_6_4289 vgnd vpwr scs8hd_decap_12
XFILLER_6_3533 vgnd vpwr scs8hd_decap_12
XFILLER_6_690 vgnd vpwr scs8hd_decap_12
XFILLER_0_1730 vgnd vpwr scs8hd_decap_6
XFILLER_0_2431 vgnd vpwr scs8hd_decap_12
XFILLER_0_3132 vgnd vpwr scs8hd_decap_12
XFILLER_0_3187 vgnd vpwr scs8hd_decap_6
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3319 vgnd vpwr scs8hd_decap_12
XFILLER_4_605 vgnd vpwr scs8hd_decap_12
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
XFILLER_7_1928 vgnd vpwr scs8hd_decap_12
XFILLER_5_3087 vgnd vpwr scs8hd_decap_12
XFILLER_5_2353 vpwr vgnd scs8hd_fill_2
XFILLER_0_800 vgnd vpwr scs8hd_decap_6
XFILLER_5_1696 vgnd vpwr scs8hd_decap_12
XFILLER_1_1538 vgnd vpwr scs8hd_decap_12
XFILLER_2_3997 vgnd vpwr scs8hd_decap_12
XPHY_795 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_784 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_773 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_762 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_751 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_740 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_955 vgnd vpwr scs8hd_decap_12
XFILLER_8_922 vgnd vpwr scs8hd_decap_12
XFILLER_7_476 vgnd vpwr scs8hd_decap_12
XFILLER_7_4576 vgnd vpwr scs8hd_decap_4
XFILLER_7_3831 vgnd vpwr scs8hd_decap_12
XFILLER_6_2106 vgnd vpwr scs8hd_decap_12
XFILLER_3_4429 vgnd vpwr scs8hd_decap_12
XFILLER_1_3441 vgnd vpwr scs8hd_decap_12
XFILLER_1_4197 vgnd vpwr scs8hd_decap_12
XFILLER_0_1048 vgnd vpwr scs8hd_decap_6
XFILLER_8_3606 vgnd vpwr scs8hd_decap_12
XFILLER_6_3374 vgnd vpwr scs8hd_decap_12
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XFILLER_2_3216 vgnd vpwr scs8hd_decap_12
XFILLER_0_1582 vgnd vpwr scs8hd_decap_12
XFILLER_2_1825 vgnd vpwr scs8hd_decap_12
XFILLER_5_903 vgnd vpwr scs8hd_decap_12
XFILLER_7_2404 vgnd vpwr scs8hd_decap_12
XFILLER_4_446 vgnd vpwr scs8hd_decap_12
XFILLER_5_2172 vgnd vpwr scs8hd_decap_12
XFILLER_0_652 vgnd vpwr scs8hd_decap_12
XFILLER_1_2014 vgnd vpwr scs8hd_decap_12
XPHY_570 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_1379 vgnd vpwr scs8hd_decap_12
XPHY_592 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_581 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_3661 vgnd vpwr scs8hd_decap_12
XFILLER_3_3514 vgnd vpwr scs8hd_decap_12
XFILLER_3_2868 vgnd vpwr scs8hd_decap_12
XFILLER_1_3282 vgnd vpwr scs8hd_decap_12
XFILLER_2_2323 vpwr vgnd scs8hd_fill_2
XFILLER_2_3057 vgnd vpwr scs8hd_decap_12
XFILLER_2_1666 vgnd vpwr scs8hd_decap_12
XFILLER_5_733 vgnd vpwr scs8hd_decap_12
XFILLER_7_2245 vgnd vpwr scs8hd_decap_12
XFILLER_4_4546 vgnd vpwr scs8hd_decap_12
XFILLER_4_3801 vgnd vpwr scs8hd_decap_12
XFILLER_4_276 vgnd vpwr scs8hd_decap_12
XFILLER_7_1599 vgnd vpwr scs8hd_decap_12
XFILLER_9_4446 vgnd vpwr scs8hd_decap_12
XFILLER_9_3745 vgnd vpwr scs8hd_decap_6
XFILLER_8_593 vgnd vpwr scs8hd_decap_12
XFILLER_6_1032 vgnd vpwr scs8hd_decap_12
XPHY_15 vgnd vpwr scs8hd_decap_3
XFILLER_3_1953 vgnd vpwr scs8hd_decap_12
XPHY_59 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_48 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_37 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_26 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__14__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_8_3277 vgnd vpwr scs8hd_decap_12
XFILLER_4_2407 vgnd vpwr scs8hd_decap_3
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_2_703 vgnd vpwr scs8hd_decap_12
XFILLER_8_1886 vgnd vpwr scs8hd_decap_12
XFILLER_2_2142 vgnd vpwr scs8hd_decap_12
XFILLER_9_335 vgnd vpwr scs8hd_decap_6
XFILLER_2_1496 vgnd vpwr scs8hd_decap_12
XFILLER_9_3008 vgnd vpwr scs8hd_decap_12
XFILLER_9_2307 vgnd vpwr scs8hd_decap_12
XFILLER_9_1606 vgnd vpwr scs8hd_decap_6
XFILLER_5_574 vgnd vpwr scs8hd_decap_12
XFILLER_7_2075 vgnd vpwr scs8hd_decap_12
XFILLER_7_1330 vgnd vpwr scs8hd_decap_12
XFILLER_4_4387 vgnd vpwr scs8hd_decap_12
XFILLER_4_3631 vgnd vpwr scs8hd_decap_12
XFILLER_0_3528 vgnd vpwr scs8hd_decap_6
XFILLER_0_4229 vgnd vpwr scs8hd_decap_12
XFILLER_4_2996 vgnd vpwr scs8hd_decap_12
XFILLER_9_4210 vgnd vpwr scs8hd_decap_6
XFILLER_9_3597 vgnd vpwr scs8hd_decap_12
XFILLER_9_2896 vgnd vpwr scs8hd_decap_12
XFILLER_8_1105 vgnd vpwr scs8hd_decap_12
XFILLER_5_3417 vgnd vpwr scs8hd_decap_12
XFILLER_3_3185 vgnd vpwr scs8hd_decap_12
XANTENNA__09__D _10_/D vgnd vpwr scs8hd_diode_2
XFILLER_7_806 vgnd vpwr scs8hd_decap_12
XFILLER_3_1794 vgnd vpwr scs8hd_decap_12
XFILLER_6_349 vgnd vpwr scs8hd_decap_12
XFILLER_8_2362 vgnd vpwr scs8hd_decap_12
XFILLER_4_2215 vgnd vpwr scs8hd_decap_12
XFILLER_1_4527 vgnd vpwr scs8hd_decap_12
XFILLER_2_544 vgnd vpwr scs8hd_decap_12
XFILLER_4_1569 vgnd vpwr scs8hd_decap_12
XFILLER_9_187 vgnd vpwr scs8hd_decap_12
XFILLER_6_3704 vgnd vpwr scs8hd_decap_12
XFILLER_6_861 vgnd vpwr scs8hd_decap_12
XFILLER_9_1458 vgnd vpwr scs8hd_decap_12
XFILLER_7_1160 vgnd vpwr scs8hd_decap_12
XFILLER_4_3472 vgnd vpwr scs8hd_decap_12
XFILLER_3_1013 vgnd vpwr scs8hd_decap_12
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XFILLER_0_1923 vgnd vpwr scs8hd_decap_12
XFILLER_0_3369 vgnd vpwr scs8hd_decap_8
XFILLER_0_1978 vgnd vpwr scs8hd_decap_6
XFILLER_0_2679 vgnd vpwr scs8hd_decap_12
XFILLER_9_4062 vgnd vpwr scs8hd_decap_12
XFILLER_9_3361 vgnd vpwr scs8hd_decap_12
XFILLER_9_2660 vgnd vpwr scs8hd_decap_6
XFILLER_5_3258 vgnd vpwr scs8hd_decap_12
XFILLER_5_2502 vgnd vpwr scs8hd_decap_12
XPHY_911 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_900 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_1867 vgnd vpwr scs8hd_decap_12
XFILLER_3_2270 vgnd vpwr scs8hd_decap_12
XFILLER_1_1709 vgnd vpwr scs8hd_decap_12
XFILLER_7_647 vgnd vpwr scs8hd_decap_12
XFILLER_3_842 vgnd vpwr scs8hd_decap_12
X_11_ enable _11_/Y vgnd vpwr scs8hd_inv_8
XFILLER_5_3770 vgnd vpwr scs8hd_decap_12
XFILLER_4_2045 vgnd vpwr scs8hd_decap_12
XFILLER_4_1300 vgnd vpwr scs8hd_decap_12
XFILLER_1_3612 vgnd vpwr scs8hd_decap_12
XFILLER_1_4368 vgnd vpwr scs8hd_decap_12
XFILLER_2_385 vgnd vpwr scs8hd_decap_12
XFILLER_1_2977 vgnd vpwr scs8hd_decap_12
XFILLER_9_1222 vgnd vpwr scs8hd_decap_12
XFILLER_6_3545 vgnd vpwr scs8hd_decap_12
XFILLER_6_2899 vgnd vpwr scs8hd_decap_12
XFILLER_0_2443 vgnd vpwr scs8hd_decap_6
XFILLER_0_2476 vgnd vpwr scs8hd_decap_4
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_3144 vgnd vpwr scs8hd_decap_12
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_617 vgnd vpwr scs8hd_decap_12
XFILLER_5_3099 vgnd vpwr scs8hd_decap_12
XPHY_763 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_752 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_741 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_730 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_796 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_785 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_774 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_967 vgnd vpwr scs8hd_decap_12
XFILLER_8_934 vgnd vpwr scs8hd_decap_12
XFILLER_6_2118 vgnd vpwr scs8hd_decap_12
XFILLER_3_672 vgnd vpwr scs8hd_decap_12
XFILLER_4_1130 vgnd vpwr scs8hd_decap_12
XFILLER_0_1005 vgnd vpwr scs8hd_decap_12
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_1_3453 vgnd vpwr scs8hd_decap_12
XFILLER_9_94 vgnd vpwr scs8hd_decap_12
XFILLER_8_3618 vgnd vpwr scs8hd_decap_12
XFILLER_6_4021 vgnd vpwr scs8hd_decap_12
XFILLER_6_2630 vgnd vpwr scs8hd_decap_12
XFILLER_6_1984 vgnd vpwr scs8hd_decap_12
XFILLER_2_3228 vgnd vpwr scs8hd_decap_12
XFILLER_0_1594 vgnd vpwr scs8hd_decap_12
XFILLER_2_1837 vgnd vpwr scs8hd_decap_12
XFILLER_7_2416 vgnd vpwr scs8hd_decap_12
XFILLER_0_664 vgnd vpwr scs8hd_decap_12
XFILLER_5_2184 vgnd vpwr scs8hd_decap_12
XFILLER_2_4485 vgnd vpwr scs8hd_decap_12
XFILLER_1_2026 vgnd vpwr scs8hd_decap_12
XFILLER_2_3740 vgnd vpwr scs8hd_decap_12
XPHY_593 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_582 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_571 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_560 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3938 vgnd vpwr scs8hd_decap_12
XFILLER_8_764 vgnd vpwr scs8hd_decap_12
XFILLER_7_3673 vgnd vpwr scs8hd_decap_12
XFILLER_6_1203 vgnd vpwr scs8hd_decap_12
XFILLER_3_3526 vgnd vpwr scs8hd_decap_12
XFILLER_1_1892 vgnd vpwr scs8hd_decap_12
XFILLER_8_3448 vgnd vpwr scs8hd_decap_12
XFILLER_8_2703 vgnd vpwr scs8hd_decap_12
XFILLER_1_428 vgnd vpwr scs8hd_decap_12
XFILLER_2_3069 vgnd vpwr scs8hd_decap_12
XFILLER_9_528 vgnd vpwr scs8hd_decap_12
XFILLER_5_745 vgnd vpwr scs8hd_decap_12
XFILLER_8_3960 vgnd vpwr scs8hd_decap_12
XFILLER_7_1501 vgnd vpwr scs8hd_decap_12
XFILLER_4_4558 vgnd vpwr scs8hd_decap_12
XFILLER_4_288 vgnd vpwr scs8hd_decap_12
XFILLER_1_940 vgnd vpwr scs8hd_decap_12
XFILLER_1_1111 vgnd vpwr scs8hd_decap_12
XFILLER_2_3570 vgnd vpwr scs8hd_decap_12
XFILLER_9_4403 vgnd vpwr scs8hd_decap_12
XPHY_390 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_4458 vgnd vpwr scs8hd_decap_6
XFILLER_9_3702 vgnd vpwr scs8hd_decap_12
XFILLER_3_4002 vgnd vpwr scs8hd_decap_12
XFILLER_6_1044 vgnd vpwr scs8hd_decap_12
XFILLER_3_3356 vgnd vpwr scs8hd_decap_12
XFILLER_3_2611 vgnd vpwr scs8hd_decap_12
XFILLER_3_1965 vgnd vpwr scs8hd_decap_12
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_38 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_27 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_715 vgnd vpwr scs8hd_decap_12
XFILLER_8_3289 vgnd vpwr scs8hd_decap_12
XFILLER_8_2533 vgnd vpwr scs8hd_decap_12
XFILLER_3_4580 vgnd vpwr scs8hd_fill_1
XFILLER_1_269 vgnd vpwr scs8hd_decap_12
XFILLER_8_1898 vgnd vpwr scs8hd_decap_12
XFILLER_2_2154 vgnd vpwr scs8hd_decap_12
XFILLER_9_2319 vgnd vpwr scs8hd_decap_6
XFILLER_5_586 vgnd vpwr scs8hd_decap_12
XFILLER_7_2087 vgnd vpwr scs8hd_decap_12
XFILLER_4_4399 vgnd vpwr scs8hd_decap_12
XFILLER_4_3643 vgnd vpwr scs8hd_decap_12
XFILLER_1_781 vgnd vpwr scs8hd_decap_12
XFILLER_0_280 vgnd vpwr scs8hd_decap_12
XFILLER_9_881 vgnd vpwr scs8hd_decap_12
XFILLER_9_2853 vgnd vpwr scs8hd_decap_12
XFILLER_8_1117 vgnd vpwr scs8hd_decap_12
XFILLER_5_3429 vgnd vpwr scs8hd_decap_12
XFILLER_3_3197 vgnd vpwr scs8hd_decap_12
XFILLER_3_2441 vgnd vpwr scs8hd_decap_12
XFILLER_7_818 vgnd vpwr scs8hd_decap_12
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_556 vgnd vpwr scs8hd_decap_12
XFILLER_8_2374 vgnd vpwr scs8hd_decap_12
XFILLER_5_3941 vgnd vpwr scs8hd_decap_12
XFILLER_1_4539 vgnd vpwr scs8hd_decap_12
XFILLER_9_199 vgnd vpwr scs8hd_decap_12
XFILLER_6_873 vgnd vpwr scs8hd_decap_12
XFILLER_6_3716 vgnd vpwr scs8hd_decap_12
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XFILLER_7_1172 vgnd vpwr scs8hd_decap_12
XFILLER_4_3484 vgnd vpwr scs8hd_decap_12
XFILLER_3_1025 vgnd vpwr scs8hd_decap_12
XFILLER_0_1935 vgnd vpwr scs8hd_decap_12
XFILLER_0_2636 vgnd vpwr scs8hd_decap_12
XFILLER_9_4074 vgnd vpwr scs8hd_decap_12
XFILLER_9_3373 vgnd vpwr scs8hd_decap_6
XFILLER_5_2514 vgnd vpwr scs8hd_decap_12
XPHY_912 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_901 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_1879 vgnd vpwr scs8hd_decap_12
XFILLER_3_2282 vgnd vpwr scs8hd_decap_12
XFILLER_7_659 vgnd vpwr scs8hd_decap_12
X_10_ _10_/A enable address[3] _10_/D _10_/X vgnd vpwr scs8hd_and4_4
XFILLER_4_2057 vgnd vpwr scs8hd_decap_12
XFILLER_1_3624 vgnd vpwr scs8hd_decap_12
XFILLER_9_1234 vgnd vpwr scs8hd_decap_6
XFILLER_6_3557 vgnd vpwr scs8hd_decap_12
XFILLER_6_2801 vgnd vpwr scs8hd_decap_12
XFILLER_0_3101 vgnd vpwr scs8hd_decap_12
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_3156 vgnd vpwr scs8hd_decap_6
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_629 vgnd vpwr scs8hd_decap_12
XFILLER_0_3690 vgnd vpwr scs8hd_decap_12
XFILLER_2_3911 vgnd vpwr scs8hd_decap_12
XPHY_786 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_775 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_764 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_753 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_742 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_731 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_720 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_797 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_979 vgnd vpwr scs8hd_decap_12
XFILLER_7_489 vgnd vpwr scs8hd_decap_12
XFILLER_7_3844 vgnd vpwr scs8hd_decap_12
XFILLER_3_684 vgnd vpwr scs8hd_decap_12
XFILLER_1_4100 vgnd vpwr scs8hd_decap_12
XFILLER_4_1142 vgnd vpwr scs8hd_decap_12
XFILLER_0_1017 vgnd vpwr scs8hd_decap_6
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_1_3465 vgnd vpwr scs8hd_decap_12
XFILLER_6_4033 vgnd vpwr scs8hd_decap_12
XFILLER_9_1086 vgnd vpwr scs8hd_decap_12
XFILLER_6_3387 vgnd vpwr scs8hd_decap_12
XFILLER_6_2642 vgnd vpwr scs8hd_decap_12
XFILLER_6_1996 vgnd vpwr scs8hd_decap_12
XFILLER_2_1849 vgnd vpwr scs8hd_decap_12
XFILLER_0_1551 vgnd vpwr scs8hd_decap_12
XFILLER_5_916 vgnd vpwr scs8hd_decap_12
XFILLER_7_2439 vgnd vpwr scs8hd_fill_1
XFILLER_7_2428 vgnd vpwr scs8hd_decap_8
XFILLER_4_459 vgnd vpwr scs8hd_decap_12
XFILLER_0_676 vgnd vpwr scs8hd_decap_6
XFILLER_0_621 vgnd vpwr scs8hd_decap_12
XFILLER_5_1440 vgnd vpwr scs8hd_decap_12
XFILLER_2_4497 vgnd vpwr scs8hd_decap_12
XFILLER_1_2038 vgnd vpwr scs8hd_decap_12
XPHY_594 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_583 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_572 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_561 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_550 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_776 vgnd vpwr scs8hd_decap_12
XFILLER_4_971 vgnd vpwr scs8hd_decap_12
XFILLER_7_3685 vgnd vpwr scs8hd_decap_12
XFILLER_6_1215 vgnd vpwr scs8hd_decap_12
XFILLER_1_2550 vgnd vpwr scs8hd_decap_12
XFILLER_1_3295 vgnd vpwr scs8hd_decap_12
XFILLER_8_4106 vgnd vpwr scs8hd_decap_12
XFILLER_6_2472 vgnd vpwr scs8hd_decap_12
XFILLER_0_2071 vgnd vpwr scs8hd_decap_6
XFILLER_2_1679 vgnd vpwr scs8hd_decap_12
XFILLER_2_2303 vgnd vpwr scs8hd_decap_3
XFILLER_5_757 vgnd vpwr scs8hd_decap_12
XFILLER_8_3972 vgnd vpwr scs8hd_decap_12
XFILLER_7_2258 vgnd vpwr scs8hd_decap_12
XFILLER_7_1513 vgnd vpwr scs8hd_decap_12
XFILLER_4_3814 vgnd vpwr scs8hd_decap_12
XFILLER_1_952 vgnd vpwr scs8hd_decap_12
XFILLER_2_3582 vgnd vpwr scs8hd_decap_12
XFILLER_1_1123 vgnd vpwr scs8hd_decap_12
XFILLER_9_4415 vgnd vpwr scs8hd_decap_12
XFILLER_9_3714 vgnd vpwr scs8hd_decap_6
XPHY_391 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_380 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4161 vgnd vpwr scs8hd_decap_12
XFILLER_7_2770 vgnd vpwr scs8hd_decap_12
XFILLER_3_4014 vgnd vpwr scs8hd_decap_12
XPHY_17 vgnd vpwr scs8hd_decap_3
XFILLER_6_1056 vgnd vpwr scs8hd_decap_12
XFILLER_3_3368 vgnd vpwr scs8hd_decap_12
XFILLER_3_1977 vgnd vpwr scs8hd_decap_12
XPHY_28 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_2391 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_727 vgnd vpwr scs8hd_decap_12
XFILLER_8_2545 vgnd vpwr scs8hd_decap_12
XFILLER_3_3880 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _10_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_1410 vgnd vpwr scs8hd_decap_12
XFILLER_9_304 vgnd vpwr scs8hd_decap_6
XFILLER_5_598 vgnd vpwr scs8hd_decap_12
XFILLER_7_2099 vgnd vpwr scs8hd_decap_12
XFILLER_7_1343 vgnd vpwr scs8hd_decap_12
XFILLER_4_3655 vgnd vpwr scs8hd_decap_12
XFILLER_0_292 vgnd vpwr scs8hd_decap_12
XFILLER_9_3566 vgnd vpwr scs8hd_decap_12
XFILLER_9_893 vgnd vpwr scs8hd_decap_6
XFILLER_9_2865 vgnd vpwr scs8hd_decap_12
XFILLER_3_2453 vgnd vpwr scs8hd_decap_12
XFILLER_8_3021 vgnd vpwr scs8hd_decap_12
XFILLER_5_3953 vgnd vpwr scs8hd_decap_12
XFILLER_2_568 vgnd vpwr scs8hd_decap_12
XFILLER_8_2386 vgnd vpwr scs8hd_decap_12
XFILLER_8_1630 vgnd vpwr scs8hd_decap_12
XFILLER_4_2228 vgnd vpwr scs8hd_decap_12
XFILLER_9_156 vgnd vpwr scs8hd_decap_12
XFILLER_9_1427 vgnd vpwr scs8hd_decap_12
XFILLER_6_3728 vgnd vpwr scs8hd_decap_12
XFILLER_4_4131 vgnd vpwr scs8hd_decap_12
XFILLER_4_3496 vgnd vpwr scs8hd_decap_12
XFILLER_4_2740 vgnd vpwr scs8hd_decap_12
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
XFILLER_7_1184 vgnd vpwr scs8hd_decap_12
XFILLER_0_1947 vgnd vpwr scs8hd_decap_6
XFILLER_0_2648 vgnd vpwr scs8hd_decap_12
XFILLER_9_4086 vgnd vpwr scs8hd_decap_6
XFILLER_9_4031 vgnd vpwr scs8hd_decap_12
XFILLER_9_3330 vgnd vpwr scs8hd_decap_12
XFILLER_5_2526 vgnd vpwr scs8hd_decap_12
XFILLER_3_2294 vgnd vpwr scs8hd_fill_1
XFILLER_0_4551 vgnd vpwr scs8hd_decap_6
XPHY_913 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_902 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_3783 vgnd vpwr scs8hd_decap_12
XFILLER_3_855 vgnd vpwr scs8hd_decap_12
XFILLER_2_398 vgnd vpwr scs8hd_decap_12
XFILLER_8_1471 vgnd vpwr scs8hd_decap_12
XFILLER_4_2069 vgnd vpwr scs8hd_decap_12
XFILLER_4_1313 vgnd vpwr scs8hd_decap_12
XFILLER_1_3636 vgnd vpwr scs8hd_decap_12
XFILLER_2_1081 vgnd vpwr scs8hd_decap_12
XFILLER_6_4204 vgnd vpwr scs8hd_decap_12
XFILLER_6_2813 vgnd vpwr scs8hd_decap_12
XFILLER_4_2581 vgnd vpwr scs8hd_decap_12
XFILLER_0_2401 vgnd vpwr scs8hd_decap_12
XFILLER_0_3113 vgnd vpwr scs8hd_decap_12
XFILLER_0_1799 vgnd vpwr scs8hd_decap_12
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_3002 vgnd vpwr scs8hd_decap_12
XFILLER_0_869 vgnd vpwr scs8hd_decap_12
XFILLER_2_3923 vgnd vpwr scs8hd_decap_12
XFILLER_9_1780 vgnd vpwr scs8hd_decap_12
XFILLER_5_1611 vgnd vpwr scs8hd_decap_12
XFILLER_1_2209 vgnd vpwr scs8hd_decap_12
XPHY_798 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_787 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_776 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_765 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_754 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_743 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_732 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_721 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_710 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4502 vgnd vpwr scs8hd_decap_12
XFILLER_7_3856 vgnd vpwr scs8hd_decap_12
XFILLER_3_3709 vgnd vpwr scs8hd_decap_12
XFILLER_3_696 vgnd vpwr scs8hd_decap_12
XFILLER_1_2721 vgnd vpwr scs8hd_decap_12
XFILLER_1_4112 vgnd vpwr scs8hd_decap_12
XFILLER_4_1154 vgnd vpwr scs8hd_decap_12
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XFILLER_9_63 vgnd vpwr scs8hd_decap_12
XFILLER_6_4045 vgnd vpwr scs8hd_decap_12
XFILLER_9_1098 vgnd vpwr scs8hd_decap_12
XFILLER_6_3399 vgnd vpwr scs8hd_decap_12
XFILLER_0_2264 vgnd vpwr scs8hd_decap_12
XFILLER_0_1563 vgnd vpwr scs8hd_decap_12
XFILLER_0_2286 vpwr vgnd scs8hd_fill_2
XFILLER_5_928 vgnd vpwr scs8hd_decap_12
XFILLER_5_1452 vgnd vpwr scs8hd_decap_12
XFILLER_0_633 vgnd vpwr scs8hd_decap_12
XFILLER_2_3753 vgnd vpwr scs8hd_decap_12
XFILLER_5_2197 vgnd vpwr scs8hd_decap_12
XFILLER_8_788 vgnd vpwr scs8hd_decap_12
XPHY_595 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_584 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_573 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_562 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_551 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_232 vgnd vpwr scs8hd_decap_12
XPHY_540 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3907 vgnd vpwr scs8hd_decap_12
XFILLER_7_4332 vgnd vpwr scs8hd_decap_12
XFILLER_7_3697 vgnd vpwr scs8hd_decap_12
XFILLER_7_2941 vgnd vpwr scs8hd_decap_12
XFILLER_4_983 vgnd vpwr scs8hd_decap_12
XFILLER_6_1227 vgnd vpwr scs8hd_decap_12
XFILLER_3_3539 vgnd vpwr scs8hd_decap_12
XFILLER_8_2716 vgnd vpwr scs8hd_decap_12
XFILLER_6_3130 vgnd vpwr scs8hd_decap_12
XFILLER_6_2484 vgnd vpwr scs8hd_decap_12
XFILLER_2_2348 vgnd vpwr scs8hd_fill_1
XFILLER_2_2359 vgnd vpwr scs8hd_decap_12
XFILLER_8_3984 vgnd vpwr scs8hd_decap_12
XFILLER_5_769 vgnd vpwr scs8hd_decap_12
XFILLER_4_3826 vgnd vpwr scs8hd_decap_12
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XFILLER_5_1282 vgnd vpwr scs8hd_decap_12
XFILLER_1_964 vgnd vpwr scs8hd_decap_12
XFILLER_2_3594 vgnd vpwr scs8hd_decap_12
XPHY_370 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_1135 vgnd vpwr scs8hd_decap_12
XFILLER_9_4427 vgnd vpwr scs8hd_decap_6
XPHY_392 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_381 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4173 vgnd vpwr scs8hd_decap_12
XFILLER_7_2782 vgnd vpwr scs8hd_decap_12
XFILLER_3_2624 vgnd vpwr scs8hd_decap_12
XPHY_18 vgnd vpwr scs8hd_decap_3
XFILLER_3_1989 vgnd vpwr scs8hd_decap_12
XPHY_29 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_2370 vgnd vpwr scs8hd_decap_3
XFILLER_8_1801 vgnd vpwr scs8hd_decap_12
XFILLER_2_739 vgnd vpwr scs8hd_decap_12
XFILLER_8_2557 vgnd vpwr scs8hd_decap_12
XFILLER_3_3892 vgnd vpwr scs8hd_decap_12
XFILLER_2_1422 vgnd vpwr scs8hd_decap_12
XFILLER_2_2167 vgnd vpwr scs8hd_decap_12
XFILLER_8_4460 vgnd vpwr scs8hd_decap_12
XFILLER_7_2001 vgnd vpwr scs8hd_decap_12
XFILLER_4_4302 vgnd vpwr scs8hd_decap_12
XFILLER_4_3667 vgnd vpwr scs8hd_decap_12
XFILLER_4_2911 vgnd vpwr scs8hd_decap_12
XFILLER_1_794 vgnd vpwr scs8hd_decap_12
XFILLER_2_4070 vgnd vpwr scs8hd_decap_12
XFILLER_7_1355 vgnd vpwr scs8hd_decap_12
XFILLER_3_1208 vgnd vpwr scs8hd_decap_12
XFILLER_9_850 vgnd vpwr scs8hd_decap_12
XFILLER_9_4279 vgnd vpwr scs8hd_decap_12
XFILLER_9_3578 vgnd vpwr scs8hd_decap_12
XFILLER_9_2822 vgnd vpwr scs8hd_decap_12
XFILLER_9_2877 vgnd vpwr scs8hd_decap_6
XFILLER_3_2465 vgnd vpwr scs8hd_decap_12
XFILLER_8_3033 vgnd vpwr scs8hd_decap_12
XFILLER_8_2398 vgnd vpwr scs8hd_decap_12
XFILLER_8_1642 vgnd vpwr scs8hd_decap_12
XFILLER_1_3807 vgnd vpwr scs8hd_decap_12
XFILLER_2_1252 vgnd vpwr scs8hd_decap_12
XFILLER_9_168 vgnd vpwr scs8hd_decap_12
XFILLER_6_886 vgnd vpwr scs8hd_decap_12
XFILLER_5_330 vgnd vpwr scs8hd_decap_12
XFILLER_9_1439 vgnd vpwr scs8hd_decap_12
XFILLER_7_1196 vgnd vpwr scs8hd_decap_12
XFILLER_4_4143 vgnd vpwr scs8hd_decap_12
XFILLER_4_2752 vgnd vpwr scs8hd_decap_12
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_0_2605 vgnd vpwr scs8hd_decap_12
XFILLER_3_1038 vgnd vpwr scs8hd_decap_12
XFILLER_0_1904 vgnd vpwr scs8hd_decap_12
XFILLER_9_4043 vgnd vpwr scs8hd_decap_12
XFILLER_8_190 vgnd vpwr scs8hd_decap_12
XFILLER_9_3342 vgnd vpwr scs8hd_decap_6
XFILLER_9_1951 vpwr vgnd scs8hd_fill_2
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _15_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_2538 vgnd vpwr scs8hd_decap_12
XFILLER_3_1550 vgnd vpwr scs8hd_decap_12
XPHY_903 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_2_300 vgnd vpwr scs8hd_decap_12
XFILLER_8_1483 vgnd vpwr scs8hd_decap_12
XFILLER_5_4441 vgnd vpwr scs8hd_decap_12
XFILLER_5_3795 vgnd vpwr scs8hd_decap_12
XFILLER_4_1325 vgnd vpwr scs8hd_decap_12
XFILLER_3_867 vgnd vpwr scs8hd_decap_12
XFILLER_1_3648 vgnd vpwr scs8hd_decap_12
XFILLER_2_1093 vgnd vpwr scs8hd_decap_12
XFILLER_9_1203 vgnd vpwr scs8hd_decap_6
XFILLER_6_4216 vgnd vpwr scs8hd_decap_12
XFILLER_6_2825 vgnd vpwr scs8hd_decap_12
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
XFILLER_0_2413 vgnd vpwr scs8hd_decap_4
XFILLER_0_3125 vgnd vpwr scs8hd_decap_6
XFILLER_9_3194 vgnd vpwr scs8hd_decap_12
XFILLER_9_1792 vgnd vpwr scs8hd_decap_6
XFILLER_5_3014 vgnd vpwr scs8hd_decap_12
XFILLER_5_2357 vpwr vgnd scs8hd_fill_2
XFILLER_5_1623 vgnd vpwr scs8hd_decap_12
XPHY_711 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_700 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_1391 vgnd vpwr scs8hd_decap_12
XPHY_799 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_788 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_777 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_766 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_755 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_744 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_733 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_722 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_403 vgnd vpwr scs8hd_decap_12
XFILLER_7_3868 vgnd vpwr scs8hd_decap_12
XFILLER_5_4271 vgnd vpwr scs8hd_decap_12
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XFILLER_5_2880 vgnd vpwr scs8hd_decap_12
XFILLER_4_1166 vgnd vpwr scs8hd_decap_12
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_1_2733 vgnd vpwr scs8hd_decap_12
XFILLER_1_3478 vgnd vpwr scs8hd_decap_12
XFILLER_1_4124 vgnd vpwr scs8hd_decap_12
XFILLER_9_75 vgnd vpwr scs8hd_decap_12
XFILLER_9_1055 vgnd vpwr scs8hd_decap_12
XFILLER_9_1022 vgnd vpwr scs8hd_fill_1
XFILLER_9_1000 vpwr vgnd scs8hd_fill_2
XFILLER_6_3301 vgnd vpwr scs8hd_decap_12
XFILLER_6_2655 vgnd vpwr scs8hd_decap_12
XFILLER_6_1910 vgnd vpwr scs8hd_decap_12
XFILLER_2_2508 vgnd vpwr scs8hd_decap_12
XFILLER_0_1520 vgnd vpwr scs8hd_decap_12
XFILLER_0_2276 vgnd vpwr scs8hd_decap_8
XFILLER_1_3990 vgnd vpwr scs8hd_decap_12
XFILLER_0_1575 vgnd vpwr scs8hd_decap_6
XFILLER_2_4411 vgnd vpwr scs8hd_decap_12
XFILLER_1_1306 vgnd vpwr scs8hd_decap_12
XFILLER_0_645 vgnd vpwr scs8hd_decap_6
XFILLER_2_3765 vgnd vpwr scs8hd_decap_12
XPHY_552 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_541 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_530 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3919 vgnd vpwr scs8hd_decap_12
XPHY_596 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_585 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_574 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_563 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4344 vgnd vpwr scs8hd_decap_12
XFILLER_7_2953 vgnd vpwr scs8hd_decap_12
XFILLER_4_995 vgnd vpwr scs8hd_decap_12
XFILLER_6_1239 vgnd vpwr scs8hd_decap_12
XFILLER_1_2563 vgnd vpwr scs8hd_decap_12
XFILLER_8_4119 vgnd vpwr scs8hd_decap_12
XFILLER_8_2728 vgnd vpwr scs8hd_decap_12
XFILLER_6_2496 vgnd vpwr scs8hd_decap_12
XFILLER_6_1740 vgnd vpwr scs8hd_decap_12
XFILLER_2_2327 vpwr vgnd scs8hd_fill_2
XFILLER_0_2040 vgnd vpwr scs8hd_decap_6
XFILLER_9_509 vgnd vpwr scs8hd_decap_12
XFILLER_7_1526 vgnd vpwr scs8hd_decap_12
XFILLER_4_3838 vgnd vpwr scs8hd_decap_12
XFILLER_2_4241 vgnd vpwr scs8hd_decap_12
XFILLER_5_1294 vgnd vpwr scs8hd_decap_12
XFILLER_1_1147 vgnd vpwr scs8hd_decap_12
XFILLER_0_497 vgnd vpwr scs8hd_decap_12
XFILLER_2_2850 vgnd vpwr scs8hd_decap_12
XFILLER_8_520 vgnd vpwr scs8hd_decap_12
XPHY_393 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_382 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_371 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_360 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ top_width_0_height_0__pin_6_ logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[3] vgnd vpwr scs8hd_ebufn_1
XFILLER_7_4185 vgnd vpwr scs8hd_decap_12
XFILLER_7_2794 vgnd vpwr scs8hd_decap_12
XFILLER_6_1069 vgnd vpwr scs8hd_decap_12
XFILLER_3_4027 vgnd vpwr scs8hd_decap_12
XFILLER_3_2636 vgnd vpwr scs8hd_decap_12
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_8_3204 vgnd vpwr scs8hd_decap_12
XFILLER_8_2569 vgnd vpwr scs8hd_decap_12
XFILLER_8_1813 vgnd vpwr scs8hd_decap_12
XFILLER_8_1846 vgnd vpwr scs8hd_decap_12
XFILLER_6_1581 vgnd vpwr scs8hd_decap_12
XFILLER_2_2179 vgnd vpwr scs8hd_decap_12
XFILLER_0_1191 vgnd vpwr scs8hd_decap_12
XFILLER_8_4472 vgnd vpwr scs8hd_decap_12
XFILLER_5_501 vgnd vpwr scs8hd_decap_12
XFILLER_7_1367 vgnd vpwr scs8hd_decap_12
XFILLER_4_4314 vgnd vpwr scs8hd_decap_12
XFILLER_4_3679 vgnd vpwr scs8hd_decap_12
XFILLER_4_2923 vgnd vpwr scs8hd_decap_12
XFILLER_0_261 vgnd vpwr scs8hd_decap_12
XFILLER_2_4082 vgnd vpwr scs8hd_decap_12
XFILLER_2_2691 vgnd vpwr scs8hd_decap_12
XFILLER_9_862 vgnd vpwr scs8hd_decap_6
XFILLER_8_361 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3535 vgnd vpwr scs8hd_decap_12
XFILLER_9_2834 vgnd vpwr scs8hd_decap_12
XFILLER_7_3270 vgnd vpwr scs8hd_decap_12
XFILLER_5_2709 vgnd vpwr scs8hd_decap_12
XFILLER_3_3112 vgnd vpwr scs8hd_decap_12
XFILLER_3_2477 vgnd vpwr scs8hd_decap_12
XFILLER_3_1721 vgnd vpwr scs8hd_decap_12
XFILLER_8_3045 vgnd vpwr scs8hd_decap_12
XFILLER_8_2333 vgnd vpwr scs8hd_decap_12
XFILLER_8_1654 vgnd vpwr scs8hd_decap_12
XFILLER_5_3966 vgnd vpwr scs8hd_decap_12
XFILLER_3_4380 vgnd vpwr scs8hd_decap_12
XFILLER_1_3819 vgnd vpwr scs8hd_decap_12
XFILLER_2_1264 vgnd vpwr scs8hd_decap_12
XFILLER_9_125 vgnd vpwr scs8hd_decap_12
XFILLER_6_898 vgnd vpwr scs8hd_decap_12
XFILLER_5_342 vgnd vpwr scs8hd_decap_12
XFILLER_4_4155 vgnd vpwr scs8hd_decap_12
XFILLER_4_2764 vgnd vpwr scs8hd_decap_12
XFILLER_0_2617 vgnd vpwr scs8hd_decap_12
XFILLER_0_3318 vgnd vpwr scs8hd_decap_12
XFILLER_0_1916 vgnd vpwr scs8hd_decap_6
XFILLER_9_4055 vgnd vpwr scs8hd_decap_6
XFILLER_9_4000 vgnd vpwr scs8hd_decap_12
XFILLER_9_1985 vgnd vpwr scs8hd_decap_12
XFILLER_0_4520 vgnd vpwr scs8hd_decap_6
XFILLER_3_1562 vgnd vpwr scs8hd_decap_12
XPHY_904 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XFILLER_8_2130 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_879 vgnd vpwr scs8hd_decap_12
XFILLER_2_312 vgnd vpwr scs8hd_decap_12
XFILLER_4_1337 vgnd vpwr scs8hd_decap_12
XFILLER_1_2904 vgnd vpwr scs8hd_decap_12
XFILLER_6_4228 vgnd vpwr scs8hd_decap_12
XFILLER_4_3240 vgnd vpwr scs8hd_decap_12
XFILLER_4_2594 vgnd vpwr scs8hd_decap_12
XFILLER_0_1768 vgnd vpwr scs8hd_decap_12
XFILLER_9_2450 vgnd vpwr scs8hd_decap_12
XFILLER_5_3026 vgnd vpwr scs8hd_decap_12
XFILLER_5_2336 vpwr vgnd scs8hd_fill_2
XFILLER_5_2314 vpwr vgnd scs8hd_fill_2
XFILLER_5_1635 vgnd vpwr scs8hd_decap_12
XFILLER_0_838 vgnd vpwr scs8hd_decap_12
XFILLER_0_4372 vgnd vpwr scs8hd_decap_12
XFILLER_2_3936 vgnd vpwr scs8hd_decap_12
XPHY_745 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_734 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_723 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_712 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_701 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_2970 vgnd vpwr scs8hd_decap_6
XFILLER_0_3671 vgnd vpwr scs8hd_decap_12
XPHY_789 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_778 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_767 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_756 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4515 vgnd vpwr scs8hd_decap_12
XFILLER_7_415 vgnd vpwr scs8hd_decap_12
XFILLER_5_4283 vgnd vpwr scs8hd_decap_12
XFILLER_1_4136 vgnd vpwr scs8hd_decap_12
XFILLER_5_2892 vgnd vpwr scs8hd_decap_12
XFILLER_4_1178 vgnd vpwr scs8hd_decap_12
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_9_87 vgnd vpwr scs8hd_decap_6
XFILLER_9_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_4058 vgnd vpwr scs8hd_decap_12
XFILLER_6_3313 vgnd vpwr scs8hd_decap_12
XFILLER_9_1067 vgnd vpwr scs8hd_decap_12
XFILLER_6_2667 vgnd vpwr scs8hd_decap_12
XFILLER_4_2380 vgnd vpwr scs8hd_decap_4
XFILLER_0_1532 vgnd vpwr scs8hd_decap_12
XFILLER_0_2233 vgnd vpwr scs8hd_decap_12
XFILLER_0_2299 vgnd vpwr scs8hd_decap_3
XFILLER_6_4570 vgnd vpwr scs8hd_decap_8
XFILLER_5_2111 vgnd vpwr scs8hd_decap_12
XFILLER_0_602 vgnd vpwr scs8hd_decap_12
XFILLER_5_1465 vgnd vpwr scs8hd_decap_12
XFILLER_1_1318 vgnd vpwr scs8hd_decap_12
XFILLER_2_3777 vgnd vpwr scs8hd_decap_12
XPHY_586 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_575 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_564 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_553 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_542 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_531 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_520 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4356 vgnd vpwr scs8hd_decap_12
XFILLER_7_3600 vgnd vpwr scs8hd_decap_12
XPHY_597 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
XFILLER_7_2965 vgnd vpwr scs8hd_decap_12
XFILLER_3_2807 vgnd vpwr scs8hd_decap_12
XFILLER_3_440 vgnd vpwr scs8hd_decap_12
XFILLER_1_3221 vgnd vpwr scs8hd_decap_12
XFILLER_1_2575 vgnd vpwr scs8hd_decap_12
XFILLER_6_3143 vgnd vpwr scs8hd_decap_12
XFILLER_6_1752 vgnd vpwr scs8hd_decap_12
XFILLER_2_1605 vgnd vpwr scs8hd_decap_12
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_3997 vgnd vpwr scs8hd_decap_12
XFILLER_7_1538 vgnd vpwr scs8hd_decap_12
XFILLER_2_4253 vgnd vpwr scs8hd_decap_12
XFILLER_1_977 vgnd vpwr scs8hd_decap_12
XFILLER_2_2862 vgnd vpwr scs8hd_decap_12
XFILLER_8_532 vgnd vpwr scs8hd_decap_12
XPHY_394 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_383 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_372 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_361 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_350 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_4197 vgnd vpwr scs8hd_decap_12
XFILLER_7_3441 vgnd vpwr scs8hd_decap_12
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_4039 vgnd vpwr scs8hd_decap_12
XFILLER_3_281 vgnd vpwr scs8hd_decap_12
XFILLER_3_2648 vgnd vpwr scs8hd_decap_12
XFILLER_1_3051 vgnd vpwr scs8hd_decap_12
XFILLER_1_1660 vgnd vpwr scs8hd_decap_12
XFILLER_1_2350 vpwr vgnd scs8hd_fill_2
XFILLER_8_3216 vgnd vpwr scs8hd_decap_12
XFILLER_8_1858 vgnd vpwr scs8hd_decap_3
XFILLER_8_1825 vgnd vpwr scs8hd_decap_12
XFILLER_3_4551 vgnd vpwr scs8hd_decap_12
XFILLER_6_1593 vgnd vpwr scs8hd_decap_12
XFILLER_2_1435 vgnd vpwr scs8hd_decap_12
XFILLER_5_513 vgnd vpwr scs8hd_decap_12
XFILLER_4_4326 vgnd vpwr scs8hd_decap_12
XFILLER_7_2014 vgnd vpwr scs8hd_decap_12
XFILLER_7_1379 vgnd vpwr scs8hd_decap_12
XFILLER_4_2935 vgnd vpwr scs8hd_decap_12
XFILLER_0_273 vgnd vpwr scs8hd_decap_6
XFILLER_2_4094 vgnd vpwr scs8hd_decap_12
XFILLER_9_4248 vgnd vpwr scs8hd_decap_12
XFILLER_8_373 vgnd vpwr scs8hd_decap_12
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3547 vgnd vpwr scs8hd_decap_12
XFILLER_9_2846 vgnd vpwr scs8hd_decap_6
XFILLER_7_3282 vgnd vpwr scs8hd_decap_12
XFILLER_3_3124 vgnd vpwr scs8hd_decap_12
.ends

