magic
tech EFS8A
magscale 1 2
timestamp 1604337443
<< locali >>
rect 3341 21879 3375 22049
rect 12081 20247 12115 20349
rect 14657 20247 14691 20349
rect 4905 17119 4939 17289
rect 6745 14263 6779 14433
rect 8861 10999 8895 11101
rect 12449 10455 12483 10625
rect 8861 10047 8895 10149
rect 6469 9367 6503 9605
rect 3525 8347 3559 8517
rect 7941 8279 7975 8517
rect 13645 7191 13679 7293
rect 6561 2295 6595 2533
<< viali >>
rect 4721 25381 4755 25415
rect 4905 25381 4939 25415
rect 8125 25381 8159 25415
rect 11345 25381 11379 25415
rect 4997 25313 5031 25347
rect 7941 25313 7975 25347
rect 11161 25313 11195 25347
rect 13921 25313 13955 25347
rect 8217 25245 8251 25279
rect 11437 25245 11471 25279
rect 7297 25177 7331 25211
rect 4445 25109 4479 25143
rect 7665 25109 7699 25143
rect 10149 25109 10183 25143
rect 10885 25109 10919 25143
rect 14105 25109 14139 25143
rect 5089 24905 5123 24939
rect 2053 24837 2087 24871
rect 3525 24837 3559 24871
rect 8677 24837 8711 24871
rect 1593 24769 1627 24803
rect 4537 24769 4571 24803
rect 5733 24769 5767 24803
rect 7757 24769 7791 24803
rect 8953 24769 8987 24803
rect 9965 24769 9999 24803
rect 10609 24769 10643 24803
rect 3801 24701 3835 24735
rect 6653 24701 6687 24735
rect 7849 24701 7883 24735
rect 13001 24701 13035 24735
rect 13277 24701 13311 24735
rect 14289 24701 14323 24735
rect 14841 24701 14875 24735
rect 15393 24701 15427 24735
rect 3157 24633 3191 24667
rect 4629 24633 4663 24667
rect 5365 24633 5399 24667
rect 7757 24633 7791 24667
rect 10701 24633 10735 24667
rect 4067 24565 4101 24599
rect 4537 24565 4571 24599
rect 7021 24565 7055 24599
rect 7287 24565 7321 24599
rect 8309 24565 8343 24599
rect 10131 24565 10165 24599
rect 10609 24565 10643 24599
rect 11069 24565 11103 24599
rect 11529 24565 11563 24599
rect 11897 24565 11931 24599
rect 12817 24565 12851 24599
rect 14013 24565 14047 24599
rect 14473 24565 14507 24599
rect 15577 24565 15611 24599
rect 16037 24565 16071 24599
rect 2881 24361 2915 24395
rect 8585 24361 8619 24395
rect 10057 24361 10091 24395
rect 15485 24361 15519 24395
rect 16589 24361 16623 24395
rect 17693 24361 17727 24395
rect 19717 24361 19751 24395
rect 1746 24293 1780 24327
rect 4905 24293 4939 24327
rect 6561 24293 6595 24327
rect 8125 24293 8159 24327
rect 8217 24293 8251 24327
rect 11060 24293 11094 24327
rect 1501 24225 1535 24259
rect 4997 24225 5031 24259
rect 6653 24225 6687 24259
rect 7113 24225 7147 24259
rect 13921 24225 13955 24259
rect 14197 24225 14231 24259
rect 15301 24225 15335 24259
rect 16405 24225 16439 24259
rect 17509 24225 17543 24259
rect 19533 24225 19567 24259
rect 4905 24157 4939 24191
rect 6469 24157 6503 24191
rect 8033 24157 8067 24191
rect 10793 24157 10827 24191
rect 6101 24089 6135 24123
rect 7389 24089 7423 24123
rect 7665 24089 7699 24123
rect 4445 24021 4479 24055
rect 5917 24021 5951 24055
rect 12173 24021 12207 24055
rect 1501 23817 1535 23851
rect 4353 23817 4387 23851
rect 6469 23817 6503 23851
rect 8309 23817 8343 23851
rect 11345 23817 11379 23851
rect 12173 23817 12207 23851
rect 15301 23817 15335 23851
rect 16405 23817 16439 23851
rect 17049 23817 17083 23851
rect 17785 23817 17819 23851
rect 18705 23817 18739 23851
rect 19809 23817 19843 23851
rect 22017 23817 22051 23851
rect 6009 23749 6043 23783
rect 6929 23749 6963 23783
rect 20913 23749 20947 23783
rect 2053 23681 2087 23715
rect 8401 23681 8435 23715
rect 10885 23681 10919 23715
rect 12449 23681 12483 23715
rect 15853 23681 15887 23715
rect 1777 23613 1811 23647
rect 2973 23613 3007 23647
rect 3229 23613 3263 23647
rect 4997 23613 5031 23647
rect 7205 23613 7239 23647
rect 8668 23613 8702 23647
rect 15577 23613 15611 23647
rect 16865 23613 16899 23647
rect 17417 23613 17451 23647
rect 18521 23613 18555 23647
rect 19073 23613 19107 23647
rect 19625 23613 19659 23647
rect 20729 23613 20763 23647
rect 21281 23613 21315 23647
rect 21833 23613 21867 23647
rect 22385 23613 22419 23647
rect 2513 23545 2547 23579
rect 2881 23545 2915 23579
rect 5365 23545 5399 23579
rect 7389 23545 7423 23579
rect 7481 23545 7515 23579
rect 11805 23545 11839 23579
rect 12694 23545 12728 23579
rect 1961 23477 1995 23511
rect 5733 23477 5767 23511
rect 7849 23477 7883 23511
rect 9781 23477 9815 23511
rect 10701 23477 10735 23511
rect 13829 23477 13863 23511
rect 14381 23477 14415 23511
rect 14933 23477 14967 23511
rect 19533 23477 19567 23511
rect 20177 23477 20211 23511
rect 1685 23273 1719 23307
rect 1961 23273 1995 23307
rect 5089 23273 5123 23307
rect 6101 23273 6135 23307
rect 6929 23273 6963 23307
rect 8493 23273 8527 23307
rect 10333 23273 10367 23307
rect 11069 23273 11103 23307
rect 17049 23273 17083 23307
rect 18153 23273 18187 23307
rect 22017 23273 22051 23307
rect 2973 23205 3007 23239
rect 3065 23205 3099 23239
rect 3433 23205 3467 23239
rect 5917 23205 5951 23239
rect 12633 23205 12667 23239
rect 12725 23205 12759 23239
rect 13185 23205 13219 23239
rect 14197 23205 14231 23239
rect 15853 23205 15887 23239
rect 4445 23137 4479 23171
rect 7113 23137 7147 23171
rect 7380 23137 7414 23171
rect 10057 23137 10091 23171
rect 10885 23137 10919 23171
rect 12449 23137 12483 23171
rect 13553 23137 13587 23171
rect 14289 23137 14323 23171
rect 16865 23137 16899 23171
rect 17969 23137 18003 23171
rect 21833 23137 21867 23171
rect 2973 23069 3007 23103
rect 6193 23069 6227 23103
rect 11161 23069 11195 23103
rect 14197 23069 14231 23103
rect 15853 23069 15887 23103
rect 15945 23069 15979 23103
rect 2513 23001 2547 23035
rect 4721 23001 4755 23035
rect 10609 23001 10643 23035
rect 12173 23001 12207 23035
rect 5641 22933 5675 22967
rect 13737 22933 13771 22967
rect 15393 22933 15427 22967
rect 2237 22729 2271 22763
rect 4261 22729 4295 22763
rect 5825 22729 5859 22763
rect 6193 22729 6227 22763
rect 7113 22729 7147 22763
rect 7297 22729 7331 22763
rect 8309 22729 8343 22763
rect 9781 22729 9815 22763
rect 10057 22729 10091 22763
rect 11069 22729 11103 22763
rect 11437 22729 11471 22763
rect 13277 22729 13311 22763
rect 15117 22729 15151 22763
rect 16405 22729 16439 22763
rect 18245 22729 18279 22763
rect 21833 22729 21867 22763
rect 4905 22661 4939 22695
rect 6653 22661 6687 22695
rect 11805 22661 11839 22695
rect 12081 22661 12115 22695
rect 13553 22661 13587 22695
rect 7849 22593 7883 22627
rect 10609 22593 10643 22627
rect 13737 22593 13771 22627
rect 1869 22525 1903 22559
rect 2329 22525 2363 22559
rect 5181 22525 5215 22559
rect 7573 22525 7607 22559
rect 8585 22525 8619 22559
rect 10333 22525 10367 22559
rect 12449 22525 12483 22559
rect 16221 22525 16255 22559
rect 2596 22457 2630 22491
rect 4721 22457 4755 22491
rect 5457 22457 5491 22491
rect 7757 22457 7791 22491
rect 9505 22457 9539 22491
rect 10517 22457 10551 22491
rect 12725 22457 12759 22491
rect 14004 22457 14038 22491
rect 15761 22457 15795 22491
rect 3709 22389 3743 22423
rect 5365 22389 5399 22423
rect 16037 22389 16071 22423
rect 16865 22389 16899 22423
rect 1961 22185 1995 22219
rect 2973 22185 3007 22219
rect 4261 22185 4295 22219
rect 8033 22185 8067 22219
rect 9965 22185 9999 22219
rect 13737 22185 13771 22219
rect 14197 22185 14231 22219
rect 15025 22185 15059 22219
rect 15853 22185 15887 22219
rect 16313 22185 16347 22219
rect 5641 22117 5675 22151
rect 7205 22117 7239 22151
rect 2329 22049 2363 22083
rect 3341 22049 3375 22083
rect 3525 22049 3559 22083
rect 7021 22049 7055 22083
rect 7757 22049 7791 22083
rect 10517 22049 10551 22083
rect 10957 22049 10991 22083
rect 12633 22049 12667 22083
rect 13553 22049 13587 22083
rect 15669 22049 15703 22083
rect 16865 22049 16899 22083
rect 2973 21981 3007 22015
rect 3065 21981 3099 22015
rect 2513 21913 2547 21947
rect 5641 21981 5675 22015
rect 5733 21981 5767 22015
rect 7297 21981 7331 22015
rect 10701 21981 10735 22015
rect 13829 21981 13863 22015
rect 15945 21981 15979 22015
rect 3801 21913 3835 21947
rect 5181 21913 5215 21947
rect 12081 21913 12115 21947
rect 17049 21913 17083 21947
rect 3341 21845 3375 21879
rect 4997 21845 5031 21879
rect 6745 21845 6779 21879
rect 9045 21845 9079 21879
rect 9413 21845 9447 21879
rect 13277 21845 13311 21879
rect 15393 21845 15427 21879
rect 5549 21641 5583 21675
rect 6285 21641 6319 21675
rect 8309 21641 8343 21675
rect 9137 21641 9171 21675
rect 10701 21641 10735 21675
rect 11897 21641 11931 21675
rect 12541 21641 12575 21675
rect 13829 21641 13863 21675
rect 14473 21641 14507 21675
rect 15025 21641 15059 21675
rect 16957 21641 16991 21675
rect 18337 21641 18371 21675
rect 2053 21573 2087 21607
rect 6929 21573 6963 21607
rect 13461 21573 13495 21607
rect 2513 21505 2547 21539
rect 11253 21505 11287 21539
rect 1869 21437 1903 21471
rect 2605 21437 2639 21471
rect 3433 21437 3467 21471
rect 3525 21437 3559 21471
rect 3792 21437 3826 21471
rect 7481 21437 7515 21471
rect 7849 21437 7883 21471
rect 8953 21437 8987 21471
rect 9689 21437 9723 21471
rect 10057 21437 10091 21471
rect 13093 21437 13127 21471
rect 15301 21437 15335 21471
rect 16313 21437 16347 21471
rect 18153 21437 18187 21471
rect 18705 21437 18739 21471
rect 3065 21369 3099 21403
rect 7205 21369 7239 21403
rect 9413 21369 9447 21403
rect 10977 21369 11011 21403
rect 12817 21369 12851 21403
rect 14841 21369 14875 21403
rect 15577 21369 15611 21403
rect 16497 21369 16531 21403
rect 2513 21301 2547 21335
rect 4905 21301 4939 21335
rect 5917 21301 5951 21335
rect 6653 21301 6687 21335
rect 7389 21301 7423 21335
rect 9597 21301 9631 21335
rect 10517 21301 10551 21335
rect 11161 21301 11195 21335
rect 12173 21301 12207 21335
rect 13001 21301 13035 21335
rect 15485 21301 15519 21335
rect 16037 21301 16071 21335
rect 2421 21097 2455 21131
rect 3617 21097 3651 21131
rect 4261 21097 4295 21131
rect 4721 21097 4755 21131
rect 6285 21097 6319 21131
rect 6929 21097 6963 21131
rect 8401 21097 8435 21131
rect 11069 21097 11103 21131
rect 12541 21097 12575 21131
rect 13185 21097 13219 21131
rect 15025 21097 15059 21131
rect 15577 21097 15611 21131
rect 17049 21097 17083 21131
rect 21097 21097 21131 21131
rect 5172 21029 5206 21063
rect 7757 21029 7791 21063
rect 7941 21029 7975 21063
rect 14197 21029 14231 21063
rect 14289 21029 14323 21063
rect 4905 20961 4939 20995
rect 9689 20961 9723 20995
rect 9956 20961 9990 20995
rect 14013 20961 14047 20995
rect 15936 20961 15970 20995
rect 20913 20961 20947 20995
rect 2329 20893 2363 20927
rect 2513 20893 2547 20927
rect 8033 20893 8067 20927
rect 15669 20893 15703 20927
rect 7481 20825 7515 20859
rect 1685 20757 1719 20791
rect 1961 20757 1995 20791
rect 3157 20757 3191 20791
rect 7297 20757 7331 20791
rect 9413 20757 9447 20791
rect 12909 20757 12943 20791
rect 13737 20757 13771 20791
rect 1593 20553 1627 20587
rect 2513 20553 2547 20587
rect 2973 20553 3007 20587
rect 4537 20553 4571 20587
rect 6285 20553 6319 20587
rect 6653 20553 6687 20587
rect 8769 20553 8803 20587
rect 9137 20553 9171 20587
rect 9413 20553 9447 20587
rect 10793 20553 10827 20587
rect 11161 20553 11195 20587
rect 13645 20553 13679 20587
rect 14105 20553 14139 20587
rect 14381 20553 14415 20587
rect 3157 20485 3191 20519
rect 4721 20485 4755 20519
rect 12541 20485 12575 20519
rect 3617 20417 3651 20451
rect 5181 20417 5215 20451
rect 9965 20417 9999 20451
rect 13001 20417 13035 20451
rect 18337 20417 18371 20451
rect 1869 20349 1903 20383
rect 3709 20349 3743 20383
rect 5733 20349 5767 20383
rect 6837 20349 6871 20383
rect 12081 20349 12115 20383
rect 13093 20349 13127 20383
rect 14657 20349 14691 20383
rect 14933 20349 14967 20383
rect 18061 20349 18095 20383
rect 18797 20349 18831 20383
rect 2145 20281 2179 20315
rect 3617 20281 3651 20315
rect 5273 20281 5307 20315
rect 7082 20281 7116 20315
rect 9689 20281 9723 20315
rect 13001 20281 13035 20315
rect 15178 20281 15212 20315
rect 2053 20213 2087 20247
rect 4169 20213 4203 20247
rect 5181 20213 5215 20247
rect 8217 20213 8251 20247
rect 9873 20213 9907 20247
rect 10425 20213 10459 20247
rect 11805 20213 11839 20247
rect 12081 20213 12115 20247
rect 12173 20213 12207 20247
rect 14657 20213 14691 20247
rect 14749 20213 14783 20247
rect 16313 20213 16347 20247
rect 20913 20213 20947 20247
rect 1869 20009 1903 20043
rect 2329 20009 2363 20043
rect 3157 20009 3191 20043
rect 5273 20009 5307 20043
rect 6561 20009 6595 20043
rect 6929 20009 6963 20043
rect 8493 20009 8527 20043
rect 10149 20009 10183 20043
rect 10793 20009 10827 20043
rect 13553 20009 13587 20043
rect 15669 20009 15703 20043
rect 3433 19941 3467 19975
rect 4721 19941 4755 19975
rect 14197 19941 14231 19975
rect 14289 19941 14323 19975
rect 14933 19941 14967 19975
rect 16488 19941 16522 19975
rect 19441 19941 19475 19975
rect 7113 19873 7147 19907
rect 7380 19873 7414 19907
rect 11161 19873 11195 19907
rect 11428 19873 11462 19907
rect 14013 19873 14047 19907
rect 16221 19873 16255 19907
rect 19165 19873 19199 19907
rect 4629 19805 4663 19839
rect 4813 19805 4847 19839
rect 9689 19805 9723 19839
rect 17601 19737 17635 19771
rect 1685 19669 1719 19703
rect 2697 19669 2731 19703
rect 3801 19669 3835 19703
rect 4261 19669 4295 19703
rect 9413 19669 9447 19703
rect 12541 19669 12575 19703
rect 13737 19669 13771 19703
rect 16037 19669 16071 19703
rect 1685 19465 1719 19499
rect 5181 19465 5215 19499
rect 7849 19465 7883 19499
rect 9045 19465 9079 19499
rect 10885 19465 10919 19499
rect 14381 19465 14415 19499
rect 15025 19465 15059 19499
rect 16313 19465 16347 19499
rect 16589 19465 16623 19499
rect 2329 19397 2363 19431
rect 4813 19329 4847 19363
rect 9505 19329 9539 19363
rect 4169 19261 4203 19295
rect 5641 19261 5675 19295
rect 6285 19261 6319 19295
rect 7205 19261 7239 19295
rect 10609 19261 10643 19295
rect 12449 19261 12483 19295
rect 15301 19261 15335 19295
rect 16957 19261 16991 19295
rect 22293 19261 22327 19295
rect 22845 19261 22879 19295
rect 2605 19193 2639 19227
rect 2881 19193 2915 19227
rect 3875 19193 3909 19227
rect 4353 19193 4387 19227
rect 4445 19193 4479 19227
rect 6653 19193 6687 19227
rect 7389 19193 7423 19227
rect 7481 19193 7515 19227
rect 8493 19193 8527 19227
rect 9597 19193 9631 19227
rect 10333 19193 10367 19227
rect 11161 19193 11195 19227
rect 11437 19193 11471 19227
rect 12716 19193 12750 19227
rect 15485 19193 15519 19227
rect 15577 19193 15611 19227
rect 2145 19125 2179 19159
rect 2789 19125 2823 19159
rect 3341 19125 3375 19159
rect 3709 19125 3743 19159
rect 6919 19125 6953 19159
rect 8769 19125 8803 19159
rect 9505 19125 9539 19159
rect 11345 19125 11379 19159
rect 11897 19125 11931 19159
rect 12265 19125 12299 19159
rect 13829 19125 13863 19159
rect 14749 19125 14783 19159
rect 19165 19125 19199 19159
rect 22477 19125 22511 19159
rect 2329 18921 2363 18955
rect 3893 18921 3927 18955
rect 5457 18921 5491 18955
rect 7573 18921 7607 18955
rect 9045 18921 9079 18955
rect 10885 18921 10919 18955
rect 15025 18921 15059 18955
rect 16313 18921 16347 18955
rect 2973 18853 3007 18887
rect 7113 18853 7147 18887
rect 10241 18853 10275 18887
rect 11253 18853 11287 18887
rect 15853 18853 15887 18887
rect 15945 18853 15979 18887
rect 2789 18785 2823 18819
rect 4333 18785 4367 18819
rect 6469 18785 6503 18819
rect 6929 18785 6963 18819
rect 10333 18785 10367 18819
rect 12992 18785 13026 18819
rect 15669 18785 15703 18819
rect 3065 18717 3099 18751
rect 4077 18717 4111 18751
rect 7205 18717 7239 18751
rect 10241 18717 10275 18751
rect 12725 18717 12759 18751
rect 2513 18649 2547 18683
rect 9781 18649 9815 18683
rect 6653 18581 6687 18615
rect 11713 18581 11747 18615
rect 12541 18581 12575 18615
rect 14105 18581 14139 18615
rect 15393 18581 15427 18615
rect 2053 18377 2087 18411
rect 4537 18377 4571 18411
rect 5089 18377 5123 18411
rect 8217 18377 8251 18411
rect 11897 18377 11931 18411
rect 12541 18377 12575 18411
rect 14105 18377 14139 18411
rect 15025 18377 15059 18411
rect 16957 18377 16991 18411
rect 2973 18309 3007 18343
rect 6929 18309 6963 18343
rect 9321 18309 9355 18343
rect 10885 18309 10919 18343
rect 15669 18309 15703 18343
rect 2145 18241 2179 18275
rect 3157 18241 3191 18275
rect 6285 18241 6319 18275
rect 7481 18241 7515 18275
rect 7849 18241 7883 18275
rect 9689 18241 9723 18275
rect 11345 18241 11379 18275
rect 13093 18241 13127 18275
rect 14565 18241 14599 18275
rect 16221 18241 16255 18275
rect 21557 18241 21591 18275
rect 2697 18173 2731 18207
rect 3424 18173 3458 18207
rect 5641 18173 5675 18207
rect 8769 18173 8803 18207
rect 9873 18173 9907 18207
rect 16589 18173 16623 18207
rect 21281 18173 21315 18207
rect 22017 18173 22051 18207
rect 1685 18105 1719 18139
rect 5733 18105 5767 18139
rect 6653 18105 6687 18139
rect 7205 18105 7239 18139
rect 7389 18105 7423 18139
rect 10241 18105 10275 18139
rect 10701 18105 10735 18139
rect 11437 18105 11471 18139
rect 12817 18105 12851 18139
rect 14565 18105 14599 18139
rect 14657 18105 14691 18139
rect 15393 18105 15427 18139
rect 15945 18105 15979 18139
rect 16129 18105 16163 18139
rect 9045 18037 9079 18071
rect 9781 18037 9815 18071
rect 11345 18037 11379 18071
rect 12173 18037 12207 18071
rect 13001 18037 13035 18071
rect 13461 18037 13495 18071
rect 13921 18037 13955 18071
rect 2329 17833 2363 17867
rect 4261 17833 4295 17867
rect 6469 17833 6503 17867
rect 7389 17833 7423 17867
rect 8585 17833 8619 17867
rect 9229 17833 9263 17867
rect 10333 17833 10367 17867
rect 10783 17833 10817 17867
rect 11713 17833 11747 17867
rect 12081 17833 12115 17867
rect 13737 17833 13771 17867
rect 14197 17833 14231 17867
rect 14565 17833 14599 17867
rect 15117 17833 15151 17867
rect 2973 17765 3007 17799
rect 3065 17765 3099 17799
rect 5356 17765 5390 17799
rect 7113 17765 7147 17799
rect 7941 17765 7975 17799
rect 8125 17765 8159 17799
rect 11253 17765 11287 17799
rect 12541 17765 12575 17799
rect 13277 17765 13311 17799
rect 15853 17765 15887 17799
rect 15945 17765 15979 17799
rect 16313 17765 16347 17799
rect 13369 17697 13403 17731
rect 15669 17697 15703 17731
rect 2881 17629 2915 17663
rect 5089 17629 5123 17663
rect 8217 17629 8251 17663
rect 11253 17629 11287 17663
rect 11345 17629 11379 17663
rect 13185 17629 13219 17663
rect 2513 17561 2547 17595
rect 7665 17561 7699 17595
rect 15393 17561 15427 17595
rect 9965 17493 9999 17527
rect 12817 17493 12851 17527
rect 2513 17289 2547 17323
rect 2881 17289 2915 17323
rect 3157 17289 3191 17323
rect 4905 17289 4939 17323
rect 4997 17289 5031 17323
rect 5273 17289 5307 17323
rect 6285 17289 6319 17323
rect 8769 17289 8803 17323
rect 9137 17289 9171 17323
rect 10885 17289 10919 17323
rect 12265 17289 12299 17323
rect 14473 17289 14507 17323
rect 16037 17289 16071 17323
rect 16405 17289 16439 17323
rect 4353 17221 4387 17255
rect 4629 17153 4663 17187
rect 10701 17221 10735 17255
rect 5825 17153 5859 17187
rect 4905 17085 4939 17119
rect 5549 17085 5583 17119
rect 6561 17085 6595 17119
rect 6837 17085 6871 17119
rect 7093 17085 7127 17119
rect 9965 17085 9999 17119
rect 11805 17085 11839 17119
rect 13093 17085 13127 17119
rect 13360 17085 13394 17119
rect 11161 17017 11195 17051
rect 11437 17017 11471 17051
rect 1685 16949 1719 16983
rect 5733 16949 5767 16983
rect 8217 16949 8251 16983
rect 10241 16949 10275 16983
rect 11345 16949 11379 16983
rect 12909 16949 12943 16983
rect 15301 16949 15335 16983
rect 15577 16949 15611 16983
rect 5181 16745 5215 16779
rect 8493 16745 8527 16779
rect 10885 16745 10919 16779
rect 11161 16745 11195 16779
rect 13277 16745 13311 16779
rect 15853 16745 15887 16779
rect 5917 16677 5951 16711
rect 6101 16677 6135 16711
rect 7380 16677 7414 16711
rect 10241 16677 10275 16711
rect 10333 16677 10367 16711
rect 12142 16677 12176 16711
rect 13921 16677 13955 16711
rect 2421 16609 2455 16643
rect 7113 16609 7147 16643
rect 9763 16609 9797 16643
rect 15945 16609 15979 16643
rect 6193 16541 6227 16575
rect 10149 16541 10183 16575
rect 11897 16541 11931 16575
rect 15853 16541 15887 16575
rect 1961 16473 1995 16507
rect 1593 16405 1627 16439
rect 4905 16405 4939 16439
rect 5641 16405 5675 16439
rect 6929 16405 6963 16439
rect 15393 16405 15427 16439
rect 1869 16201 1903 16235
rect 4997 16201 5031 16235
rect 6929 16201 6963 16235
rect 11069 16201 11103 16235
rect 13093 16201 13127 16235
rect 16221 16201 16255 16235
rect 2053 16133 2087 16167
rect 5273 16133 5307 16167
rect 7849 16133 7883 16167
rect 8493 16133 8527 16167
rect 10609 16133 10643 16167
rect 13369 16133 13403 16167
rect 2421 16065 2455 16099
rect 5733 16065 5767 16099
rect 7481 16065 7515 16099
rect 8677 16065 8711 16099
rect 11161 16065 11195 16099
rect 15853 16065 15887 16099
rect 2605 15997 2639 16031
rect 4721 15997 4755 16031
rect 8933 15997 8967 16031
rect 13921 15997 13955 16031
rect 14177 15997 14211 16031
rect 16681 15997 16715 16031
rect 17417 15997 17451 16031
rect 3433 15929 3467 15963
rect 5733 15929 5767 15963
rect 5825 15929 5859 15963
rect 7205 15929 7239 15963
rect 7389 15929 7423 15963
rect 11989 15929 12023 15963
rect 16957 15929 16991 15963
rect 2513 15861 2547 15895
rect 3065 15861 3099 15895
rect 3525 15861 3559 15895
rect 4353 15861 4387 15895
rect 6193 15861 6227 15895
rect 6561 15861 6595 15895
rect 10057 15861 10091 15895
rect 12725 15861 12759 15895
rect 13829 15861 13863 15895
rect 15301 15861 15335 15895
rect 1961 15657 1995 15691
rect 5273 15657 5307 15691
rect 7389 15657 7423 15691
rect 8953 15657 8987 15691
rect 11621 15657 11655 15691
rect 13921 15657 13955 15691
rect 8493 15589 8527 15623
rect 15853 15589 15887 15623
rect 16939 15589 16973 15623
rect 17233 15589 17267 15623
rect 17417 15589 17451 15623
rect 1409 15521 1443 15555
rect 2513 15521 2547 15555
rect 4445 15521 4479 15555
rect 5457 15521 5491 15555
rect 5724 15521 5758 15555
rect 8309 15521 8343 15555
rect 9689 15521 9723 15555
rect 9956 15521 9990 15555
rect 15669 15521 15703 15555
rect 18429 15521 18463 15555
rect 8585 15453 8619 15487
rect 13921 15453 13955 15487
rect 14013 15453 14047 15487
rect 15945 15453 15979 15487
rect 17509 15453 17543 15487
rect 3157 15385 3191 15419
rect 6837 15385 6871 15419
rect 15117 15385 15151 15419
rect 1593 15317 1627 15351
rect 2329 15317 2363 15351
rect 2697 15317 2731 15351
rect 3433 15317 3467 15351
rect 3801 15317 3835 15351
rect 7757 15317 7791 15351
rect 8033 15317 8067 15351
rect 9505 15317 9539 15351
rect 11069 15317 11103 15351
rect 12633 15317 12667 15351
rect 13461 15317 13495 15351
rect 15393 15317 15427 15351
rect 18613 15317 18647 15351
rect 2053 15113 2087 15147
rect 2605 15113 2639 15147
rect 3893 15113 3927 15147
rect 5457 15113 5491 15147
rect 5917 15113 5951 15147
rect 7941 15113 7975 15147
rect 8309 15113 8343 15147
rect 8769 15113 8803 15147
rect 10333 15113 10367 15147
rect 12633 15113 12667 15147
rect 13645 15113 13679 15147
rect 14013 15113 14047 15147
rect 16589 15113 16623 15147
rect 17233 15113 17267 15147
rect 17509 15113 17543 15147
rect 18245 15113 18279 15147
rect 18613 15113 18647 15147
rect 2973 15045 3007 15079
rect 4537 15045 4571 15079
rect 6929 15045 6963 15079
rect 9321 15045 9355 15079
rect 10885 15045 10919 15079
rect 12265 15045 12299 15079
rect 4261 14977 4295 15011
rect 4905 14977 4939 15011
rect 7389 14977 7423 15011
rect 9873 14977 9907 15011
rect 1409 14909 1443 14943
rect 3249 14909 3283 14943
rect 3525 14909 3559 14943
rect 15209 14909 15243 14943
rect 3433 14841 3467 14875
rect 5089 14841 5123 14875
rect 6193 14841 6227 14875
rect 7481 14841 7515 14875
rect 9597 14841 9631 14875
rect 10701 14841 10735 14875
rect 11161 14841 11195 14875
rect 11437 14841 11471 14875
rect 11897 14841 11931 14875
rect 12909 14841 12943 14875
rect 13093 14841 13127 14875
rect 13185 14841 13219 14875
rect 14749 14841 14783 14875
rect 15476 14841 15510 14875
rect 1593 14773 1627 14807
rect 4997 14773 5031 14807
rect 6653 14773 6687 14807
rect 7389 14773 7423 14807
rect 9045 14773 9079 14807
rect 9781 14773 9815 14807
rect 11345 14773 11379 14807
rect 14381 14773 14415 14807
rect 15117 14773 15151 14807
rect 2973 14569 3007 14603
rect 3525 14569 3559 14603
rect 5457 14569 5491 14603
rect 6193 14569 6227 14603
rect 8401 14569 8435 14603
rect 9781 14569 9815 14603
rect 10241 14569 10275 14603
rect 12817 14569 12851 14603
rect 13185 14569 13219 14603
rect 15117 14569 15151 14603
rect 15945 14569 15979 14603
rect 17509 14569 17543 14603
rect 2789 14501 2823 14535
rect 3065 14501 3099 14535
rect 4322 14501 4356 14535
rect 6469 14501 6503 14535
rect 13829 14501 13863 14535
rect 13921 14501 13955 14535
rect 15577 14501 15611 14535
rect 4077 14433 4111 14467
rect 6745 14433 6779 14467
rect 7277 14433 7311 14467
rect 11060 14433 11094 14467
rect 16396 14433 16430 14467
rect 2513 14297 2547 14331
rect 7021 14365 7055 14399
rect 10793 14365 10827 14399
rect 13829 14365 13863 14399
rect 16129 14365 16163 14399
rect 13369 14297 13403 14331
rect 1685 14229 1719 14263
rect 2053 14229 2087 14263
rect 3893 14229 3927 14263
rect 6745 14229 6779 14263
rect 6837 14229 6871 14263
rect 9321 14229 9355 14263
rect 10701 14229 10735 14263
rect 12173 14229 12207 14263
rect 14657 14229 14691 14263
rect 2605 14025 2639 14059
rect 2973 14025 3007 14059
rect 4537 14025 4571 14059
rect 5457 14025 5491 14059
rect 8769 14025 8803 14059
rect 9965 14025 9999 14059
rect 10609 14025 10643 14059
rect 14381 14025 14415 14059
rect 14749 14025 14783 14059
rect 1685 13957 1719 13991
rect 5825 13957 5859 13991
rect 10885 13957 10919 13991
rect 15025 13957 15059 13991
rect 2145 13889 2179 13923
rect 3157 13889 3191 13923
rect 5181 13889 5215 13923
rect 6561 13889 6595 13923
rect 6837 13889 6871 13923
rect 15393 13889 15427 13923
rect 3413 13821 3447 13855
rect 5641 13821 5675 13855
rect 6193 13821 6227 13855
rect 7093 13821 7127 13855
rect 11161 13821 11195 13855
rect 12265 13821 12299 13855
rect 12449 13821 12483 13855
rect 15577 13821 15611 13855
rect 16497 13821 16531 13855
rect 2237 13753 2271 13787
rect 10333 13753 10367 13787
rect 11437 13753 11471 13787
rect 12694 13753 12728 13787
rect 2145 13685 2179 13719
rect 8217 13685 8251 13719
rect 11345 13685 11379 13719
rect 11805 13685 11839 13719
rect 13829 13685 13863 13719
rect 15485 13685 15519 13719
rect 16129 13685 16163 13719
rect 1685 13481 1719 13515
rect 2329 13481 2363 13515
rect 3525 13481 3559 13515
rect 6745 13481 6779 13515
rect 7481 13481 7515 13515
rect 9229 13481 9263 13515
rect 11621 13481 11655 13515
rect 14657 13481 14691 13515
rect 17049 13481 17083 13515
rect 2927 13413 2961 13447
rect 3065 13413 3099 13447
rect 4445 13413 4479 13447
rect 4629 13413 4663 13447
rect 5457 13413 5491 13447
rect 6469 13413 6503 13447
rect 7297 13413 7331 13447
rect 12878 13413 12912 13447
rect 15025 13413 15059 13447
rect 15936 13413 15970 13447
rect 2789 13345 2823 13379
rect 4721 13345 4755 13379
rect 5641 13345 5675 13379
rect 12633 13345 12667 13379
rect 18521 13345 18555 13379
rect 7573 13277 7607 13311
rect 11529 13277 11563 13311
rect 11713 13277 11747 13311
rect 12449 13277 12483 13311
rect 15669 13277 15703 13311
rect 18797 13277 18831 13311
rect 4169 13209 4203 13243
rect 11161 13209 11195 13243
rect 2513 13141 2547 13175
rect 3893 13141 3927 13175
rect 5089 13141 5123 13175
rect 5825 13141 5859 13175
rect 7021 13141 7055 13175
rect 7941 13141 7975 13175
rect 8401 13141 8435 13175
rect 10333 13141 10367 13175
rect 10793 13141 10827 13175
rect 14013 13141 14047 13175
rect 15485 13141 15519 13175
rect 2053 12937 2087 12971
rect 2605 12937 2639 12971
rect 3893 12937 3927 12971
rect 4169 12937 4203 12971
rect 5089 12937 5123 12971
rect 5549 12937 5583 12971
rect 8217 12937 8251 12971
rect 9229 12937 9263 12971
rect 10793 12937 10827 12971
rect 11897 12937 11931 12971
rect 12909 12937 12943 12971
rect 14105 12937 14139 12971
rect 14749 12937 14783 12971
rect 16129 12937 16163 12971
rect 18521 12937 18555 12971
rect 2421 12869 2455 12903
rect 6929 12869 6963 12903
rect 10241 12869 10275 12903
rect 13185 12869 13219 12903
rect 3157 12801 3191 12835
rect 4629 12801 4663 12835
rect 6285 12801 6319 12835
rect 6653 12801 6687 12835
rect 7389 12801 7423 12835
rect 9781 12801 9815 12835
rect 11345 12801 11379 12835
rect 12265 12801 12299 12835
rect 13553 12801 13587 12835
rect 15117 12801 15151 12835
rect 16405 12801 16439 12835
rect 1409 12733 1443 12767
rect 2881 12733 2915 12767
rect 4721 12733 4755 12767
rect 5641 12733 5675 12767
rect 7849 12733 7883 12767
rect 14565 12733 14599 12767
rect 15301 12733 15335 12767
rect 3617 12665 3651 12699
rect 4629 12665 4663 12699
rect 7389 12665 7423 12699
rect 7481 12665 7515 12699
rect 8585 12665 8619 12699
rect 9505 12665 9539 12699
rect 11069 12665 11103 12699
rect 13645 12665 13679 12699
rect 13737 12665 13771 12699
rect 1593 12597 1627 12631
rect 3065 12597 3099 12631
rect 5825 12597 5859 12631
rect 8953 12597 8987 12631
rect 9689 12597 9723 12631
rect 10517 12597 10551 12631
rect 11253 12597 11287 12631
rect 15209 12597 15243 12631
rect 15761 12597 15795 12631
rect 1869 12393 1903 12427
rect 3433 12393 3467 12427
rect 3893 12393 3927 12427
rect 5365 12393 5399 12427
rect 7757 12393 7791 12427
rect 11161 12393 11195 12427
rect 14197 12393 14231 12427
rect 2789 12325 2823 12359
rect 2973 12325 3007 12359
rect 4813 12325 4847 12359
rect 10241 12325 10275 12359
rect 11805 12325 11839 12359
rect 13369 12325 13403 12359
rect 15853 12325 15887 12359
rect 3065 12257 3099 12291
rect 4905 12257 4939 12291
rect 5825 12257 5859 12291
rect 6092 12257 6126 12291
rect 10057 12257 10091 12291
rect 10701 12257 10735 12291
rect 11621 12257 11655 12291
rect 13185 12257 13219 12291
rect 13921 12257 13955 12291
rect 15945 12257 15979 12291
rect 19533 12257 19567 12291
rect 4721 12189 4755 12223
rect 5733 12189 5767 12223
rect 8401 12189 8435 12223
rect 10333 12189 10367 12223
rect 11897 12189 11931 12223
rect 13461 12189 13495 12223
rect 15853 12189 15887 12223
rect 2237 12121 2271 12155
rect 4353 12121 4387 12155
rect 12909 12121 12943 12155
rect 15393 12121 15427 12155
rect 2513 12053 2547 12087
rect 7205 12053 7239 12087
rect 8125 12053 8159 12087
rect 9137 12053 9171 12087
rect 9781 12053 9815 12087
rect 11345 12053 11379 12087
rect 12541 12053 12575 12087
rect 14749 12053 14783 12087
rect 15117 12053 15151 12087
rect 19717 12053 19751 12087
rect 1961 11849 1995 11883
rect 5273 11849 5307 11883
rect 6193 11849 6227 11883
rect 6561 11849 6595 11883
rect 8217 11849 8251 11883
rect 9137 11849 9171 11883
rect 10977 11849 11011 11883
rect 11713 11849 11747 11883
rect 13461 11849 13495 11883
rect 13829 11849 13863 11883
rect 15301 11849 15335 11883
rect 16773 11849 16807 11883
rect 19533 11849 19567 11883
rect 4813 11781 4847 11815
rect 9413 11781 9447 11815
rect 9689 11781 9723 11815
rect 12541 11781 12575 11815
rect 6837 11713 6871 11747
rect 10241 11713 10275 11747
rect 12173 11713 12207 11747
rect 2421 11645 2455 11679
rect 5825 11645 5859 11679
rect 7104 11645 7138 11679
rect 9965 11645 9999 11679
rect 12817 11645 12851 11679
rect 14013 11645 14047 11679
rect 14933 11645 14967 11679
rect 15393 11645 15427 11679
rect 2666 11577 2700 11611
rect 5549 11577 5583 11611
rect 10149 11577 10183 11611
rect 10701 11577 10735 11611
rect 11161 11577 11195 11611
rect 13001 11577 13035 11611
rect 13093 11577 13127 11611
rect 14289 11577 14323 11611
rect 15638 11577 15672 11611
rect 1409 11509 1443 11543
rect 2329 11509 2363 11543
rect 3801 11509 3835 11543
rect 4353 11509 4387 11543
rect 5733 11509 5767 11543
rect 2145 11305 2179 11339
rect 2789 11305 2823 11339
rect 5549 11305 5583 11339
rect 5807 11305 5841 11339
rect 6285 11305 6319 11339
rect 7849 11305 7883 11339
rect 9413 11305 9447 11339
rect 10701 11305 10735 11339
rect 11069 11305 11103 11339
rect 13553 11305 13587 11339
rect 15117 11305 15151 11339
rect 16681 11305 16715 11339
rect 2605 11237 2639 11271
rect 2881 11237 2915 11271
rect 4721 11237 4755 11271
rect 4813 11237 4847 11271
rect 6377 11237 6411 11271
rect 8585 11237 8619 11271
rect 10057 11237 10091 11271
rect 10241 11237 10275 11271
rect 14749 11237 14783 11271
rect 3893 11169 3927 11203
rect 5181 11169 5215 11203
rect 8401 11169 8435 11203
rect 11509 11169 11543 11203
rect 13737 11169 13771 11203
rect 15557 11169 15591 11203
rect 3341 11101 3375 11135
rect 4721 11101 4755 11135
rect 6193 11101 6227 11135
rect 8677 11101 8711 11135
rect 8861 11101 8895 11135
rect 10333 11101 10367 11135
rect 11253 11101 11287 11135
rect 14013 11101 14047 11135
rect 15301 11101 15335 11135
rect 2329 11033 2363 11067
rect 4261 11033 4295 11067
rect 7021 11033 7055 11067
rect 8125 11033 8159 11067
rect 9781 11033 9815 11067
rect 13277 11033 13311 11067
rect 1685 10965 1719 10999
rect 7389 10965 7423 10999
rect 8861 10965 8895 10999
rect 9137 10965 9171 10999
rect 12633 10965 12667 10999
rect 2513 10761 2547 10795
rect 2881 10761 2915 10795
rect 5457 10761 5491 10795
rect 6193 10761 6227 10795
rect 7113 10761 7147 10795
rect 9965 10761 9999 10795
rect 11069 10761 11103 10795
rect 13921 10761 13955 10795
rect 14565 10761 14599 10795
rect 15117 10761 15151 10795
rect 1593 10693 1627 10727
rect 8125 10693 8159 10727
rect 2053 10625 2087 10659
rect 3065 10625 3099 10659
rect 7665 10625 7699 10659
rect 12449 10625 12483 10659
rect 12541 10625 12575 10659
rect 15669 10625 15703 10659
rect 2145 10557 2179 10591
rect 3332 10557 3366 10591
rect 5549 10557 5583 10591
rect 7389 10557 7423 10591
rect 8585 10557 8619 10591
rect 8841 10557 8875 10591
rect 2053 10489 2087 10523
rect 6469 10489 6503 10523
rect 12797 10557 12831 10591
rect 16589 10557 16623 10591
rect 17325 10557 17359 10591
rect 14933 10489 14967 10523
rect 15393 10489 15427 10523
rect 16865 10489 16899 10523
rect 4445 10421 4479 10455
rect 5089 10421 5123 10455
rect 5733 10421 5767 10455
rect 7573 10421 7607 10455
rect 8401 10421 8435 10455
rect 10609 10421 10643 10455
rect 11161 10421 11195 10455
rect 11713 10421 11747 10455
rect 12265 10421 12299 10455
rect 12449 10421 12483 10455
rect 15577 10421 15611 10455
rect 16129 10421 16163 10455
rect 1685 10217 1719 10251
rect 2237 10217 2271 10251
rect 3433 10217 3467 10251
rect 3801 10217 3835 10251
rect 4629 10217 4663 10251
rect 4997 10217 5031 10251
rect 7573 10217 7607 10251
rect 9045 10217 9079 10251
rect 9505 10217 9539 10251
rect 9873 10217 9907 10251
rect 11529 10217 11563 10251
rect 12623 10217 12657 10251
rect 14657 10217 14691 10251
rect 2973 10149 3007 10183
rect 5733 10149 5767 10183
rect 8585 10149 8619 10183
rect 8861 10149 8895 10183
rect 10701 10149 10735 10183
rect 13093 10149 13127 10183
rect 13185 10149 13219 10183
rect 15669 10149 15703 10183
rect 15853 10149 15887 10183
rect 4077 10081 4111 10115
rect 6561 10081 6595 10115
rect 6745 10081 6779 10115
rect 10517 10081 10551 10115
rect 11161 10081 11195 10115
rect 12909 10081 12943 10115
rect 14105 10081 14139 10115
rect 2881 10013 2915 10047
rect 3065 10013 3099 10047
rect 5733 10013 5767 10047
rect 5825 10013 5859 10047
rect 6929 10013 6963 10047
rect 8585 10013 8619 10047
rect 8677 10013 8711 10047
rect 8861 10013 8895 10047
rect 10793 10013 10827 10047
rect 12449 10013 12483 10047
rect 15945 10013 15979 10047
rect 2513 9945 2547 9979
rect 6285 9945 6319 9979
rect 8125 9945 8159 9979
rect 15393 9945 15427 9979
rect 4261 9877 4295 9911
rect 5273 9877 5307 9911
rect 7941 9877 7975 9911
rect 10241 9877 10275 9911
rect 11897 9877 11931 9911
rect 13921 9877 13955 9911
rect 14289 9877 14323 9911
rect 15117 9877 15151 9911
rect 3617 9673 3651 9707
rect 9045 9673 9079 9707
rect 9689 9673 9723 9707
rect 10701 9673 10735 9707
rect 15761 9673 15795 9707
rect 16865 9673 16899 9707
rect 2513 9605 2547 9639
rect 6469 9605 6503 9639
rect 6561 9605 6595 9639
rect 6929 9605 6963 9639
rect 11805 9605 11839 9639
rect 12909 9605 12943 9639
rect 13369 9605 13403 9639
rect 3065 9537 3099 9571
rect 1593 9469 1627 9503
rect 2881 9469 2915 9503
rect 4261 9469 4295 9503
rect 4528 9469 4562 9503
rect 6285 9469 6319 9503
rect 1869 9401 1903 9435
rect 8125 9537 8159 9571
rect 9413 9537 9447 9571
rect 10149 9537 10183 9571
rect 8401 9469 8435 9503
rect 10241 9469 10275 9503
rect 12265 9469 12299 9503
rect 12725 9469 12759 9503
rect 13829 9469 13863 9503
rect 14085 9469 14119 9503
rect 16313 9469 16347 9503
rect 7205 9401 7239 9435
rect 7481 9401 7515 9435
rect 16129 9401 16163 9435
rect 4169 9333 4203 9367
rect 5641 9333 5675 9367
rect 6469 9333 6503 9367
rect 7389 9333 7423 9367
rect 8585 9333 8619 9367
rect 10149 9333 10183 9367
rect 10977 9333 11011 9367
rect 11161 9333 11195 9367
rect 13645 9333 13679 9367
rect 15209 9333 15243 9367
rect 16497 9333 16531 9367
rect 1685 9129 1719 9163
rect 3801 9129 3835 9163
rect 4353 9129 4387 9163
rect 8953 9129 8987 9163
rect 9505 9129 9539 9163
rect 9873 9129 9907 9163
rect 10701 9129 10735 9163
rect 12449 9129 12483 9163
rect 13001 9129 13035 9163
rect 14657 9129 14691 9163
rect 15945 9129 15979 9163
rect 2973 9061 3007 9095
rect 5181 9061 5215 9095
rect 14197 9061 14231 9095
rect 2329 8993 2363 9027
rect 3065 8993 3099 9027
rect 3525 8993 3559 9027
rect 4997 8993 5031 9027
rect 7021 8993 7055 9027
rect 7288 8993 7322 9027
rect 9689 8993 9723 9027
rect 11336 8993 11370 9027
rect 15025 8993 15059 9027
rect 15301 8993 15335 9027
rect 16405 8993 16439 9027
rect 2881 8925 2915 8959
rect 5273 8925 5307 8959
rect 6009 8925 6043 8959
rect 11069 8925 11103 8959
rect 14197 8925 14231 8959
rect 14289 8925 14323 8959
rect 13553 8857 13587 8891
rect 2513 8789 2547 8823
rect 4721 8789 4755 8823
rect 5641 8789 5675 8823
rect 6469 8789 6503 8823
rect 6929 8789 6963 8823
rect 8401 8789 8435 8823
rect 10333 8789 10367 8823
rect 13737 8789 13771 8823
rect 15485 8789 15519 8823
rect 16589 8789 16623 8823
rect 2513 8585 2547 8619
rect 3709 8585 3743 8619
rect 6653 8585 6687 8619
rect 7849 8585 7883 8619
rect 11069 8585 11103 8619
rect 11437 8585 11471 8619
rect 11805 8585 11839 8619
rect 16221 8585 16255 8619
rect 16589 8585 16623 8619
rect 3525 8517 3559 8551
rect 5641 8517 5675 8551
rect 7941 8517 7975 8551
rect 8401 8517 8435 8551
rect 9965 8517 9999 8551
rect 12541 8517 12575 8551
rect 14105 8517 14139 8551
rect 15669 8517 15703 8551
rect 1685 8449 1719 8483
rect 3341 8449 3375 8483
rect 1409 8381 1443 8415
rect 7297 8449 7331 8483
rect 4169 8381 4203 8415
rect 4261 8381 4295 8415
rect 6285 8381 6319 8415
rect 7021 8381 7055 8415
rect 3065 8313 3099 8347
rect 3525 8313 3559 8347
rect 4528 8313 4562 8347
rect 9321 8449 9355 8483
rect 10333 8449 10367 8483
rect 10517 8449 10551 8483
rect 13093 8449 13127 8483
rect 14289 8449 14323 8483
rect 8677 8381 8711 8415
rect 12265 8381 12299 8415
rect 12817 8381 12851 8415
rect 8217 8313 8251 8347
rect 8861 8313 8895 8347
rect 8953 8313 8987 8347
rect 13645 8313 13679 8347
rect 14556 8313 14590 8347
rect 16773 8313 16807 8347
rect 2779 8245 2813 8279
rect 3249 8245 3283 8279
rect 7941 8245 7975 8279
rect 9781 8245 9815 8279
rect 10425 8245 10459 8279
rect 13001 8245 13035 8279
rect 2329 8041 2363 8075
rect 3433 8041 3467 8075
rect 3893 8041 3927 8075
rect 4353 8041 4387 8075
rect 4721 8041 4755 8075
rect 6285 8041 6319 8075
rect 8585 8041 8619 8075
rect 8953 8041 8987 8075
rect 10425 8041 10459 8075
rect 10885 8041 10919 8075
rect 14197 8041 14231 8075
rect 15301 8041 15335 8075
rect 17693 8041 17727 8075
rect 2973 7973 3007 8007
rect 8033 7973 8067 8007
rect 11437 7973 11471 8007
rect 11621 7973 11655 8007
rect 11713 7973 11747 8007
rect 13093 7973 13127 8007
rect 13737 7973 13771 8007
rect 13829 7973 13863 8007
rect 14657 7973 14691 8007
rect 5161 7905 5195 7939
rect 7849 7905 7883 7939
rect 9689 7905 9723 7939
rect 16313 7905 16347 7939
rect 16580 7905 16614 7939
rect 2973 7837 3007 7871
rect 3065 7837 3099 7871
rect 4905 7837 4939 7871
rect 8125 7837 8159 7871
rect 9965 7837 9999 7871
rect 13645 7837 13679 7871
rect 14933 7837 14967 7871
rect 7573 7769 7607 7803
rect 12541 7769 12575 7803
rect 1777 7701 1811 7735
rect 2513 7701 2547 7735
rect 6929 7701 6963 7735
rect 7297 7701 7331 7735
rect 9321 7701 9355 7735
rect 11161 7701 11195 7735
rect 12081 7701 12115 7735
rect 13277 7701 13311 7735
rect 15853 7701 15887 7735
rect 16129 7701 16163 7735
rect 1777 7497 1811 7531
rect 3157 7497 3191 7531
rect 4813 7497 4847 7531
rect 5089 7497 5123 7531
rect 6101 7497 6135 7531
rect 7849 7497 7883 7531
rect 8309 7497 8343 7531
rect 10241 7497 10275 7531
rect 12081 7497 12115 7531
rect 14013 7497 14047 7531
rect 17601 7497 17635 7531
rect 3341 7429 3375 7463
rect 4537 7429 4571 7463
rect 6929 7429 6963 7463
rect 9229 7429 9263 7463
rect 10793 7429 10827 7463
rect 11805 7429 11839 7463
rect 14933 7429 14967 7463
rect 15577 7429 15611 7463
rect 3801 7361 3835 7395
rect 5549 7361 5583 7395
rect 5641 7361 5675 7395
rect 7481 7361 7515 7395
rect 11253 7361 11287 7395
rect 11345 7361 11379 7395
rect 12633 7361 12667 7395
rect 14565 7361 14599 7395
rect 16037 7361 16071 7395
rect 2329 7293 2363 7327
rect 3893 7293 3927 7327
rect 7205 7293 7239 7327
rect 8677 7293 8711 7327
rect 10609 7293 10643 7327
rect 12449 7293 12483 7327
rect 13645 7293 13679 7327
rect 14289 7293 14323 7327
rect 2053 7225 2087 7259
rect 2237 7225 2271 7259
rect 9505 7225 9539 7259
rect 9781 7225 9815 7259
rect 11253 7225 11287 7259
rect 13461 7225 13495 7259
rect 16037 7225 16071 7259
rect 16129 7225 16163 7259
rect 18061 7225 18095 7259
rect 2789 7157 2823 7191
rect 3801 7157 3835 7191
rect 5549 7157 5583 7191
rect 6561 7157 6595 7191
rect 7389 7157 7423 7191
rect 9045 7157 9079 7191
rect 9689 7157 9723 7191
rect 13645 7157 13679 7191
rect 13737 7157 13771 7191
rect 14473 7157 14507 7191
rect 15393 7157 15427 7191
rect 16497 7157 16531 7191
rect 16957 7157 16991 7191
rect 17233 7157 17267 7191
rect 18521 7157 18555 7191
rect 2329 6953 2363 6987
rect 2973 6953 3007 6987
rect 6101 6953 6135 6987
rect 7389 6953 7423 6987
rect 7941 6953 7975 6987
rect 9229 6953 9263 6987
rect 10425 6953 10459 6987
rect 14657 6953 14691 6987
rect 17785 6953 17819 6987
rect 4333 6885 4367 6919
rect 7205 6885 7239 6919
rect 11621 6885 11655 6919
rect 3065 6817 3099 6851
rect 3525 6817 3559 6851
rect 7481 6817 7515 6851
rect 8401 6817 8435 6851
rect 9689 6817 9723 6851
rect 10977 6817 11011 6851
rect 11437 6817 11471 6851
rect 12173 6817 12207 6851
rect 12889 6817 12923 6851
rect 14933 6817 14967 6851
rect 15301 6817 15335 6851
rect 15945 6817 15979 6851
rect 16672 6817 16706 6851
rect 1409 6749 1443 6783
rect 2973 6749 3007 6783
rect 4077 6749 4111 6783
rect 8309 6749 8343 6783
rect 9965 6749 9999 6783
rect 11713 6749 11747 6783
rect 12633 6749 12667 6783
rect 16405 6749 16439 6783
rect 18889 6749 18923 6783
rect 2513 6681 2547 6715
rect 6377 6681 6411 6715
rect 11161 6681 11195 6715
rect 1961 6613 1995 6647
rect 3893 6613 3927 6647
rect 5457 6613 5491 6647
rect 6929 6613 6963 6647
rect 8585 6613 8619 6647
rect 12449 6613 12483 6647
rect 14013 6613 14047 6647
rect 15485 6613 15519 6647
rect 16313 6613 16347 6647
rect 18337 6613 18371 6647
rect 18705 6613 18739 6647
rect 19349 6613 19383 6647
rect 4629 6409 4663 6443
rect 5181 6409 5215 6443
rect 8309 6409 8343 6443
rect 10517 6409 10551 6443
rect 13829 6409 13863 6443
rect 14381 6409 14415 6443
rect 15393 6409 15427 6443
rect 15761 6409 15795 6443
rect 15945 6409 15979 6443
rect 16865 6409 16899 6443
rect 17785 6409 17819 6443
rect 6929 6341 6963 6375
rect 10977 6341 11011 6375
rect 5733 6273 5767 6307
rect 6653 6273 6687 6307
rect 7481 6273 7515 6307
rect 8401 6273 8435 6307
rect 11253 6273 11287 6307
rect 16405 6273 16439 6307
rect 18061 6273 18095 6307
rect 1409 6205 1443 6239
rect 2513 6205 2547 6239
rect 2605 6205 2639 6239
rect 11069 6205 11103 6239
rect 12449 6205 12483 6239
rect 2145 6137 2179 6171
rect 2872 6137 2906 6171
rect 5457 6137 5491 6171
rect 6285 6137 6319 6171
rect 7205 6137 7239 6171
rect 7389 6137 7423 6171
rect 8646 6137 8680 6171
rect 12173 6137 12207 6171
rect 12694 6137 12728 6171
rect 15025 6137 15059 6171
rect 16497 6137 16531 6171
rect 18306 6137 18340 6171
rect 1593 6069 1627 6103
rect 3985 6069 4019 6103
rect 4997 6069 5031 6103
rect 5641 6069 5675 6103
rect 7849 6069 7883 6103
rect 9781 6069 9815 6103
rect 11897 6069 11931 6103
rect 16405 6069 16439 6103
rect 17417 6069 17451 6103
rect 19441 6069 19475 6103
rect 3525 5865 3559 5899
rect 3893 5865 3927 5899
rect 5089 5865 5123 5899
rect 5549 5865 5583 5899
rect 7297 5865 7331 5899
rect 9505 5865 9539 5899
rect 13277 5865 13311 5899
rect 15761 5865 15795 5899
rect 18981 5865 19015 5899
rect 19625 5865 19659 5899
rect 2973 5797 3007 5831
rect 4629 5797 4663 5831
rect 4721 5797 4755 5831
rect 11244 5797 11278 5831
rect 14013 5797 14047 5831
rect 14105 5797 14139 5831
rect 16221 5797 16255 5831
rect 16405 5797 16439 5831
rect 16497 5797 16531 5831
rect 3065 5729 3099 5763
rect 4445 5729 4479 5763
rect 6184 5729 6218 5763
rect 8401 5729 8435 5763
rect 9689 5729 9723 5763
rect 9965 5729 9999 5763
rect 10977 5729 11011 5763
rect 14841 5729 14875 5763
rect 17141 5729 17175 5763
rect 17509 5729 17543 5763
rect 17868 5729 17902 5763
rect 2973 5661 3007 5695
rect 5917 5661 5951 5695
rect 13921 5661 13955 5695
rect 17601 5661 17635 5695
rect 20361 5661 20395 5695
rect 2329 5593 2363 5627
rect 4169 5593 4203 5627
rect 7849 5593 7883 5627
rect 13553 5593 13587 5627
rect 15945 5593 15979 5627
rect 1961 5525 1995 5559
rect 2513 5525 2547 5559
rect 8309 5525 8343 5559
rect 8585 5525 8619 5559
rect 9045 5525 9079 5559
rect 10425 5525 10459 5559
rect 10885 5525 10919 5559
rect 12357 5525 12391 5559
rect 12909 5525 12943 5559
rect 14473 5525 14507 5559
rect 20085 5525 20119 5559
rect 1869 5321 1903 5355
rect 4077 5321 4111 5355
rect 5733 5321 5767 5355
rect 7021 5321 7055 5355
rect 7941 5321 7975 5355
rect 8493 5321 8527 5355
rect 10057 5321 10091 5355
rect 10977 5321 11011 5355
rect 13001 5321 13035 5355
rect 15945 5321 15979 5355
rect 16313 5321 16347 5355
rect 19073 5321 19107 5355
rect 19441 5321 19475 5355
rect 21005 5321 21039 5355
rect 2513 5253 2547 5287
rect 3525 5253 3559 5287
rect 6561 5253 6595 5287
rect 16497 5253 16531 5287
rect 18153 5253 18187 5287
rect 19717 5253 19751 5287
rect 2881 5185 2915 5219
rect 3065 5185 3099 5219
rect 4537 5185 4571 5219
rect 7389 5185 7423 5219
rect 7573 5185 7607 5219
rect 8677 5185 8711 5219
rect 13553 5185 13587 5219
rect 16957 5185 16991 5219
rect 18613 5185 18647 5219
rect 20269 5185 20303 5219
rect 2329 5117 2363 5151
rect 4629 5117 4663 5151
rect 5549 5117 5583 5151
rect 6285 5117 6319 5151
rect 11161 5117 11195 5151
rect 12081 5117 12115 5151
rect 12449 5117 12483 5151
rect 13820 5117 13854 5151
rect 15577 5117 15611 5151
rect 17049 5117 17083 5151
rect 18705 5117 18739 5151
rect 20729 5117 20763 5151
rect 4537 5049 4571 5083
rect 4997 5049 5031 5083
rect 7481 5049 7515 5083
rect 8922 5049 8956 5083
rect 13369 5049 13403 5083
rect 17785 5049 17819 5083
rect 18613 5049 18647 5083
rect 19993 5049 20027 5083
rect 2973 4981 3007 5015
rect 3893 4981 3927 5015
rect 5457 4981 5491 5015
rect 10701 4981 10735 5015
rect 11345 4981 11379 5015
rect 11713 4981 11747 5015
rect 12633 4981 12667 5015
rect 14933 4981 14967 5015
rect 16957 4981 16991 5015
rect 17417 4981 17451 5015
rect 20177 4981 20211 5015
rect 4629 4777 4663 4811
rect 5917 4777 5951 4811
rect 6285 4777 6319 4811
rect 8769 4777 8803 4811
rect 10241 4777 10275 4811
rect 12081 4777 12115 4811
rect 13645 4777 13679 4811
rect 14105 4777 14139 4811
rect 16129 4777 16163 4811
rect 19073 4777 19107 4811
rect 2973 4709 3007 4743
rect 3893 4709 3927 4743
rect 4721 4709 4755 4743
rect 6828 4709 6862 4743
rect 13001 4709 13035 4743
rect 13737 4709 13771 4743
rect 4445 4641 4479 4675
rect 6561 4641 6595 4675
rect 10057 4641 10091 4675
rect 11437 4641 11471 4675
rect 12173 4641 12207 4675
rect 13461 4641 13495 4675
rect 15117 4641 15151 4675
rect 16221 4641 16255 4675
rect 16589 4641 16623 4675
rect 17408 4641 17442 4675
rect 19625 4641 19659 4675
rect 20913 4641 20947 4675
rect 1409 4573 1443 4607
rect 2237 4573 2271 4607
rect 2881 4573 2915 4607
rect 3065 4573 3099 4607
rect 10333 4573 10367 4607
rect 12081 4573 12115 4607
rect 12541 4573 12575 4607
rect 16129 4573 16163 4607
rect 17141 4573 17175 4607
rect 20269 4573 20303 4607
rect 2513 4505 2547 4539
rect 4169 4505 4203 4539
rect 9781 4505 9815 4539
rect 14473 4505 14507 4539
rect 18521 4505 18555 4539
rect 19809 4505 19843 4539
rect 1869 4437 1903 4471
rect 3525 4437 3559 4471
rect 5089 4437 5123 4471
rect 5457 4437 5491 4471
rect 7941 4437 7975 4471
rect 9137 4437 9171 4471
rect 9413 4437 9447 4471
rect 10793 4437 10827 4471
rect 11621 4437 11655 4471
rect 13185 4437 13219 4471
rect 15669 4437 15703 4471
rect 16957 4437 16991 4471
rect 19441 4437 19475 4471
rect 20545 4437 20579 4471
rect 21097 4437 21131 4471
rect 21465 4437 21499 4471
rect 3157 4233 3191 4267
rect 4629 4233 4663 4267
rect 6285 4233 6319 4267
rect 10149 4233 10183 4267
rect 11713 4233 11747 4267
rect 13277 4233 13311 4267
rect 15761 4233 15795 4267
rect 17325 4233 17359 4267
rect 21097 4233 21131 4267
rect 6561 4165 6595 4199
rect 7941 4165 7975 4199
rect 10701 4165 10735 4199
rect 19625 4165 19659 4199
rect 3525 4097 3559 4131
rect 5089 4097 5123 4131
rect 5733 4097 5767 4131
rect 5825 4097 5859 4131
rect 7573 4097 7607 4131
rect 8125 4097 8159 4131
rect 12081 4097 12115 4131
rect 13645 4097 13679 4131
rect 13829 4097 13863 4131
rect 16773 4097 16807 4131
rect 18797 4097 18831 4131
rect 2421 4029 2455 4063
rect 2697 4029 2731 4063
rect 3985 4029 4019 4063
rect 5255 4029 5289 4063
rect 6837 4029 6871 4063
rect 11253 4029 11287 4063
rect 12449 4029 12483 4063
rect 16387 4029 16421 4063
rect 18061 4029 18095 4063
rect 19165 4029 19199 4063
rect 20177 4029 20211 4063
rect 20729 4029 20763 4063
rect 21281 4029 21315 4063
rect 21833 4029 21867 4063
rect 2127 3961 2161 3995
rect 4261 3961 4295 3995
rect 7113 3961 7147 3995
rect 8392 3961 8426 3995
rect 10977 3961 11011 3995
rect 12725 3961 12759 3995
rect 14096 3961 14130 3995
rect 16957 3961 16991 3995
rect 17693 3961 17727 3995
rect 18337 3961 18371 3995
rect 19993 3961 20027 3995
rect 1961 3893 1995 3927
rect 2605 3893 2639 3927
rect 3699 3893 3733 3927
rect 4169 3893 4203 3927
rect 5733 3893 5767 3927
rect 9505 3893 9539 3927
rect 10425 3893 10459 3927
rect 11161 3893 11195 3927
rect 15209 3893 15243 3927
rect 16221 3893 16255 3927
rect 16865 3893 16899 3927
rect 20361 3893 20395 3927
rect 21465 3893 21499 3927
rect 22385 3893 22419 3927
rect 2145 3689 2179 3723
rect 2973 3689 3007 3723
rect 3893 3689 3927 3723
rect 6469 3689 6503 3723
rect 8953 3689 8987 3723
rect 10241 3689 10275 3723
rect 12173 3689 12207 3723
rect 12725 3689 12759 3723
rect 13829 3689 13863 3723
rect 14933 3689 14967 3723
rect 16405 3689 16439 3723
rect 17969 3689 18003 3723
rect 21465 3689 21499 3723
rect 2789 3621 2823 3655
rect 4445 3621 4479 3655
rect 4629 3621 4663 3655
rect 6285 3621 6319 3655
rect 6561 3621 6595 3655
rect 7205 3621 7239 3655
rect 8033 3621 8067 3655
rect 8125 3621 8159 3655
rect 9505 3621 9539 3655
rect 10609 3621 10643 3655
rect 13185 3621 13219 3655
rect 13645 3621 13679 3655
rect 15577 3621 15611 3655
rect 18889 3621 18923 3655
rect 1409 3553 1443 3587
rect 3065 3553 3099 3587
rect 3525 3553 3559 3587
rect 5641 3553 5675 3587
rect 7849 3553 7883 3587
rect 9689 3553 9723 3587
rect 10793 3553 10827 3587
rect 11060 3553 11094 3587
rect 15301 3553 15335 3587
rect 16845 3553 16879 3587
rect 18521 3553 18555 3587
rect 19073 3553 19107 3587
rect 20913 3553 20947 3587
rect 22017 3553 22051 3587
rect 4721 3485 4755 3519
rect 13921 3485 13955 3519
rect 16589 3485 16623 3519
rect 19625 3485 19659 3519
rect 4169 3417 4203 3451
rect 5273 3417 5307 3451
rect 8493 3417 8527 3451
rect 13369 3417 13403 3451
rect 14381 3417 14415 3451
rect 21097 3417 21131 3451
rect 2513 3349 2547 3383
rect 6009 3349 6043 3383
rect 7573 3349 7607 3383
rect 9873 3349 9907 3383
rect 19257 3349 19291 3383
rect 19993 3349 20027 3383
rect 20361 3349 20395 3383
rect 21833 3349 21867 3383
rect 22201 3349 22235 3383
rect 1777 3145 1811 3179
rect 2145 3145 2179 3179
rect 3249 3145 3283 3179
rect 6009 3145 6043 3179
rect 8493 3145 8527 3179
rect 11529 3145 11563 3179
rect 12173 3145 12207 3179
rect 14473 3145 14507 3179
rect 18153 3145 18187 3179
rect 19073 3145 19107 3179
rect 19441 3145 19475 3179
rect 22017 3145 22051 3179
rect 2329 3077 2363 3111
rect 17417 3077 17451 3111
rect 22661 3077 22695 3111
rect 2881 3009 2915 3043
rect 7113 3009 7147 3043
rect 12449 3009 12483 3043
rect 17877 3009 17911 3043
rect 18521 3009 18555 3043
rect 18705 3009 18739 3043
rect 20085 3009 20119 3043
rect 20269 3009 20303 3043
rect 23673 3009 23707 3043
rect 2605 2941 2639 2975
rect 3801 2941 3835 2975
rect 6561 2941 6595 2975
rect 7380 2941 7414 2975
rect 9045 2941 9079 2975
rect 9505 2941 9539 2975
rect 9597 2941 9631 2975
rect 14749 2941 14783 2975
rect 14933 2941 14967 2975
rect 16865 2941 16899 2975
rect 19699 2941 19733 2975
rect 21189 2941 21223 2975
rect 21465 2941 21499 2975
rect 22477 2941 22511 2975
rect 23029 2941 23063 2975
rect 4046 2873 4080 2907
rect 9842 2873 9876 2907
rect 12694 2873 12728 2907
rect 15178 2873 15212 2907
rect 18613 2873 18647 2907
rect 20177 2873 20211 2907
rect 2789 2805 2823 2839
rect 3709 2805 3743 2839
rect 5181 2805 5215 2839
rect 10977 2805 11011 2839
rect 13829 2805 13863 2839
rect 16313 2805 16347 2839
rect 20913 2805 20947 2839
rect 1961 2601 1995 2635
rect 2973 2601 3007 2635
rect 6745 2601 6779 2635
rect 8309 2601 8343 2635
rect 9505 2601 9539 2635
rect 10333 2601 10367 2635
rect 10885 2601 10919 2635
rect 15209 2601 15243 2635
rect 16865 2601 16899 2635
rect 18889 2601 18923 2635
rect 19717 2601 19751 2635
rect 20821 2601 20855 2635
rect 21465 2601 21499 2635
rect 3065 2533 3099 2567
rect 4344 2533 4378 2567
rect 6561 2533 6595 2567
rect 7174 2533 7208 2567
rect 10149 2533 10183 2567
rect 10425 2533 10459 2567
rect 12449 2533 12483 2567
rect 13001 2533 13035 2567
rect 13185 2533 13219 2567
rect 13277 2533 13311 2567
rect 13645 2533 13679 2567
rect 20545 2533 20579 2567
rect 3893 2465 3927 2499
rect 4077 2465 4111 2499
rect 1409 2397 1443 2431
rect 2329 2397 2363 2431
rect 2973 2397 3007 2431
rect 6929 2465 6963 2499
rect 9229 2465 9263 2499
rect 11161 2465 11195 2499
rect 11345 2465 11379 2499
rect 12081 2465 12115 2499
rect 14197 2465 14231 2499
rect 14749 2465 14783 2499
rect 15485 2465 15519 2499
rect 15741 2465 15775 2499
rect 17693 2465 17727 2499
rect 18981 2465 19015 2499
rect 19901 2465 19935 2499
rect 21281 2465 21315 2499
rect 21833 2465 21867 2499
rect 22477 2465 22511 2499
rect 23029 2465 23063 2499
rect 24041 2465 24075 2499
rect 24593 2465 24627 2499
rect 14105 2397 14139 2431
rect 18797 2397 18831 2431
rect 9873 2329 9907 2363
rect 12725 2329 12759 2363
rect 14381 2329 14415 2363
rect 18429 2329 18463 2363
rect 20085 2329 20119 2363
rect 22661 2329 22695 2363
rect 2513 2261 2547 2295
rect 3525 2261 3559 2295
rect 5457 2261 5491 2295
rect 6285 2261 6319 2295
rect 6561 2261 6595 2295
rect 11529 2261 11563 2295
rect 18061 2261 18095 2295
rect 22201 2261 22235 2295
rect 24225 2261 24259 2295
<< metal1 >>
rect 4062 26256 4068 26308
rect 4120 26296 4126 26308
rect 12158 26296 12164 26308
rect 4120 26268 12164 26296
rect 4120 26256 4126 26268
rect 12158 26256 12164 26268
rect 12216 26256 12222 26308
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 2314 25440 2320 25492
rect 2372 25480 2378 25492
rect 5442 25480 5448 25492
rect 2372 25452 3372 25480
rect 2372 25440 2378 25452
rect 3344 25276 3372 25452
rect 4724 25452 5448 25480
rect 3418 25372 3424 25424
rect 3476 25412 3482 25424
rect 4724 25421 4752 25452
rect 5442 25440 5448 25452
rect 5500 25440 5506 25492
rect 4709 25415 4767 25421
rect 4709 25412 4721 25415
rect 3476 25384 4721 25412
rect 3476 25372 3482 25384
rect 4709 25381 4721 25384
rect 4755 25381 4767 25415
rect 4709 25375 4767 25381
rect 4893 25415 4951 25421
rect 4893 25381 4905 25415
rect 4939 25412 4951 25415
rect 5166 25412 5172 25424
rect 4939 25384 5172 25412
rect 4939 25381 4951 25384
rect 4893 25375 4951 25381
rect 3510 25304 3516 25356
rect 3568 25344 3574 25356
rect 4985 25347 5043 25353
rect 4985 25344 4997 25347
rect 3568 25316 4997 25344
rect 3568 25304 3574 25316
rect 4985 25313 4997 25316
rect 5031 25313 5043 25347
rect 4985 25307 5043 25313
rect 5092 25276 5120 25384
rect 5166 25372 5172 25384
rect 5224 25412 5230 25424
rect 8113 25415 8171 25421
rect 8113 25412 8125 25415
rect 5224 25384 8125 25412
rect 5224 25372 5230 25384
rect 8113 25381 8125 25384
rect 8159 25412 8171 25415
rect 8570 25412 8576 25424
rect 8159 25384 8576 25412
rect 8159 25381 8171 25384
rect 8113 25375 8171 25381
rect 8570 25372 8576 25384
rect 8628 25372 8634 25424
rect 11333 25415 11391 25421
rect 11333 25381 11345 25415
rect 11379 25412 11391 25415
rect 11514 25412 11520 25424
rect 11379 25384 11520 25412
rect 11379 25381 11391 25384
rect 11333 25375 11391 25381
rect 11514 25372 11520 25384
rect 11572 25372 11578 25424
rect 7006 25304 7012 25356
rect 7064 25344 7070 25356
rect 7929 25347 7987 25353
rect 7929 25344 7941 25347
rect 7064 25316 7941 25344
rect 7064 25304 7070 25316
rect 7929 25313 7941 25316
rect 7975 25313 7987 25347
rect 7929 25307 7987 25313
rect 11054 25304 11060 25356
rect 11112 25344 11118 25356
rect 11149 25347 11207 25353
rect 11149 25344 11161 25347
rect 11112 25316 11161 25344
rect 11112 25304 11118 25316
rect 11149 25313 11161 25316
rect 11195 25313 11207 25347
rect 11149 25307 11207 25313
rect 13909 25347 13967 25353
rect 13909 25313 13921 25347
rect 13955 25344 13967 25347
rect 13998 25344 14004 25356
rect 13955 25316 14004 25344
rect 13955 25313 13967 25316
rect 13909 25307 13967 25313
rect 13998 25304 14004 25316
rect 14056 25304 14062 25356
rect 3344 25248 5120 25276
rect 8205 25279 8263 25285
rect 8205 25245 8217 25279
rect 8251 25276 8263 25279
rect 8478 25276 8484 25288
rect 8251 25248 8484 25276
rect 8251 25245 8263 25248
rect 8205 25239 8263 25245
rect 8478 25236 8484 25248
rect 8536 25236 8542 25288
rect 11425 25279 11483 25285
rect 11425 25245 11437 25279
rect 11471 25276 11483 25279
rect 11882 25276 11888 25288
rect 11471 25248 11888 25276
rect 11471 25245 11483 25248
rect 11425 25239 11483 25245
rect 11882 25236 11888 25248
rect 11940 25236 11946 25288
rect 5626 25168 5632 25220
rect 5684 25208 5690 25220
rect 6454 25208 6460 25220
rect 5684 25180 6460 25208
rect 5684 25168 5690 25180
rect 6454 25168 6460 25180
rect 6512 25168 6518 25220
rect 7285 25211 7343 25217
rect 7285 25177 7297 25211
rect 7331 25208 7343 25211
rect 7926 25208 7932 25220
rect 7331 25180 7932 25208
rect 7331 25177 7343 25180
rect 7285 25171 7343 25177
rect 7926 25168 7932 25180
rect 7984 25168 7990 25220
rect 23474 25168 23480 25220
rect 23532 25208 23538 25220
rect 24302 25208 24308 25220
rect 23532 25180 24308 25208
rect 23532 25168 23538 25180
rect 24302 25168 24308 25180
rect 24360 25168 24366 25220
rect 4430 25140 4436 25152
rect 4391 25112 4436 25140
rect 4430 25100 4436 25112
rect 4488 25100 4494 25152
rect 7653 25143 7711 25149
rect 7653 25109 7665 25143
rect 7699 25140 7711 25143
rect 7742 25140 7748 25152
rect 7699 25112 7748 25140
rect 7699 25109 7711 25112
rect 7653 25103 7711 25109
rect 7742 25100 7748 25112
rect 7800 25100 7806 25152
rect 10137 25143 10195 25149
rect 10137 25109 10149 25143
rect 10183 25140 10195 25143
rect 10778 25140 10784 25152
rect 10183 25112 10784 25140
rect 10183 25109 10195 25112
rect 10137 25103 10195 25109
rect 10778 25100 10784 25112
rect 10836 25100 10842 25152
rect 10873 25143 10931 25149
rect 10873 25109 10885 25143
rect 10919 25140 10931 25143
rect 10962 25140 10968 25152
rect 10919 25112 10968 25140
rect 10919 25109 10931 25112
rect 10873 25103 10931 25109
rect 10962 25100 10968 25112
rect 11020 25100 11026 25152
rect 14093 25143 14151 25149
rect 14093 25109 14105 25143
rect 14139 25140 14151 25143
rect 25958 25140 25964 25152
rect 14139 25112 25964 25140
rect 14139 25109 14151 25112
rect 14093 25103 14151 25109
rect 25958 25100 25964 25112
rect 26016 25100 26022 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 2866 24896 2872 24948
rect 2924 24936 2930 24948
rect 3602 24936 3608 24948
rect 2924 24908 3608 24936
rect 2924 24896 2930 24908
rect 3602 24896 3608 24908
rect 3660 24896 3666 24948
rect 5077 24939 5135 24945
rect 5077 24905 5089 24939
rect 5123 24936 5135 24939
rect 5166 24936 5172 24948
rect 5123 24908 5172 24936
rect 5123 24905 5135 24908
rect 5077 24899 5135 24905
rect 5166 24896 5172 24908
rect 5224 24896 5230 24948
rect 11974 24936 11980 24948
rect 5276 24908 11980 24936
rect 2041 24871 2099 24877
rect 2041 24837 2053 24871
rect 2087 24868 2099 24871
rect 3510 24868 3516 24880
rect 2087 24840 3516 24868
rect 2087 24837 2099 24840
rect 2041 24831 2099 24837
rect 3510 24828 3516 24840
rect 3568 24828 3574 24880
rect 4062 24828 4068 24880
rect 4120 24868 4126 24880
rect 5276 24868 5304 24908
rect 11974 24896 11980 24908
rect 12032 24896 12038 24948
rect 4120 24840 5304 24868
rect 4120 24828 4126 24840
rect 8478 24828 8484 24880
rect 8536 24868 8542 24880
rect 8665 24871 8723 24877
rect 8665 24868 8677 24871
rect 8536 24840 8677 24868
rect 8536 24828 8542 24840
rect 8665 24837 8677 24840
rect 8711 24868 8723 24871
rect 11882 24868 11888 24880
rect 8711 24840 11888 24868
rect 8711 24837 8723 24840
rect 8665 24831 8723 24837
rect 11882 24828 11888 24840
rect 11940 24828 11946 24880
rect 1394 24760 1400 24812
rect 1452 24800 1458 24812
rect 1581 24803 1639 24809
rect 1581 24800 1593 24803
rect 1452 24772 1593 24800
rect 1452 24760 1458 24772
rect 1581 24769 1593 24772
rect 1627 24769 1639 24803
rect 1581 24763 1639 24769
rect 4430 24760 4436 24812
rect 4488 24800 4494 24812
rect 4525 24803 4583 24809
rect 4525 24800 4537 24803
rect 4488 24772 4537 24800
rect 4488 24760 4494 24772
rect 4525 24769 4537 24772
rect 4571 24800 4583 24803
rect 5721 24803 5779 24809
rect 5721 24800 5733 24803
rect 4571 24772 5733 24800
rect 4571 24769 4583 24772
rect 4525 24763 4583 24769
rect 5721 24769 5733 24772
rect 5767 24769 5779 24803
rect 5721 24763 5779 24769
rect 6086 24760 6092 24812
rect 6144 24800 6150 24812
rect 7745 24803 7803 24809
rect 7745 24800 7757 24803
rect 6144 24772 7757 24800
rect 6144 24760 6150 24772
rect 7745 24769 7757 24772
rect 7791 24800 7803 24803
rect 8941 24803 8999 24809
rect 8941 24800 8953 24803
rect 7791 24772 8953 24800
rect 7791 24769 7803 24772
rect 7745 24763 7803 24769
rect 8941 24769 8953 24772
rect 8987 24769 8999 24803
rect 8941 24763 8999 24769
rect 9953 24803 10011 24809
rect 9953 24769 9965 24803
rect 9999 24800 10011 24803
rect 10597 24803 10655 24809
rect 10597 24800 10609 24803
rect 9999 24772 10609 24800
rect 9999 24769 10011 24772
rect 9953 24763 10011 24769
rect 10597 24769 10609 24772
rect 10643 24800 10655 24803
rect 10870 24800 10876 24812
rect 10643 24772 10876 24800
rect 10643 24769 10655 24772
rect 10597 24763 10655 24769
rect 10870 24760 10876 24772
rect 10928 24760 10934 24812
rect 3418 24692 3424 24744
rect 3476 24732 3482 24744
rect 3789 24735 3847 24741
rect 3789 24732 3801 24735
rect 3476 24704 3801 24732
rect 3476 24692 3482 24704
rect 3789 24701 3801 24704
rect 3835 24701 3847 24735
rect 3789 24695 3847 24701
rect 6641 24735 6699 24741
rect 6641 24701 6653 24735
rect 6687 24732 6699 24735
rect 7650 24732 7656 24744
rect 6687 24704 7656 24732
rect 6687 24701 6699 24704
rect 6641 24695 6699 24701
rect 7650 24692 7656 24704
rect 7708 24732 7714 24744
rect 7837 24735 7895 24741
rect 7708 24704 7788 24732
rect 7708 24692 7714 24704
rect 3145 24667 3203 24673
rect 3145 24633 3157 24667
rect 3191 24664 3203 24667
rect 4614 24664 4620 24676
rect 3191 24636 4620 24664
rect 3191 24633 3203 24636
rect 3145 24627 3203 24633
rect 4614 24624 4620 24636
rect 4672 24624 4678 24676
rect 7760 24673 7788 24704
rect 7837 24701 7849 24735
rect 7883 24732 7895 24735
rect 7926 24732 7932 24744
rect 7883 24704 7932 24732
rect 7883 24701 7895 24704
rect 7837 24695 7895 24701
rect 7926 24692 7932 24704
rect 7984 24692 7990 24744
rect 12989 24735 13047 24741
rect 12989 24732 13001 24735
rect 12820 24704 13001 24732
rect 5353 24667 5411 24673
rect 5353 24664 5365 24667
rect 4724 24636 5365 24664
rect 4062 24605 4068 24608
rect 4055 24599 4068 24605
rect 4055 24565 4067 24599
rect 4120 24596 4126 24608
rect 4120 24568 4155 24596
rect 4055 24559 4068 24565
rect 4062 24556 4068 24559
rect 4120 24556 4126 24568
rect 4430 24556 4436 24608
rect 4488 24596 4494 24608
rect 4525 24599 4583 24605
rect 4525 24596 4537 24599
rect 4488 24568 4537 24596
rect 4488 24556 4494 24568
rect 4525 24565 4537 24568
rect 4571 24596 4583 24599
rect 4724 24596 4752 24636
rect 5353 24633 5365 24636
rect 5399 24633 5411 24667
rect 5353 24627 5411 24633
rect 7745 24667 7803 24673
rect 7745 24633 7757 24667
rect 7791 24633 7803 24667
rect 7745 24627 7803 24633
rect 9858 24624 9864 24676
rect 9916 24664 9922 24676
rect 10689 24667 10747 24673
rect 10689 24664 10701 24667
rect 9916 24636 10701 24664
rect 9916 24624 9922 24636
rect 10689 24633 10701 24636
rect 10735 24633 10747 24667
rect 10689 24627 10747 24633
rect 7006 24596 7012 24608
rect 4571 24568 4752 24596
rect 6967 24568 7012 24596
rect 4571 24565 4583 24568
rect 4525 24559 4583 24565
rect 7006 24556 7012 24568
rect 7064 24556 7070 24608
rect 7275 24599 7333 24605
rect 7275 24565 7287 24599
rect 7321 24596 7333 24599
rect 7374 24596 7380 24608
rect 7321 24568 7380 24596
rect 7321 24565 7333 24568
rect 7275 24559 7333 24565
rect 7374 24556 7380 24568
rect 7432 24556 7438 24608
rect 8297 24599 8355 24605
rect 8297 24565 8309 24599
rect 8343 24596 8355 24599
rect 8570 24596 8576 24608
rect 8343 24568 8576 24596
rect 8343 24565 8355 24568
rect 8297 24559 8355 24565
rect 8570 24556 8576 24568
rect 8628 24556 8634 24608
rect 9950 24556 9956 24608
rect 10008 24596 10014 24608
rect 10119 24599 10177 24605
rect 10119 24596 10131 24599
rect 10008 24568 10131 24596
rect 10008 24556 10014 24568
rect 10119 24565 10131 24568
rect 10165 24565 10177 24599
rect 10119 24559 10177 24565
rect 10597 24599 10655 24605
rect 10597 24565 10609 24599
rect 10643 24596 10655 24599
rect 10778 24596 10784 24608
rect 10643 24568 10784 24596
rect 10643 24565 10655 24568
rect 10597 24559 10655 24565
rect 10778 24556 10784 24568
rect 10836 24556 10842 24608
rect 11054 24596 11060 24608
rect 11015 24568 11060 24596
rect 11054 24556 11060 24568
rect 11112 24556 11118 24608
rect 11514 24596 11520 24608
rect 11475 24568 11520 24596
rect 11514 24556 11520 24568
rect 11572 24556 11578 24608
rect 11882 24596 11888 24608
rect 11843 24568 11888 24596
rect 11882 24556 11888 24568
rect 11940 24556 11946 24608
rect 12434 24556 12440 24608
rect 12492 24596 12498 24608
rect 12820 24605 12848 24704
rect 12989 24701 13001 24704
rect 13035 24701 13047 24735
rect 12989 24695 13047 24701
rect 13265 24735 13323 24741
rect 13265 24701 13277 24735
rect 13311 24732 13323 24735
rect 14277 24735 14335 24741
rect 14277 24732 14289 24735
rect 13311 24704 14289 24732
rect 13311 24701 13323 24704
rect 13265 24695 13323 24701
rect 14277 24701 14289 24704
rect 14323 24732 14335 24735
rect 14829 24735 14887 24741
rect 14829 24732 14841 24735
rect 14323 24704 14841 24732
rect 14323 24701 14335 24704
rect 14277 24695 14335 24701
rect 14829 24701 14841 24704
rect 14875 24701 14887 24735
rect 14829 24695 14887 24701
rect 15381 24735 15439 24741
rect 15381 24701 15393 24735
rect 15427 24732 15439 24735
rect 15427 24704 16068 24732
rect 15427 24701 15439 24704
rect 15381 24695 15439 24701
rect 12805 24599 12863 24605
rect 12805 24596 12817 24599
rect 12492 24568 12817 24596
rect 12492 24556 12498 24568
rect 12805 24565 12817 24568
rect 12851 24565 12863 24599
rect 13998 24596 14004 24608
rect 13959 24568 14004 24596
rect 12805 24559 12863 24565
rect 13998 24556 14004 24568
rect 14056 24556 14062 24608
rect 14461 24599 14519 24605
rect 14461 24565 14473 24599
rect 14507 24596 14519 24599
rect 15102 24596 15108 24608
rect 14507 24568 15108 24596
rect 14507 24565 14519 24568
rect 14461 24559 14519 24565
rect 15102 24556 15108 24568
rect 15160 24556 15166 24608
rect 15562 24596 15568 24608
rect 15523 24568 15568 24596
rect 15562 24556 15568 24568
rect 15620 24556 15626 24608
rect 16040 24605 16068 24704
rect 16025 24599 16083 24605
rect 16025 24565 16037 24599
rect 16071 24596 16083 24599
rect 16114 24596 16120 24608
rect 16071 24568 16120 24596
rect 16071 24565 16083 24568
rect 16025 24559 16083 24565
rect 16114 24556 16120 24568
rect 16172 24556 16178 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 2869 24395 2927 24401
rect 2869 24361 2881 24395
rect 2915 24392 2927 24395
rect 3050 24392 3056 24404
rect 2915 24364 3056 24392
rect 2915 24361 2927 24364
rect 2869 24355 2927 24361
rect 3050 24352 3056 24364
rect 3108 24392 3114 24404
rect 3510 24392 3516 24404
rect 3108 24364 3516 24392
rect 3108 24352 3114 24364
rect 3510 24352 3516 24364
rect 3568 24352 3574 24404
rect 7926 24352 7932 24404
rect 7984 24392 7990 24404
rect 8573 24395 8631 24401
rect 8573 24392 8585 24395
rect 7984 24364 8585 24392
rect 7984 24352 7990 24364
rect 8573 24361 8585 24364
rect 8619 24392 8631 24395
rect 8662 24392 8668 24404
rect 8619 24364 8668 24392
rect 8619 24361 8631 24364
rect 8573 24355 8631 24361
rect 8662 24352 8668 24364
rect 8720 24392 8726 24404
rect 9858 24392 9864 24404
rect 8720 24364 9864 24392
rect 8720 24352 8726 24364
rect 9858 24352 9864 24364
rect 9916 24392 9922 24404
rect 10045 24395 10103 24401
rect 10045 24392 10057 24395
rect 9916 24364 10057 24392
rect 9916 24352 9922 24364
rect 10045 24361 10057 24364
rect 10091 24361 10103 24395
rect 10045 24355 10103 24361
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 16482 24392 16488 24404
rect 15519 24364 16488 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 16482 24352 16488 24364
rect 16540 24352 16546 24404
rect 16577 24395 16635 24401
rect 16577 24361 16589 24395
rect 16623 24392 16635 24395
rect 17494 24392 17500 24404
rect 16623 24364 17500 24392
rect 16623 24361 16635 24364
rect 16577 24355 16635 24361
rect 17494 24352 17500 24364
rect 17552 24352 17558 24404
rect 17678 24392 17684 24404
rect 17639 24364 17684 24392
rect 17678 24352 17684 24364
rect 17736 24352 17742 24404
rect 19705 24395 19763 24401
rect 19705 24361 19717 24395
rect 19751 24392 19763 24395
rect 19978 24392 19984 24404
rect 19751 24364 19984 24392
rect 19751 24361 19763 24364
rect 19705 24355 19763 24361
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 1670 24284 1676 24336
rect 1728 24333 1734 24336
rect 1728 24327 1792 24333
rect 1728 24293 1746 24327
rect 1780 24293 1792 24327
rect 4890 24324 4896 24336
rect 4851 24296 4896 24324
rect 1728 24287 1792 24293
rect 1728 24284 1734 24287
rect 4890 24284 4896 24296
rect 4948 24284 4954 24336
rect 6362 24284 6368 24336
rect 6420 24324 6426 24336
rect 6549 24327 6607 24333
rect 6549 24324 6561 24327
rect 6420 24296 6561 24324
rect 6420 24284 6426 24296
rect 6549 24293 6561 24296
rect 6595 24293 6607 24327
rect 8110 24324 8116 24336
rect 8071 24296 8116 24324
rect 6549 24287 6607 24293
rect 8110 24284 8116 24296
rect 8168 24284 8174 24336
rect 8205 24327 8263 24333
rect 8205 24293 8217 24327
rect 8251 24324 8263 24327
rect 8478 24324 8484 24336
rect 8251 24296 8484 24324
rect 8251 24293 8263 24296
rect 8205 24287 8263 24293
rect 1489 24259 1547 24265
rect 1489 24225 1501 24259
rect 1535 24256 1547 24259
rect 2498 24256 2504 24268
rect 1535 24228 2504 24256
rect 1535 24225 1547 24228
rect 1489 24219 1547 24225
rect 2498 24216 2504 24228
rect 2556 24216 2562 24268
rect 4614 24216 4620 24268
rect 4672 24256 4678 24268
rect 4985 24259 5043 24265
rect 4985 24256 4997 24259
rect 4672 24228 4997 24256
rect 4672 24216 4678 24228
rect 4985 24225 4997 24228
rect 5031 24225 5043 24259
rect 4985 24219 5043 24225
rect 6641 24259 6699 24265
rect 6641 24225 6653 24259
rect 6687 24256 6699 24259
rect 7101 24259 7159 24265
rect 7101 24256 7113 24259
rect 6687 24228 7113 24256
rect 6687 24225 6699 24228
rect 6641 24219 6699 24225
rect 7101 24225 7113 24228
rect 7147 24256 7159 24259
rect 8220 24256 8248 24287
rect 8478 24284 8484 24296
rect 8536 24284 8542 24336
rect 11048 24327 11106 24333
rect 11048 24293 11060 24327
rect 11094 24324 11106 24327
rect 11146 24324 11152 24336
rect 11094 24296 11152 24324
rect 11094 24293 11106 24296
rect 11048 24287 11106 24293
rect 11146 24284 11152 24296
rect 11204 24284 11210 24336
rect 7147 24228 8248 24256
rect 13909 24259 13967 24265
rect 7147 24225 7159 24228
rect 7101 24219 7159 24225
rect 13909 24225 13921 24259
rect 13955 24225 13967 24259
rect 13909 24219 13967 24225
rect 14185 24259 14243 24265
rect 14185 24225 14197 24259
rect 14231 24256 14243 24259
rect 15286 24256 15292 24268
rect 14231 24228 15292 24256
rect 14231 24225 14243 24228
rect 14185 24219 14243 24225
rect 4893 24191 4951 24197
rect 4893 24157 4905 24191
rect 4939 24157 4951 24191
rect 4893 24151 4951 24157
rect 4908 24120 4936 24151
rect 6270 24148 6276 24200
rect 6328 24188 6334 24200
rect 6457 24191 6515 24197
rect 6457 24188 6469 24191
rect 6328 24160 6469 24188
rect 6328 24148 6334 24160
rect 6457 24157 6469 24160
rect 6503 24157 6515 24191
rect 8021 24191 8079 24197
rect 8021 24188 8033 24191
rect 6457 24151 6515 24157
rect 7392 24160 8033 24188
rect 4982 24120 4988 24132
rect 4908 24092 4988 24120
rect 4982 24080 4988 24092
rect 5040 24080 5046 24132
rect 6086 24120 6092 24132
rect 6047 24092 6092 24120
rect 6086 24080 6092 24092
rect 6144 24080 6150 24132
rect 6914 24080 6920 24132
rect 6972 24120 6978 24132
rect 7392 24129 7420 24160
rect 8021 24157 8033 24160
rect 8067 24157 8079 24191
rect 8021 24151 8079 24157
rect 8294 24148 8300 24200
rect 8352 24188 8358 24200
rect 10594 24188 10600 24200
rect 8352 24160 10600 24188
rect 8352 24148 8358 24160
rect 10594 24148 10600 24160
rect 10652 24188 10658 24200
rect 10781 24191 10839 24197
rect 10781 24188 10793 24191
rect 10652 24160 10793 24188
rect 10652 24148 10658 24160
rect 10781 24157 10793 24160
rect 10827 24157 10839 24191
rect 13924 24188 13952 24219
rect 15286 24216 15292 24228
rect 15344 24216 15350 24268
rect 16390 24256 16396 24268
rect 16351 24228 16396 24256
rect 16390 24216 16396 24228
rect 16448 24216 16454 24268
rect 17402 24216 17408 24268
rect 17460 24256 17466 24268
rect 17497 24259 17555 24265
rect 17497 24256 17509 24259
rect 17460 24228 17509 24256
rect 17460 24216 17466 24228
rect 17497 24225 17509 24228
rect 17543 24225 17555 24259
rect 17497 24219 17555 24225
rect 19521 24259 19579 24265
rect 19521 24225 19533 24259
rect 19567 24256 19579 24259
rect 20162 24256 20168 24268
rect 19567 24228 20168 24256
rect 19567 24225 19579 24228
rect 19521 24219 19579 24225
rect 20162 24216 20168 24228
rect 20220 24216 20226 24268
rect 14274 24188 14280 24200
rect 13924 24160 14280 24188
rect 10781 24151 10839 24157
rect 14274 24148 14280 24160
rect 14332 24148 14338 24200
rect 7377 24123 7435 24129
rect 7377 24120 7389 24123
rect 6972 24092 7389 24120
rect 6972 24080 6978 24092
rect 7377 24089 7389 24092
rect 7423 24089 7435 24123
rect 7650 24120 7656 24132
rect 7611 24092 7656 24120
rect 7377 24083 7435 24089
rect 7650 24080 7656 24092
rect 7708 24080 7714 24132
rect 4430 24052 4436 24064
rect 4391 24024 4436 24052
rect 4430 24012 4436 24024
rect 4488 24012 4494 24064
rect 5905 24055 5963 24061
rect 5905 24021 5917 24055
rect 5951 24052 5963 24055
rect 5994 24052 6000 24064
rect 5951 24024 6000 24052
rect 5951 24021 5963 24024
rect 5905 24015 5963 24021
rect 5994 24012 6000 24024
rect 6052 24012 6058 24064
rect 12066 24012 12072 24064
rect 12124 24052 12130 24064
rect 12161 24055 12219 24061
rect 12161 24052 12173 24055
rect 12124 24024 12173 24052
rect 12124 24012 12130 24024
rect 12161 24021 12173 24024
rect 12207 24021 12219 24055
rect 12161 24015 12219 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1486 23848 1492 23860
rect 1447 23820 1492 23848
rect 1486 23808 1492 23820
rect 1544 23808 1550 23860
rect 4341 23851 4399 23857
rect 4341 23817 4353 23851
rect 4387 23848 4399 23851
rect 4614 23848 4620 23860
rect 4387 23820 4620 23848
rect 4387 23817 4399 23820
rect 4341 23811 4399 23817
rect 4614 23808 4620 23820
rect 4672 23808 4678 23860
rect 6086 23808 6092 23860
rect 6144 23848 6150 23860
rect 6270 23848 6276 23860
rect 6144 23820 6276 23848
rect 6144 23808 6150 23820
rect 6270 23808 6276 23820
rect 6328 23848 6334 23860
rect 6457 23851 6515 23857
rect 6457 23848 6469 23851
rect 6328 23820 6469 23848
rect 6328 23808 6334 23820
rect 6457 23817 6469 23820
rect 6503 23817 6515 23851
rect 8294 23848 8300 23860
rect 8255 23820 8300 23848
rect 6457 23811 6515 23817
rect 8294 23808 8300 23820
rect 8352 23808 8358 23860
rect 10594 23808 10600 23860
rect 10652 23848 10658 23860
rect 11333 23851 11391 23857
rect 11333 23848 11345 23851
rect 10652 23820 11345 23848
rect 10652 23808 10658 23820
rect 11333 23817 11345 23820
rect 11379 23848 11391 23851
rect 12161 23851 12219 23857
rect 12161 23848 12173 23851
rect 11379 23820 12173 23848
rect 11379 23817 11391 23820
rect 11333 23811 11391 23817
rect 12161 23817 12173 23820
rect 12207 23817 12219 23851
rect 15286 23848 15292 23860
rect 15247 23820 15292 23848
rect 12161 23811 12219 23817
rect 5902 23740 5908 23792
rect 5960 23780 5966 23792
rect 5997 23783 6055 23789
rect 5997 23780 6009 23783
rect 5960 23752 6009 23780
rect 5960 23740 5966 23752
rect 5997 23749 6009 23752
rect 6043 23780 6055 23783
rect 6362 23780 6368 23792
rect 6043 23752 6368 23780
rect 6043 23749 6055 23752
rect 5997 23743 6055 23749
rect 6362 23740 6368 23752
rect 6420 23740 6426 23792
rect 6914 23780 6920 23792
rect 6875 23752 6920 23780
rect 6914 23740 6920 23752
rect 6972 23740 6978 23792
rect 2038 23712 2044 23724
rect 1951 23684 2044 23712
rect 2038 23672 2044 23684
rect 2096 23712 2102 23724
rect 2096 23684 3096 23712
rect 2096 23672 2102 23684
rect 3068 23656 3096 23684
rect 7098 23672 7104 23724
rect 7156 23712 7162 23724
rect 8312 23712 8340 23808
rect 8389 23715 8447 23721
rect 8389 23712 8401 23715
rect 7156 23684 8401 23712
rect 7156 23672 7162 23684
rect 8389 23681 8401 23684
rect 8435 23681 8447 23715
rect 10870 23712 10876 23724
rect 10831 23684 10876 23712
rect 8389 23675 8447 23681
rect 10870 23672 10876 23684
rect 10928 23672 10934 23724
rect 12176 23712 12204 23811
rect 15286 23808 15292 23820
rect 15344 23808 15350 23860
rect 16390 23848 16396 23860
rect 16351 23820 16396 23848
rect 16390 23808 16396 23820
rect 16448 23808 16454 23860
rect 17037 23851 17095 23857
rect 17037 23817 17049 23851
rect 17083 23848 17095 23851
rect 17126 23848 17132 23860
rect 17083 23820 17132 23848
rect 17083 23817 17095 23820
rect 17037 23811 17095 23817
rect 17126 23808 17132 23820
rect 17184 23808 17190 23860
rect 17402 23808 17408 23860
rect 17460 23848 17466 23860
rect 17773 23851 17831 23857
rect 17773 23848 17785 23851
rect 17460 23820 17785 23848
rect 17460 23808 17466 23820
rect 17773 23817 17785 23820
rect 17819 23817 17831 23851
rect 18690 23848 18696 23860
rect 18651 23820 18696 23848
rect 17773 23811 17831 23817
rect 18690 23808 18696 23820
rect 18748 23808 18754 23860
rect 19797 23851 19855 23857
rect 19797 23817 19809 23851
rect 19843 23848 19855 23851
rect 20990 23848 20996 23860
rect 19843 23820 20996 23848
rect 19843 23817 19855 23820
rect 19797 23811 19855 23817
rect 20990 23808 20996 23820
rect 21048 23808 21054 23860
rect 22002 23848 22008 23860
rect 21963 23820 22008 23848
rect 22002 23808 22008 23820
rect 22060 23808 22066 23860
rect 12434 23712 12440 23724
rect 12176 23684 12440 23712
rect 12434 23672 12440 23684
rect 12492 23672 12498 23724
rect 15841 23715 15899 23721
rect 15841 23681 15853 23715
rect 15887 23712 15899 23715
rect 16408 23712 16436 23808
rect 20901 23783 20959 23789
rect 20901 23749 20913 23783
rect 20947 23780 20959 23783
rect 22646 23780 22652 23792
rect 20947 23752 22652 23780
rect 20947 23749 20959 23752
rect 20901 23743 20959 23749
rect 22646 23740 22652 23752
rect 22704 23740 22710 23792
rect 15887 23684 16436 23712
rect 15887 23681 15899 23684
rect 15841 23675 15899 23681
rect 1394 23604 1400 23656
rect 1452 23644 1458 23656
rect 1765 23647 1823 23653
rect 1765 23644 1777 23647
rect 1452 23616 1777 23644
rect 1452 23604 1458 23616
rect 1765 23613 1777 23616
rect 1811 23613 1823 23647
rect 1765 23607 1823 23613
rect 2961 23647 3019 23653
rect 2961 23613 2973 23647
rect 3007 23613 3019 23647
rect 2961 23607 3019 23613
rect 2498 23576 2504 23588
rect 2411 23548 2504 23576
rect 2498 23536 2504 23548
rect 2556 23576 2562 23588
rect 2869 23579 2927 23585
rect 2869 23576 2881 23579
rect 2556 23548 2881 23576
rect 2556 23536 2562 23548
rect 2869 23545 2881 23548
rect 2915 23576 2927 23579
rect 2976 23576 3004 23607
rect 3050 23604 3056 23656
rect 3108 23644 3114 23656
rect 3217 23647 3275 23653
rect 3217 23644 3229 23647
rect 3108 23616 3229 23644
rect 3108 23604 3114 23616
rect 3217 23613 3229 23616
rect 3263 23613 3275 23647
rect 4982 23644 4988 23656
rect 4943 23616 4988 23644
rect 3217 23607 3275 23613
rect 4982 23604 4988 23616
rect 5040 23604 5046 23656
rect 5994 23604 6000 23656
rect 6052 23644 6058 23656
rect 7190 23644 7196 23656
rect 6052 23616 7196 23644
rect 6052 23604 6058 23616
rect 7190 23604 7196 23616
rect 7248 23604 7254 23656
rect 8662 23653 8668 23656
rect 8656 23644 8668 23653
rect 8623 23616 8668 23644
rect 8656 23607 8668 23616
rect 8662 23604 8668 23607
rect 8720 23604 8726 23656
rect 15565 23647 15623 23653
rect 15565 23644 15577 23647
rect 14936 23616 15577 23644
rect 3510 23576 3516 23588
rect 2915 23548 3516 23576
rect 2915 23545 2927 23548
rect 2869 23539 2927 23545
rect 3510 23536 3516 23548
rect 3568 23536 3574 23588
rect 5353 23579 5411 23585
rect 5353 23545 5365 23579
rect 5399 23576 5411 23579
rect 7374 23576 7380 23588
rect 5399 23548 7380 23576
rect 5399 23545 5411 23548
rect 5353 23539 5411 23545
rect 7374 23536 7380 23548
rect 7432 23536 7438 23588
rect 7466 23536 7472 23588
rect 7524 23576 7530 23588
rect 7524 23548 9812 23576
rect 7524 23536 7530 23548
rect 9784 23520 9812 23548
rect 11054 23536 11060 23588
rect 11112 23576 11118 23588
rect 11793 23579 11851 23585
rect 11793 23576 11805 23579
rect 11112 23548 11805 23576
rect 11112 23536 11118 23548
rect 11793 23545 11805 23548
rect 11839 23576 11851 23579
rect 12066 23576 12072 23588
rect 11839 23548 12072 23576
rect 11839 23545 11851 23548
rect 11793 23539 11851 23545
rect 12066 23536 12072 23548
rect 12124 23576 12130 23588
rect 12682 23579 12740 23585
rect 12682 23576 12694 23579
rect 12124 23548 12694 23576
rect 12124 23536 12130 23548
rect 12682 23545 12694 23548
rect 12728 23545 12740 23579
rect 12682 23539 12740 23545
rect 1946 23508 1952 23520
rect 1907 23480 1952 23508
rect 1946 23468 1952 23480
rect 2004 23468 2010 23520
rect 5721 23511 5779 23517
rect 5721 23477 5733 23511
rect 5767 23508 5779 23511
rect 6270 23508 6276 23520
rect 5767 23480 6276 23508
rect 5767 23477 5779 23480
rect 5721 23471 5779 23477
rect 6270 23468 6276 23480
rect 6328 23468 6334 23520
rect 7650 23468 7656 23520
rect 7708 23508 7714 23520
rect 7837 23511 7895 23517
rect 7837 23508 7849 23511
rect 7708 23480 7849 23508
rect 7708 23468 7714 23480
rect 7837 23477 7849 23480
rect 7883 23508 7895 23511
rect 8110 23508 8116 23520
rect 7883 23480 8116 23508
rect 7883 23477 7895 23480
rect 7837 23471 7895 23477
rect 8110 23468 8116 23480
rect 8168 23468 8174 23520
rect 9766 23508 9772 23520
rect 9679 23480 9772 23508
rect 9766 23468 9772 23480
rect 9824 23508 9830 23520
rect 10689 23511 10747 23517
rect 10689 23508 10701 23511
rect 9824 23480 10701 23508
rect 9824 23468 9830 23480
rect 10689 23477 10701 23480
rect 10735 23508 10747 23511
rect 11146 23508 11152 23520
rect 10735 23480 11152 23508
rect 10735 23477 10747 23480
rect 10689 23471 10747 23477
rect 11146 23468 11152 23480
rect 11204 23468 11210 23520
rect 13814 23508 13820 23520
rect 13727 23480 13820 23508
rect 13814 23468 13820 23480
rect 13872 23508 13878 23520
rect 14182 23508 14188 23520
rect 13872 23480 14188 23508
rect 13872 23468 13878 23480
rect 14182 23468 14188 23480
rect 14240 23468 14246 23520
rect 14274 23468 14280 23520
rect 14332 23508 14338 23520
rect 14369 23511 14427 23517
rect 14369 23508 14381 23511
rect 14332 23480 14381 23508
rect 14332 23468 14338 23480
rect 14369 23477 14381 23480
rect 14415 23477 14427 23511
rect 14369 23471 14427 23477
rect 14734 23468 14740 23520
rect 14792 23508 14798 23520
rect 14936 23517 14964 23616
rect 15565 23613 15577 23616
rect 15611 23613 15623 23647
rect 16850 23644 16856 23656
rect 16811 23616 16856 23644
rect 15565 23607 15623 23613
rect 16850 23604 16856 23616
rect 16908 23644 16914 23656
rect 17405 23647 17463 23653
rect 17405 23644 17417 23647
rect 16908 23616 17417 23644
rect 16908 23604 16914 23616
rect 17405 23613 17417 23616
rect 17451 23613 17463 23647
rect 18506 23644 18512 23656
rect 18467 23616 18512 23644
rect 17405 23607 17463 23613
rect 18506 23604 18512 23616
rect 18564 23644 18570 23656
rect 19061 23647 19119 23653
rect 19061 23644 19073 23647
rect 18564 23616 19073 23644
rect 18564 23604 18570 23616
rect 19061 23613 19073 23616
rect 19107 23613 19119 23647
rect 19613 23647 19671 23653
rect 19613 23644 19625 23647
rect 19061 23607 19119 23613
rect 19536 23616 19625 23644
rect 19536 23520 19564 23616
rect 19613 23613 19625 23616
rect 19659 23613 19671 23647
rect 20714 23644 20720 23656
rect 20675 23616 20720 23644
rect 19613 23607 19671 23613
rect 20714 23604 20720 23616
rect 20772 23644 20778 23656
rect 21269 23647 21327 23653
rect 21269 23644 21281 23647
rect 20772 23616 21281 23644
rect 20772 23604 20778 23616
rect 21269 23613 21281 23616
rect 21315 23613 21327 23647
rect 21818 23644 21824 23656
rect 21731 23616 21824 23644
rect 21269 23607 21327 23613
rect 21818 23604 21824 23616
rect 21876 23644 21882 23656
rect 22373 23647 22431 23653
rect 22373 23644 22385 23647
rect 21876 23616 22385 23644
rect 21876 23604 21882 23616
rect 22373 23613 22385 23616
rect 22419 23613 22431 23647
rect 22373 23607 22431 23613
rect 14921 23511 14979 23517
rect 14921 23508 14933 23511
rect 14792 23480 14933 23508
rect 14792 23468 14798 23480
rect 14921 23477 14933 23480
rect 14967 23477 14979 23511
rect 19518 23508 19524 23520
rect 19479 23480 19524 23508
rect 14921 23471 14979 23477
rect 19518 23468 19524 23480
rect 19576 23468 19582 23520
rect 20162 23508 20168 23520
rect 20123 23480 20168 23508
rect 20162 23468 20168 23480
rect 20220 23468 20226 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1670 23304 1676 23316
rect 1631 23276 1676 23304
rect 1670 23264 1676 23276
rect 1728 23264 1734 23316
rect 1946 23304 1952 23316
rect 1907 23276 1952 23304
rect 1946 23264 1952 23276
rect 2004 23264 2010 23316
rect 4430 23264 4436 23316
rect 4488 23304 4494 23316
rect 5077 23307 5135 23313
rect 5077 23304 5089 23307
rect 4488 23276 5089 23304
rect 4488 23264 4494 23276
rect 5077 23273 5089 23276
rect 5123 23304 5135 23307
rect 5166 23304 5172 23316
rect 5123 23276 5172 23304
rect 5123 23273 5135 23276
rect 5077 23267 5135 23273
rect 5166 23264 5172 23276
rect 5224 23264 5230 23316
rect 5534 23264 5540 23316
rect 5592 23304 5598 23316
rect 6089 23307 6147 23313
rect 6089 23304 6101 23307
rect 5592 23276 6101 23304
rect 5592 23264 5598 23276
rect 6089 23273 6101 23276
rect 6135 23273 6147 23307
rect 6089 23267 6147 23273
rect 6917 23307 6975 23313
rect 6917 23273 6929 23307
rect 6963 23304 6975 23307
rect 7466 23304 7472 23316
rect 6963 23276 7472 23304
rect 6963 23273 6975 23276
rect 6917 23267 6975 23273
rect 7466 23264 7472 23276
rect 7524 23264 7530 23316
rect 8481 23307 8539 23313
rect 8481 23273 8493 23307
rect 8527 23304 8539 23307
rect 8662 23304 8668 23316
rect 8527 23276 8668 23304
rect 8527 23273 8539 23276
rect 8481 23267 8539 23273
rect 8662 23264 8668 23276
rect 8720 23264 8726 23316
rect 10042 23264 10048 23316
rect 10100 23304 10106 23316
rect 10321 23307 10379 23313
rect 10321 23304 10333 23307
rect 10100 23276 10333 23304
rect 10100 23264 10106 23276
rect 10321 23273 10333 23276
rect 10367 23304 10379 23307
rect 11057 23307 11115 23313
rect 11057 23304 11069 23307
rect 10367 23276 11069 23304
rect 10367 23273 10379 23276
rect 10321 23267 10379 23273
rect 11057 23273 11069 23276
rect 11103 23273 11115 23307
rect 13814 23304 13820 23316
rect 11057 23267 11115 23273
rect 12728 23276 13820 23304
rect 12728 23248 12756 23276
rect 13814 23264 13820 23276
rect 13872 23264 13878 23316
rect 17037 23307 17095 23313
rect 17037 23273 17049 23307
rect 17083 23304 17095 23307
rect 17862 23304 17868 23316
rect 17083 23276 17868 23304
rect 17083 23273 17095 23276
rect 17037 23267 17095 23273
rect 17862 23264 17868 23276
rect 17920 23264 17926 23316
rect 18141 23307 18199 23313
rect 18141 23273 18153 23307
rect 18187 23304 18199 23307
rect 19242 23304 19248 23316
rect 18187 23276 19248 23304
rect 18187 23273 18199 23276
rect 18141 23267 18199 23273
rect 19242 23264 19248 23276
rect 19300 23264 19306 23316
rect 22002 23304 22008 23316
rect 21963 23276 22008 23304
rect 22002 23264 22008 23276
rect 22060 23264 22066 23316
rect 2961 23239 3019 23245
rect 2961 23205 2973 23239
rect 3007 23205 3019 23239
rect 2961 23199 3019 23205
rect 2866 23128 2872 23180
rect 2924 23168 2930 23180
rect 2976 23168 3004 23199
rect 3050 23196 3056 23248
rect 3108 23236 3114 23248
rect 3421 23239 3479 23245
rect 3421 23236 3433 23239
rect 3108 23208 3433 23236
rect 3108 23196 3114 23208
rect 3421 23205 3433 23208
rect 3467 23205 3479 23239
rect 5902 23236 5908 23248
rect 5863 23208 5908 23236
rect 3421 23199 3479 23205
rect 5902 23196 5908 23208
rect 5960 23196 5966 23248
rect 12066 23196 12072 23248
rect 12124 23236 12130 23248
rect 12621 23239 12679 23245
rect 12621 23236 12633 23239
rect 12124 23208 12633 23236
rect 12124 23196 12130 23208
rect 12621 23205 12633 23208
rect 12667 23205 12679 23239
rect 12621 23199 12679 23205
rect 12710 23196 12716 23248
rect 12768 23236 12774 23248
rect 13173 23239 13231 23245
rect 12768 23208 12861 23236
rect 12768 23196 12774 23208
rect 13173 23205 13185 23239
rect 13219 23236 13231 23239
rect 14185 23239 14243 23245
rect 14185 23236 14197 23239
rect 13219 23208 14197 23236
rect 13219 23205 13231 23208
rect 13173 23199 13231 23205
rect 14185 23205 14197 23208
rect 14231 23205 14243 23239
rect 14185 23199 14243 23205
rect 15841 23239 15899 23245
rect 15841 23205 15853 23239
rect 15887 23236 15899 23239
rect 15930 23236 15936 23248
rect 15887 23208 15936 23236
rect 15887 23205 15899 23208
rect 15841 23199 15899 23205
rect 2924 23140 3004 23168
rect 2924 23128 2930 23140
rect 4246 23128 4252 23180
rect 4304 23168 4310 23180
rect 4433 23171 4491 23177
rect 4433 23168 4445 23171
rect 4304 23140 4445 23168
rect 4304 23128 4310 23140
rect 4433 23137 4445 23140
rect 4479 23168 4491 23171
rect 4614 23168 4620 23180
rect 4479 23140 4620 23168
rect 4479 23137 4491 23140
rect 4433 23131 4491 23137
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 7098 23168 7104 23180
rect 7059 23140 7104 23168
rect 7098 23128 7104 23140
rect 7156 23128 7162 23180
rect 7374 23177 7380 23180
rect 7368 23168 7380 23177
rect 7287 23140 7380 23168
rect 7368 23131 7380 23140
rect 7432 23168 7438 23180
rect 8110 23168 8116 23180
rect 7432 23140 8116 23168
rect 7374 23128 7380 23131
rect 7432 23128 7438 23140
rect 8110 23128 8116 23140
rect 8168 23128 8174 23180
rect 10042 23168 10048 23180
rect 9955 23140 10048 23168
rect 10042 23128 10048 23140
rect 10100 23168 10106 23180
rect 10873 23171 10931 23177
rect 10873 23168 10885 23171
rect 10100 23140 10885 23168
rect 10100 23128 10106 23140
rect 10873 23137 10885 23140
rect 10919 23137 10931 23171
rect 10873 23131 10931 23137
rect 11790 23128 11796 23180
rect 11848 23168 11854 23180
rect 12437 23171 12495 23177
rect 12437 23168 12449 23171
rect 11848 23140 12449 23168
rect 11848 23128 11854 23140
rect 12437 23137 12449 23140
rect 12483 23137 12495 23171
rect 12437 23131 12495 23137
rect 2958 23100 2964 23112
rect 2919 23072 2964 23100
rect 2958 23060 2964 23072
rect 3016 23060 3022 23112
rect 6181 23103 6239 23109
rect 6181 23069 6193 23103
rect 6227 23100 6239 23103
rect 6270 23100 6276 23112
rect 6227 23072 6276 23100
rect 6227 23069 6239 23072
rect 6181 23063 6239 23069
rect 6270 23060 6276 23072
rect 6328 23060 6334 23112
rect 11054 23060 11060 23112
rect 11112 23100 11118 23112
rect 11149 23103 11207 23109
rect 11149 23100 11161 23103
rect 11112 23072 11161 23100
rect 11112 23060 11118 23072
rect 11149 23069 11161 23072
rect 11195 23069 11207 23103
rect 11149 23063 11207 23069
rect 2501 23035 2559 23041
rect 2501 23001 2513 23035
rect 2547 23032 2559 23035
rect 4709 23035 4767 23041
rect 4709 23032 4721 23035
rect 2547 23004 4721 23032
rect 2547 23001 2559 23004
rect 2501 22995 2559 23001
rect 4709 23001 4721 23004
rect 4755 23032 4767 23035
rect 4890 23032 4896 23044
rect 4755 23004 4896 23032
rect 4755 23001 4767 23004
rect 4709 22995 4767 23001
rect 4890 22992 4896 23004
rect 4948 22992 4954 23044
rect 10594 23032 10600 23044
rect 10555 23004 10600 23032
rect 10594 22992 10600 23004
rect 10652 22992 10658 23044
rect 12161 23035 12219 23041
rect 12161 23001 12173 23035
rect 12207 23032 12219 23035
rect 13188 23032 13216 23199
rect 15930 23196 15936 23208
rect 15988 23196 15994 23248
rect 13541 23171 13599 23177
rect 13541 23137 13553 23171
rect 13587 23168 13599 23171
rect 14277 23171 14335 23177
rect 14277 23168 14289 23171
rect 13587 23140 14289 23168
rect 13587 23137 13599 23140
rect 13541 23131 13599 23137
rect 14277 23137 14289 23140
rect 14323 23168 14335 23171
rect 14642 23168 14648 23180
rect 14323 23140 14648 23168
rect 14323 23137 14335 23140
rect 14277 23131 14335 23137
rect 14642 23128 14648 23140
rect 14700 23168 14706 23180
rect 14700 23140 15976 23168
rect 14700 23128 14706 23140
rect 14185 23103 14243 23109
rect 14185 23069 14197 23103
rect 14231 23100 14243 23103
rect 14458 23100 14464 23112
rect 14231 23072 14464 23100
rect 14231 23069 14243 23072
rect 14185 23063 14243 23069
rect 14458 23060 14464 23072
rect 14516 23060 14522 23112
rect 15838 23100 15844 23112
rect 15799 23072 15844 23100
rect 15838 23060 15844 23072
rect 15896 23060 15902 23112
rect 15948 23109 15976 23140
rect 16758 23128 16764 23180
rect 16816 23168 16822 23180
rect 16853 23171 16911 23177
rect 16853 23168 16865 23171
rect 16816 23140 16865 23168
rect 16816 23128 16822 23140
rect 16853 23137 16865 23140
rect 16899 23137 16911 23171
rect 17954 23168 17960 23180
rect 17915 23140 17960 23168
rect 16853 23131 16911 23137
rect 17954 23128 17960 23140
rect 18012 23128 18018 23180
rect 21726 23128 21732 23180
rect 21784 23168 21790 23180
rect 21821 23171 21879 23177
rect 21821 23168 21833 23171
rect 21784 23140 21833 23168
rect 21784 23128 21790 23140
rect 21821 23137 21833 23140
rect 21867 23137 21879 23171
rect 21821 23131 21879 23137
rect 15933 23103 15991 23109
rect 15933 23069 15945 23103
rect 15979 23069 15991 23103
rect 15933 23063 15991 23069
rect 12207 23004 13216 23032
rect 12207 23001 12219 23004
rect 12161 22995 12219 23001
rect 5629 22967 5687 22973
rect 5629 22933 5641 22967
rect 5675 22964 5687 22967
rect 6730 22964 6736 22976
rect 5675 22936 6736 22964
rect 5675 22933 5687 22936
rect 5629 22927 5687 22933
rect 6730 22924 6736 22936
rect 6788 22924 6794 22976
rect 13722 22964 13728 22976
rect 13683 22936 13728 22964
rect 13722 22924 13728 22936
rect 13780 22924 13786 22976
rect 15378 22964 15384 22976
rect 15339 22936 15384 22964
rect 15378 22924 15384 22936
rect 15436 22924 15442 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2225 22763 2283 22769
rect 2225 22729 2237 22763
rect 2271 22760 2283 22763
rect 2958 22760 2964 22772
rect 2271 22732 2964 22760
rect 2271 22729 2283 22732
rect 2225 22723 2283 22729
rect 2958 22720 2964 22732
rect 3016 22760 3022 22772
rect 3970 22760 3976 22772
rect 3016 22732 3976 22760
rect 3016 22720 3022 22732
rect 3970 22720 3976 22732
rect 4028 22720 4034 22772
rect 4154 22720 4160 22772
rect 4212 22760 4218 22772
rect 4249 22763 4307 22769
rect 4249 22760 4261 22763
rect 4212 22732 4261 22760
rect 4212 22720 4218 22732
rect 4249 22729 4261 22732
rect 4295 22729 4307 22763
rect 4249 22723 4307 22729
rect 5534 22720 5540 22772
rect 5592 22760 5598 22772
rect 5813 22763 5871 22769
rect 5813 22760 5825 22763
rect 5592 22732 5825 22760
rect 5592 22720 5598 22732
rect 5813 22729 5825 22732
rect 5859 22729 5871 22763
rect 5813 22723 5871 22729
rect 5994 22720 6000 22772
rect 6052 22760 6058 22772
rect 6181 22763 6239 22769
rect 6181 22760 6193 22763
rect 6052 22732 6193 22760
rect 6052 22720 6058 22732
rect 6181 22729 6193 22732
rect 6227 22760 6239 22763
rect 6914 22760 6920 22772
rect 6227 22732 6920 22760
rect 6227 22729 6239 22732
rect 6181 22723 6239 22729
rect 6914 22720 6920 22732
rect 6972 22720 6978 22772
rect 7098 22760 7104 22772
rect 7059 22732 7104 22760
rect 7098 22720 7104 22732
rect 7156 22720 7162 22772
rect 7190 22720 7196 22772
rect 7248 22760 7254 22772
rect 7285 22763 7343 22769
rect 7285 22760 7297 22763
rect 7248 22732 7297 22760
rect 7248 22720 7254 22732
rect 7285 22729 7297 22732
rect 7331 22729 7343 22763
rect 8297 22763 8355 22769
rect 8297 22760 8309 22763
rect 7285 22723 7343 22729
rect 7852 22732 8309 22760
rect 4890 22692 4896 22704
rect 4851 22664 4896 22692
rect 4890 22652 4896 22664
rect 4948 22652 4954 22704
rect 6270 22652 6276 22704
rect 6328 22692 6334 22704
rect 6641 22695 6699 22701
rect 6641 22692 6653 22695
rect 6328 22664 6653 22692
rect 6328 22652 6334 22664
rect 6641 22661 6653 22664
rect 6687 22692 6699 22695
rect 7374 22692 7380 22704
rect 6687 22664 7380 22692
rect 6687 22661 6699 22664
rect 6641 22655 6699 22661
rect 7374 22652 7380 22664
rect 7432 22652 7438 22704
rect 3602 22584 3608 22636
rect 3660 22624 3666 22636
rect 7006 22624 7012 22636
rect 3660 22596 7012 22624
rect 3660 22584 3666 22596
rect 7006 22584 7012 22596
rect 7064 22584 7070 22636
rect 7852 22633 7880 22732
rect 8297 22729 8309 22732
rect 8343 22760 8355 22763
rect 8662 22760 8668 22772
rect 8343 22732 8668 22760
rect 8343 22729 8355 22732
rect 8297 22723 8355 22729
rect 8662 22720 8668 22732
rect 8720 22720 8726 22772
rect 9766 22760 9772 22772
rect 9727 22732 9772 22760
rect 9766 22720 9772 22732
rect 9824 22720 9830 22772
rect 10042 22760 10048 22772
rect 10003 22732 10048 22760
rect 10042 22720 10048 22732
rect 10100 22720 10106 22772
rect 11054 22760 11060 22772
rect 11015 22732 11060 22760
rect 11054 22720 11060 22732
rect 11112 22720 11118 22772
rect 11425 22763 11483 22769
rect 11425 22729 11437 22763
rect 11471 22760 11483 22763
rect 12710 22760 12716 22772
rect 11471 22732 12716 22760
rect 11471 22729 11483 22732
rect 11425 22723 11483 22729
rect 12710 22720 12716 22732
rect 12768 22720 12774 22772
rect 13265 22763 13323 22769
rect 13265 22729 13277 22763
rect 13311 22760 13323 22763
rect 14458 22760 14464 22772
rect 13311 22732 14464 22760
rect 13311 22729 13323 22732
rect 13265 22723 13323 22729
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 14642 22720 14648 22772
rect 14700 22760 14706 22772
rect 15105 22763 15163 22769
rect 15105 22760 15117 22763
rect 14700 22732 15117 22760
rect 14700 22720 14706 22732
rect 7837 22627 7895 22633
rect 7837 22593 7849 22627
rect 7883 22593 7895 22627
rect 9784 22624 9812 22720
rect 15028 22704 15056 22732
rect 15105 22729 15117 22732
rect 15151 22729 15163 22763
rect 15105 22723 15163 22729
rect 16022 22720 16028 22772
rect 16080 22760 16086 22772
rect 16393 22763 16451 22769
rect 16393 22760 16405 22763
rect 16080 22732 16405 22760
rect 16080 22720 16086 22732
rect 16393 22729 16405 22732
rect 16439 22729 16451 22763
rect 16393 22723 16451 22729
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 18233 22763 18291 22769
rect 18233 22760 18245 22763
rect 18012 22732 18245 22760
rect 18012 22720 18018 22732
rect 18233 22729 18245 22732
rect 18279 22729 18291 22763
rect 18233 22723 18291 22729
rect 21726 22720 21732 22772
rect 21784 22760 21790 22772
rect 21821 22763 21879 22769
rect 21821 22760 21833 22763
rect 21784 22732 21833 22760
rect 21784 22720 21790 22732
rect 21821 22729 21833 22732
rect 21867 22729 21879 22763
rect 21821 22723 21879 22729
rect 11790 22692 11796 22704
rect 11751 22664 11796 22692
rect 11790 22652 11796 22664
rect 11848 22652 11854 22704
rect 12066 22692 12072 22704
rect 12027 22664 12072 22692
rect 12066 22652 12072 22664
rect 12124 22652 12130 22704
rect 12434 22652 12440 22704
rect 12492 22692 12498 22704
rect 13541 22695 13599 22701
rect 13541 22692 13553 22695
rect 12492 22664 13553 22692
rect 12492 22652 12498 22664
rect 13541 22661 13553 22664
rect 13587 22692 13599 22695
rect 13587 22664 13768 22692
rect 13587 22661 13599 22664
rect 13541 22655 13599 22661
rect 13740 22633 13768 22664
rect 15010 22652 15016 22704
rect 15068 22652 15074 22704
rect 10597 22627 10655 22633
rect 10597 22624 10609 22627
rect 9784 22596 10609 22624
rect 7837 22587 7895 22593
rect 10597 22593 10609 22596
rect 10643 22593 10655 22627
rect 10597 22587 10655 22593
rect 13725 22627 13783 22633
rect 13725 22593 13737 22627
rect 13771 22593 13783 22627
rect 13725 22587 13783 22593
rect 1857 22559 1915 22565
rect 1857 22525 1869 22559
rect 1903 22556 1915 22559
rect 2317 22559 2375 22565
rect 2317 22556 2329 22559
rect 1903 22528 2329 22556
rect 1903 22525 1915 22528
rect 1857 22519 1915 22525
rect 2317 22525 2329 22528
rect 2363 22556 2375 22559
rect 3510 22556 3516 22568
rect 2363 22528 3516 22556
rect 2363 22525 2375 22528
rect 2317 22519 2375 22525
rect 3510 22516 3516 22528
rect 3568 22516 3574 22568
rect 5166 22556 5172 22568
rect 5127 22528 5172 22556
rect 5166 22516 5172 22528
rect 5224 22516 5230 22568
rect 6730 22516 6736 22568
rect 6788 22556 6794 22568
rect 7561 22559 7619 22565
rect 7561 22556 7573 22559
rect 6788 22528 7573 22556
rect 6788 22516 6794 22528
rect 7561 22525 7573 22528
rect 7607 22556 7619 22559
rect 8573 22559 8631 22565
rect 8573 22556 8585 22559
rect 7607 22528 8585 22556
rect 7607 22525 7619 22528
rect 7561 22519 7619 22525
rect 8573 22525 8585 22528
rect 8619 22525 8631 22559
rect 8573 22519 8631 22525
rect 9950 22516 9956 22568
rect 10008 22556 10014 22568
rect 10321 22559 10379 22565
rect 10321 22556 10333 22559
rect 10008 22528 10333 22556
rect 10008 22516 10014 22528
rect 10321 22525 10333 22528
rect 10367 22525 10379 22559
rect 10321 22519 10379 22525
rect 12437 22559 12495 22565
rect 12437 22525 12449 22559
rect 12483 22556 12495 22559
rect 12618 22556 12624 22568
rect 12483 22528 12624 22556
rect 12483 22525 12495 22528
rect 12437 22519 12495 22525
rect 12618 22516 12624 22528
rect 12676 22516 12682 22568
rect 16209 22559 16267 22565
rect 16209 22556 16221 22559
rect 13832 22528 16221 22556
rect 2584 22491 2642 22497
rect 2584 22457 2596 22491
rect 2630 22488 2642 22491
rect 2682 22488 2688 22500
rect 2630 22460 2688 22488
rect 2630 22457 2642 22460
rect 2584 22451 2642 22457
rect 2682 22448 2688 22460
rect 2740 22448 2746 22500
rect 3786 22488 3792 22500
rect 3699 22460 3792 22488
rect 3712 22429 3740 22460
rect 3786 22448 3792 22460
rect 3844 22488 3850 22500
rect 4709 22491 4767 22497
rect 4709 22488 4721 22491
rect 3844 22460 4721 22488
rect 3844 22448 3850 22460
rect 4709 22457 4721 22460
rect 4755 22488 4767 22491
rect 5445 22491 5503 22497
rect 5445 22488 5457 22491
rect 4755 22460 5457 22488
rect 4755 22457 4767 22460
rect 4709 22451 4767 22457
rect 5445 22457 5457 22460
rect 5491 22457 5503 22491
rect 7742 22488 7748 22500
rect 7703 22460 7748 22488
rect 5445 22451 5503 22457
rect 7742 22448 7748 22460
rect 7800 22448 7806 22500
rect 9493 22491 9551 22497
rect 9493 22457 9505 22491
rect 9539 22488 9551 22491
rect 10505 22491 10563 22497
rect 10505 22488 10517 22491
rect 9539 22460 10517 22488
rect 9539 22457 9551 22460
rect 9493 22451 9551 22457
rect 10505 22457 10517 22460
rect 10551 22457 10563 22491
rect 10505 22451 10563 22457
rect 12713 22491 12771 22497
rect 12713 22457 12725 22491
rect 12759 22488 12771 22491
rect 13832 22488 13860 22528
rect 16209 22525 16221 22528
rect 16255 22556 16267 22559
rect 16298 22556 16304 22568
rect 16255 22528 16304 22556
rect 16255 22525 16267 22528
rect 16209 22519 16267 22525
rect 16298 22516 16304 22528
rect 16356 22516 16362 22568
rect 12759 22460 13860 22488
rect 13992 22491 14050 22497
rect 12759 22457 12771 22460
rect 12713 22451 12771 22457
rect 13992 22457 14004 22491
rect 14038 22488 14050 22491
rect 14182 22488 14188 22500
rect 14038 22460 14188 22488
rect 14038 22457 14050 22460
rect 13992 22451 14050 22457
rect 3697 22423 3755 22429
rect 3697 22389 3709 22423
rect 3743 22389 3755 22423
rect 3697 22383 3755 22389
rect 4154 22380 4160 22432
rect 4212 22420 4218 22432
rect 5353 22423 5411 22429
rect 5353 22420 5365 22423
rect 4212 22392 5365 22420
rect 4212 22380 4218 22392
rect 5353 22389 5365 22392
rect 5399 22389 5411 22423
rect 10520 22420 10548 22451
rect 14182 22448 14188 22460
rect 14240 22448 14246 22500
rect 15749 22491 15807 22497
rect 15749 22457 15761 22491
rect 15795 22488 15807 22491
rect 15838 22488 15844 22500
rect 15795 22460 15844 22488
rect 15795 22457 15807 22460
rect 15749 22451 15807 22457
rect 15838 22448 15844 22460
rect 15896 22488 15902 22500
rect 15896 22460 16252 22488
rect 15896 22448 15902 22460
rect 16224 22432 16252 22460
rect 10686 22420 10692 22432
rect 10520 22392 10692 22420
rect 5353 22383 5411 22389
rect 10686 22380 10692 22392
rect 10744 22380 10750 22432
rect 16022 22420 16028 22432
rect 15983 22392 16028 22420
rect 16022 22380 16028 22392
rect 16080 22380 16086 22432
rect 16206 22380 16212 22432
rect 16264 22380 16270 22432
rect 16758 22380 16764 22432
rect 16816 22420 16822 22432
rect 16853 22423 16911 22429
rect 16853 22420 16865 22423
rect 16816 22392 16865 22420
rect 16816 22380 16822 22392
rect 16853 22389 16865 22392
rect 16899 22389 16911 22423
rect 16853 22383 16911 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1949 22219 2007 22225
rect 1949 22185 1961 22219
rect 1995 22216 2007 22219
rect 2038 22216 2044 22228
rect 1995 22188 2044 22216
rect 1995 22185 2007 22188
rect 1949 22179 2007 22185
rect 2038 22176 2044 22188
rect 2096 22176 2102 22228
rect 2961 22219 3019 22225
rect 2961 22185 2973 22219
rect 3007 22216 3019 22219
rect 4249 22219 4307 22225
rect 4249 22216 4261 22219
rect 3007 22188 4261 22216
rect 3007 22185 3019 22188
rect 2961 22179 3019 22185
rect 4249 22185 4261 22188
rect 4295 22216 4307 22219
rect 4890 22216 4896 22228
rect 4295 22188 4896 22216
rect 4295 22185 4307 22188
rect 4249 22179 4307 22185
rect 4890 22176 4896 22188
rect 4948 22176 4954 22228
rect 6822 22216 6828 22228
rect 5644 22188 6828 22216
rect 2866 22148 2872 22160
rect 2792 22120 2872 22148
rect 2317 22083 2375 22089
rect 2317 22049 2329 22083
rect 2363 22080 2375 22083
rect 2792 22080 2820 22120
rect 2866 22108 2872 22120
rect 2924 22108 2930 22160
rect 3142 22108 3148 22160
rect 3200 22148 3206 22160
rect 5534 22148 5540 22160
rect 3200 22120 5540 22148
rect 3200 22108 3206 22120
rect 5534 22108 5540 22120
rect 5592 22148 5598 22160
rect 5644 22157 5672 22188
rect 6822 22176 6828 22188
rect 6880 22176 6886 22228
rect 7742 22176 7748 22228
rect 7800 22216 7806 22228
rect 8021 22219 8079 22225
rect 8021 22216 8033 22219
rect 7800 22188 8033 22216
rect 7800 22176 7806 22188
rect 8021 22185 8033 22188
rect 8067 22185 8079 22219
rect 9950 22216 9956 22228
rect 9911 22188 9956 22216
rect 8021 22179 8079 22185
rect 9950 22176 9956 22188
rect 10008 22176 10014 22228
rect 13725 22219 13783 22225
rect 13725 22185 13737 22219
rect 13771 22216 13783 22219
rect 13814 22216 13820 22228
rect 13771 22188 13820 22216
rect 13771 22185 13783 22188
rect 13725 22179 13783 22185
rect 13814 22176 13820 22188
rect 13872 22176 13878 22228
rect 14182 22216 14188 22228
rect 14143 22188 14188 22216
rect 14182 22176 14188 22188
rect 14240 22176 14246 22228
rect 14274 22176 14280 22228
rect 14332 22216 14338 22228
rect 15010 22216 15016 22228
rect 14332 22188 15016 22216
rect 14332 22176 14338 22188
rect 15010 22176 15016 22188
rect 15068 22176 15074 22228
rect 15838 22216 15844 22228
rect 15799 22188 15844 22216
rect 15838 22176 15844 22188
rect 15896 22176 15902 22228
rect 16298 22216 16304 22228
rect 16259 22188 16304 22216
rect 16298 22176 16304 22188
rect 16356 22176 16362 22228
rect 5629 22151 5687 22157
rect 5629 22148 5641 22151
rect 5592 22120 5641 22148
rect 5592 22108 5598 22120
rect 5629 22117 5641 22120
rect 5675 22117 5687 22151
rect 7193 22151 7251 22157
rect 7193 22148 7205 22151
rect 5629 22111 5687 22117
rect 6564 22120 7205 22148
rect 2363 22052 2820 22080
rect 3329 22083 3387 22089
rect 2363 22049 2375 22052
rect 2317 22043 2375 22049
rect 3329 22049 3341 22083
rect 3375 22080 3387 22083
rect 3513 22083 3571 22089
rect 3513 22080 3525 22083
rect 3375 22052 3525 22080
rect 3375 22049 3387 22052
rect 3329 22043 3387 22049
rect 3513 22049 3525 22052
rect 3559 22080 3571 22083
rect 4062 22080 4068 22092
rect 3559 22052 4068 22080
rect 3559 22049 3571 22052
rect 3513 22043 3571 22049
rect 4062 22040 4068 22052
rect 4120 22040 4126 22092
rect 6564 22080 6592 22120
rect 7193 22117 7205 22120
rect 7239 22148 7251 22151
rect 8202 22148 8208 22160
rect 7239 22120 8208 22148
rect 7239 22117 7251 22120
rect 7193 22111 7251 22117
rect 8202 22108 8208 22120
rect 8260 22108 8266 22160
rect 7006 22080 7012 22092
rect 5184 22052 6592 22080
rect 6967 22052 7012 22080
rect 2958 22012 2964 22024
rect 2919 21984 2964 22012
rect 2958 21972 2964 21984
rect 3016 21972 3022 22024
rect 3050 21972 3056 22024
rect 3108 22012 3114 22024
rect 3108 21984 3153 22012
rect 3108 21972 3114 21984
rect 2498 21944 2504 21956
rect 2459 21916 2504 21944
rect 2498 21904 2504 21916
rect 2556 21904 2562 21956
rect 2590 21904 2596 21956
rect 2648 21944 2654 21956
rect 5184 21953 5212 22052
rect 7006 22040 7012 22052
rect 7064 22040 7070 22092
rect 7745 22083 7803 22089
rect 7745 22049 7757 22083
rect 7791 22080 7803 22083
rect 8110 22080 8116 22092
rect 7791 22052 8116 22080
rect 7791 22049 7803 22052
rect 7745 22043 7803 22049
rect 8110 22040 8116 22052
rect 8168 22040 8174 22092
rect 9858 22040 9864 22092
rect 9916 22080 9922 22092
rect 10502 22080 10508 22092
rect 9916 22052 10508 22080
rect 9916 22040 9922 22052
rect 10502 22040 10508 22052
rect 10560 22040 10566 22092
rect 10778 22040 10784 22092
rect 10836 22080 10842 22092
rect 10945 22083 11003 22089
rect 10945 22080 10957 22083
rect 10836 22052 10957 22080
rect 10836 22040 10842 22052
rect 10945 22049 10957 22052
rect 10991 22049 11003 22083
rect 12618 22080 12624 22092
rect 12579 22052 12624 22080
rect 10945 22043 11003 22049
rect 12618 22040 12624 22052
rect 12676 22040 12682 22092
rect 13446 22040 13452 22092
rect 13504 22080 13510 22092
rect 13541 22083 13599 22089
rect 13541 22080 13553 22083
rect 13504 22052 13553 22080
rect 13504 22040 13510 22052
rect 13541 22049 13553 22052
rect 13587 22049 13599 22083
rect 13541 22043 13599 22049
rect 14458 22040 14464 22092
rect 14516 22080 14522 22092
rect 15378 22080 15384 22092
rect 14516 22052 15384 22080
rect 14516 22040 14522 22052
rect 15378 22040 15384 22052
rect 15436 22080 15442 22092
rect 15657 22083 15715 22089
rect 15657 22080 15669 22083
rect 15436 22052 15669 22080
rect 15436 22040 15442 22052
rect 15657 22049 15669 22052
rect 15703 22049 15715 22083
rect 15657 22043 15715 22049
rect 16206 22040 16212 22092
rect 16264 22080 16270 22092
rect 16853 22083 16911 22089
rect 16853 22080 16865 22083
rect 16264 22052 16865 22080
rect 16264 22040 16270 22052
rect 16853 22049 16865 22052
rect 16899 22080 16911 22083
rect 16942 22080 16948 22092
rect 16899 22052 16948 22080
rect 16899 22049 16911 22052
rect 16853 22043 16911 22049
rect 16942 22040 16948 22052
rect 17000 22040 17006 22092
rect 5626 22012 5632 22024
rect 5587 21984 5632 22012
rect 5626 21972 5632 21984
rect 5684 21972 5690 22024
rect 5721 22015 5779 22021
rect 5721 21981 5733 22015
rect 5767 21981 5779 22015
rect 5721 21975 5779 21981
rect 7285 22015 7343 22021
rect 7285 21981 7297 22015
rect 7331 22012 7343 22015
rect 7374 22012 7380 22024
rect 7331 21984 7380 22012
rect 7331 21981 7343 21984
rect 7285 21975 7343 21981
rect 3789 21947 3847 21953
rect 3789 21944 3801 21947
rect 2648 21916 3801 21944
rect 2648 21904 2654 21916
rect 3789 21913 3801 21916
rect 3835 21913 3847 21947
rect 3789 21907 3847 21913
rect 5169 21947 5227 21953
rect 5169 21913 5181 21947
rect 5215 21913 5227 21947
rect 5169 21907 5227 21913
rect 2682 21836 2688 21888
rect 2740 21876 2746 21888
rect 3329 21879 3387 21885
rect 3329 21876 3341 21879
rect 2740 21848 3341 21876
rect 2740 21836 2746 21848
rect 3329 21845 3341 21848
rect 3375 21845 3387 21879
rect 3329 21839 3387 21845
rect 4985 21879 5043 21885
rect 4985 21845 4997 21879
rect 5031 21876 5043 21879
rect 5736 21876 5764 21975
rect 7374 21972 7380 21984
rect 7432 21972 7438 22024
rect 10594 21972 10600 22024
rect 10652 22012 10658 22024
rect 10689 22015 10747 22021
rect 10689 22012 10701 22015
rect 10652 21984 10701 22012
rect 10652 21972 10658 21984
rect 10689 21981 10701 21984
rect 10735 21981 10747 22015
rect 10689 21975 10747 21981
rect 13817 22015 13875 22021
rect 13817 21981 13829 22015
rect 13863 21981 13875 22015
rect 13817 21975 13875 21981
rect 15933 22015 15991 22021
rect 15933 21981 15945 22015
rect 15979 22012 15991 22015
rect 16022 22012 16028 22024
rect 15979 21984 16028 22012
rect 15979 21981 15991 21984
rect 15933 21975 15991 21981
rect 11882 21904 11888 21956
rect 11940 21944 11946 21956
rect 12069 21947 12127 21953
rect 12069 21944 12081 21947
rect 11940 21916 12081 21944
rect 11940 21904 11946 21916
rect 12069 21913 12081 21916
rect 12115 21944 12127 21947
rect 13078 21944 13084 21956
rect 12115 21916 13084 21944
rect 12115 21913 12127 21916
rect 12069 21907 12127 21913
rect 13078 21904 13084 21916
rect 13136 21944 13142 21956
rect 13832 21944 13860 21975
rect 16022 21972 16028 21984
rect 16080 21972 16086 22024
rect 17034 21944 17040 21956
rect 13136 21916 13860 21944
rect 16995 21916 17040 21944
rect 13136 21904 13142 21916
rect 17034 21904 17040 21916
rect 17092 21904 17098 21956
rect 6270 21876 6276 21888
rect 5031 21848 6276 21876
rect 5031 21845 5043 21848
rect 4985 21839 5043 21845
rect 6270 21836 6276 21848
rect 6328 21836 6334 21888
rect 6730 21876 6736 21888
rect 6691 21848 6736 21876
rect 6730 21836 6736 21848
rect 6788 21836 6794 21888
rect 9030 21876 9036 21888
rect 8991 21848 9036 21876
rect 9030 21836 9036 21848
rect 9088 21836 9094 21888
rect 9398 21876 9404 21888
rect 9359 21848 9404 21876
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 10870 21836 10876 21888
rect 10928 21876 10934 21888
rect 11422 21876 11428 21888
rect 10928 21848 11428 21876
rect 10928 21836 10934 21848
rect 11422 21836 11428 21848
rect 11480 21836 11486 21888
rect 11790 21836 11796 21888
rect 11848 21876 11854 21888
rect 13265 21879 13323 21885
rect 13265 21876 13277 21879
rect 11848 21848 13277 21876
rect 11848 21836 11854 21848
rect 13265 21845 13277 21848
rect 13311 21845 13323 21879
rect 15378 21876 15384 21888
rect 15339 21848 15384 21876
rect 13265 21839 13323 21845
rect 15378 21836 15384 21848
rect 15436 21836 15442 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 5534 21672 5540 21684
rect 5495 21644 5540 21672
rect 5534 21632 5540 21644
rect 5592 21632 5598 21684
rect 6273 21675 6331 21681
rect 6273 21641 6285 21675
rect 6319 21672 6331 21675
rect 7006 21672 7012 21684
rect 6319 21644 7012 21672
rect 6319 21641 6331 21644
rect 6273 21635 6331 21641
rect 7006 21632 7012 21644
rect 7064 21632 7070 21684
rect 8202 21632 8208 21684
rect 8260 21672 8266 21684
rect 8297 21675 8355 21681
rect 8297 21672 8309 21675
rect 8260 21644 8309 21672
rect 8260 21632 8266 21644
rect 8297 21641 8309 21644
rect 8343 21641 8355 21675
rect 9122 21672 9128 21684
rect 9083 21644 9128 21672
rect 8297 21635 8355 21641
rect 9122 21632 9128 21644
rect 9180 21632 9186 21684
rect 10686 21672 10692 21684
rect 10647 21644 10692 21672
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 11882 21672 11888 21684
rect 11843 21644 11888 21672
rect 11882 21632 11888 21644
rect 11940 21632 11946 21684
rect 12526 21672 12532 21684
rect 12487 21644 12532 21672
rect 12526 21632 12532 21644
rect 12584 21632 12590 21684
rect 13354 21632 13360 21684
rect 13412 21672 13418 21684
rect 13814 21672 13820 21684
rect 13412 21644 13820 21672
rect 13412 21632 13418 21644
rect 13814 21632 13820 21644
rect 13872 21632 13878 21684
rect 14458 21672 14464 21684
rect 14419 21644 14464 21672
rect 14458 21632 14464 21644
rect 14516 21632 14522 21684
rect 14734 21632 14740 21684
rect 14792 21672 14798 21684
rect 15013 21675 15071 21681
rect 15013 21672 15025 21675
rect 14792 21644 15025 21672
rect 14792 21632 14798 21644
rect 15013 21641 15025 21644
rect 15059 21641 15071 21675
rect 16942 21672 16948 21684
rect 16903 21644 16948 21672
rect 15013 21635 15071 21641
rect 16942 21632 16948 21644
rect 17000 21632 17006 21684
rect 18322 21672 18328 21684
rect 18283 21644 18328 21672
rect 18322 21632 18328 21644
rect 18380 21632 18386 21684
rect 2041 21607 2099 21613
rect 2041 21573 2053 21607
rect 2087 21604 2099 21607
rect 2958 21604 2964 21616
rect 2087 21576 2964 21604
rect 2087 21573 2099 21576
rect 2041 21567 2099 21573
rect 2958 21564 2964 21576
rect 3016 21564 3022 21616
rect 6917 21607 6975 21613
rect 6917 21573 6929 21607
rect 6963 21604 6975 21607
rect 7742 21604 7748 21616
rect 6963 21576 7748 21604
rect 6963 21573 6975 21576
rect 6917 21567 6975 21573
rect 7742 21564 7748 21576
rect 7800 21564 7806 21616
rect 12434 21564 12440 21616
rect 12492 21604 12498 21616
rect 13446 21604 13452 21616
rect 12492 21576 13452 21604
rect 12492 21564 12498 21576
rect 13446 21564 13452 21576
rect 13504 21564 13510 21616
rect 2498 21536 2504 21548
rect 2459 21508 2504 21536
rect 2498 21496 2504 21508
rect 2556 21496 2562 21548
rect 2608 21508 3648 21536
rect 2608 21477 2636 21508
rect 1857 21471 1915 21477
rect 1857 21437 1869 21471
rect 1903 21468 1915 21471
rect 2593 21471 2651 21477
rect 2593 21468 2605 21471
rect 1903 21440 2605 21468
rect 1903 21437 1915 21440
rect 1857 21431 1915 21437
rect 2593 21437 2605 21440
rect 2639 21437 2651 21471
rect 2593 21431 2651 21437
rect 3421 21471 3479 21477
rect 3421 21437 3433 21471
rect 3467 21468 3479 21471
rect 3510 21468 3516 21480
rect 3467 21440 3516 21468
rect 3467 21437 3479 21440
rect 3421 21431 3479 21437
rect 3510 21428 3516 21440
rect 3568 21428 3574 21480
rect 3620 21468 3648 21508
rect 10502 21496 10508 21548
rect 10560 21536 10566 21548
rect 11241 21539 11299 21545
rect 11241 21536 11253 21539
rect 10560 21508 11253 21536
rect 10560 21496 10566 21508
rect 11241 21505 11253 21508
rect 11287 21505 11299 21539
rect 11241 21499 11299 21505
rect 3786 21477 3792 21480
rect 3780 21468 3792 21477
rect 3620 21440 3792 21468
rect 3780 21431 3792 21440
rect 3786 21428 3792 21431
rect 3844 21428 3850 21480
rect 7374 21428 7380 21480
rect 7432 21468 7438 21480
rect 7469 21471 7527 21477
rect 7469 21468 7481 21471
rect 7432 21440 7481 21468
rect 7432 21428 7438 21440
rect 7469 21437 7481 21440
rect 7515 21468 7527 21471
rect 7837 21471 7895 21477
rect 7837 21468 7849 21471
rect 7515 21440 7849 21468
rect 7515 21437 7527 21440
rect 7469 21431 7527 21437
rect 7837 21437 7849 21440
rect 7883 21437 7895 21471
rect 7837 21431 7895 21437
rect 8941 21471 8999 21477
rect 8941 21437 8953 21471
rect 8987 21468 8999 21471
rect 9677 21471 9735 21477
rect 9677 21468 9689 21471
rect 8987 21440 9689 21468
rect 8987 21437 8999 21440
rect 8941 21431 8999 21437
rect 9677 21437 9689 21440
rect 9723 21468 9735 21471
rect 10042 21468 10048 21480
rect 9723 21440 10048 21468
rect 9723 21437 9735 21440
rect 9677 21431 9735 21437
rect 10042 21428 10048 21440
rect 10100 21428 10106 21480
rect 13078 21468 13084 21480
rect 13039 21440 13084 21468
rect 13078 21428 13084 21440
rect 13136 21428 13142 21480
rect 14734 21428 14740 21480
rect 14792 21468 14798 21480
rect 15289 21471 15347 21477
rect 15289 21468 15301 21471
rect 14792 21440 15301 21468
rect 14792 21428 14798 21440
rect 15289 21437 15301 21440
rect 15335 21468 15347 21471
rect 16301 21471 16359 21477
rect 16301 21468 16313 21471
rect 15335 21440 16313 21468
rect 15335 21437 15347 21440
rect 15289 21431 15347 21437
rect 16301 21437 16313 21440
rect 16347 21437 16359 21471
rect 16301 21431 16359 21437
rect 18141 21471 18199 21477
rect 18141 21437 18153 21471
rect 18187 21468 18199 21471
rect 18322 21468 18328 21480
rect 18187 21440 18328 21468
rect 18187 21437 18199 21440
rect 18141 21431 18199 21437
rect 18322 21428 18328 21440
rect 18380 21468 18386 21480
rect 18693 21471 18751 21477
rect 18693 21468 18705 21471
rect 18380 21440 18705 21468
rect 18380 21428 18386 21440
rect 18693 21437 18705 21440
rect 18739 21437 18751 21471
rect 18693 21431 18751 21437
rect 3050 21400 3056 21412
rect 2963 21372 3056 21400
rect 3050 21360 3056 21372
rect 3108 21400 3114 21412
rect 7193 21403 7251 21409
rect 7193 21400 7205 21403
rect 3108 21372 4936 21400
rect 3108 21360 3114 21372
rect 1578 21292 1584 21344
rect 1636 21332 1642 21344
rect 2501 21335 2559 21341
rect 2501 21332 2513 21335
rect 1636 21304 2513 21332
rect 1636 21292 1642 21304
rect 2501 21301 2513 21304
rect 2547 21332 2559 21335
rect 2590 21332 2596 21344
rect 2547 21304 2596 21332
rect 2547 21301 2559 21304
rect 2501 21295 2559 21301
rect 2590 21292 2596 21304
rect 2648 21292 2654 21344
rect 4908 21341 4936 21372
rect 6840 21372 7205 21400
rect 6840 21344 6868 21372
rect 7193 21369 7205 21372
rect 7239 21369 7251 21403
rect 9398 21400 9404 21412
rect 9359 21372 9404 21400
rect 7193 21363 7251 21369
rect 9398 21360 9404 21372
rect 9456 21360 9462 21412
rect 10965 21403 11023 21409
rect 10965 21369 10977 21403
rect 11011 21400 11023 21403
rect 11238 21400 11244 21412
rect 11011 21372 11244 21400
rect 11011 21369 11023 21372
rect 10965 21363 11023 21369
rect 11238 21360 11244 21372
rect 11296 21400 11302 21412
rect 11790 21400 11796 21412
rect 11296 21372 11796 21400
rect 11296 21360 11302 21372
rect 11790 21360 11796 21372
rect 11848 21360 11854 21412
rect 12526 21360 12532 21412
rect 12584 21400 12590 21412
rect 12805 21403 12863 21409
rect 12805 21400 12817 21403
rect 12584 21372 12817 21400
rect 12584 21360 12590 21372
rect 12805 21369 12817 21372
rect 12851 21369 12863 21403
rect 12805 21363 12863 21369
rect 14829 21403 14887 21409
rect 14829 21369 14841 21403
rect 14875 21400 14887 21403
rect 15565 21403 15623 21409
rect 15565 21400 15577 21403
rect 14875 21372 15577 21400
rect 14875 21369 14887 21372
rect 14829 21363 14887 21369
rect 15565 21369 15577 21372
rect 15611 21400 15623 21403
rect 15654 21400 15660 21412
rect 15611 21372 15660 21400
rect 15611 21369 15623 21372
rect 15565 21363 15623 21369
rect 15654 21360 15660 21372
rect 15712 21360 15718 21412
rect 15746 21360 15752 21412
rect 15804 21400 15810 21412
rect 16485 21403 16543 21409
rect 16485 21400 16497 21403
rect 15804 21372 16497 21400
rect 15804 21360 15810 21372
rect 16485 21369 16497 21372
rect 16531 21369 16543 21403
rect 16485 21363 16543 21369
rect 26234 21360 26240 21412
rect 26292 21400 26298 21412
rect 27614 21400 27620 21412
rect 26292 21372 27620 21400
rect 26292 21360 26298 21372
rect 27614 21360 27620 21372
rect 27672 21360 27678 21412
rect 4893 21335 4951 21341
rect 4893 21301 4905 21335
rect 4939 21332 4951 21335
rect 5258 21332 5264 21344
rect 4939 21304 5264 21332
rect 4939 21301 4951 21304
rect 4893 21295 4951 21301
rect 5258 21292 5264 21304
rect 5316 21292 5322 21344
rect 5905 21335 5963 21341
rect 5905 21301 5917 21335
rect 5951 21332 5963 21335
rect 5994 21332 6000 21344
rect 5951 21304 6000 21332
rect 5951 21301 5963 21304
rect 5905 21295 5963 21301
rect 5994 21292 6000 21304
rect 6052 21292 6058 21344
rect 6641 21335 6699 21341
rect 6641 21301 6653 21335
rect 6687 21332 6699 21335
rect 6822 21332 6828 21344
rect 6687 21304 6828 21332
rect 6687 21301 6699 21304
rect 6641 21295 6699 21301
rect 6822 21292 6828 21304
rect 6880 21292 6886 21344
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 7377 21335 7435 21341
rect 7377 21332 7389 21335
rect 6972 21304 7389 21332
rect 6972 21292 6978 21304
rect 7377 21301 7389 21304
rect 7423 21301 7435 21335
rect 7377 21295 7435 21301
rect 9030 21292 9036 21344
rect 9088 21332 9094 21344
rect 9585 21335 9643 21341
rect 9585 21332 9597 21335
rect 9088 21304 9597 21332
rect 9088 21292 9094 21304
rect 9585 21301 9597 21304
rect 9631 21301 9643 21335
rect 9585 21295 9643 21301
rect 10505 21335 10563 21341
rect 10505 21301 10517 21335
rect 10551 21332 10563 21335
rect 10686 21332 10692 21344
rect 10551 21304 10692 21332
rect 10551 21301 10563 21304
rect 10505 21295 10563 21301
rect 10686 21292 10692 21304
rect 10744 21292 10750 21344
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 11149 21335 11207 21341
rect 11149 21332 11161 21335
rect 11112 21304 11161 21332
rect 11112 21292 11118 21304
rect 11149 21301 11161 21304
rect 11195 21301 11207 21335
rect 11149 21295 11207 21301
rect 11330 21292 11336 21344
rect 11388 21332 11394 21344
rect 12161 21335 12219 21341
rect 12161 21332 12173 21335
rect 11388 21304 12173 21332
rect 11388 21292 11394 21304
rect 12161 21301 12173 21304
rect 12207 21332 12219 21335
rect 12989 21335 13047 21341
rect 12989 21332 13001 21335
rect 12207 21304 13001 21332
rect 12207 21301 12219 21304
rect 12161 21295 12219 21301
rect 12989 21301 13001 21304
rect 13035 21301 13047 21335
rect 12989 21295 13047 21301
rect 15010 21292 15016 21344
rect 15068 21332 15074 21344
rect 15378 21332 15384 21344
rect 15068 21304 15384 21332
rect 15068 21292 15074 21304
rect 15378 21292 15384 21304
rect 15436 21332 15442 21344
rect 15473 21335 15531 21341
rect 15473 21332 15485 21335
rect 15436 21304 15485 21332
rect 15436 21292 15442 21304
rect 15473 21301 15485 21304
rect 15519 21301 15531 21335
rect 16022 21332 16028 21344
rect 15983 21304 16028 21332
rect 15473 21295 15531 21301
rect 16022 21292 16028 21304
rect 16080 21292 16086 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 2314 21088 2320 21140
rect 2372 21128 2378 21140
rect 2409 21131 2467 21137
rect 2409 21128 2421 21131
rect 2372 21100 2421 21128
rect 2372 21088 2378 21100
rect 2409 21097 2421 21100
rect 2455 21097 2467 21131
rect 2409 21091 2467 21097
rect 3605 21131 3663 21137
rect 3605 21097 3617 21131
rect 3651 21128 3663 21131
rect 3786 21128 3792 21140
rect 3651 21100 3792 21128
rect 3651 21097 3663 21100
rect 3605 21091 3663 21097
rect 3786 21088 3792 21100
rect 3844 21088 3850 21140
rect 4246 21128 4252 21140
rect 4207 21100 4252 21128
rect 4246 21088 4252 21100
rect 4304 21088 4310 21140
rect 4709 21131 4767 21137
rect 4709 21097 4721 21131
rect 4755 21128 4767 21131
rect 5442 21128 5448 21140
rect 4755 21100 5448 21128
rect 4755 21097 4767 21100
rect 4709 21091 4767 21097
rect 5442 21088 5448 21100
rect 5500 21088 5506 21140
rect 6270 21128 6276 21140
rect 6231 21100 6276 21128
rect 6270 21088 6276 21100
rect 6328 21088 6334 21140
rect 6914 21128 6920 21140
rect 6875 21100 6920 21128
rect 6914 21088 6920 21100
rect 6972 21088 6978 21140
rect 8389 21131 8447 21137
rect 8389 21128 8401 21131
rect 7760 21100 8401 21128
rect 7760 21072 7788 21100
rect 8389 21097 8401 21100
rect 8435 21097 8447 21131
rect 8389 21091 8447 21097
rect 10042 21088 10048 21140
rect 10100 21128 10106 21140
rect 10778 21128 10784 21140
rect 10100 21100 10784 21128
rect 10100 21088 10106 21100
rect 10778 21088 10784 21100
rect 10836 21128 10842 21140
rect 11057 21131 11115 21137
rect 11057 21128 11069 21131
rect 10836 21100 11069 21128
rect 10836 21088 10842 21100
rect 11057 21097 11069 21100
rect 11103 21097 11115 21131
rect 11057 21091 11115 21097
rect 11974 21088 11980 21140
rect 12032 21128 12038 21140
rect 12526 21128 12532 21140
rect 12032 21100 12532 21128
rect 12032 21088 12038 21100
rect 12526 21088 12532 21100
rect 12584 21088 12590 21140
rect 13078 21088 13084 21140
rect 13136 21128 13142 21140
rect 13173 21131 13231 21137
rect 13173 21128 13185 21131
rect 13136 21100 13185 21128
rect 13136 21088 13142 21100
rect 13173 21097 13185 21100
rect 13219 21097 13231 21131
rect 15010 21128 15016 21140
rect 14971 21100 15016 21128
rect 13173 21091 13231 21097
rect 15010 21088 15016 21100
rect 15068 21088 15074 21140
rect 15565 21131 15623 21137
rect 15565 21097 15577 21131
rect 15611 21128 15623 21131
rect 15838 21128 15844 21140
rect 15611 21100 15844 21128
rect 15611 21097 15623 21100
rect 15565 21091 15623 21097
rect 15838 21088 15844 21100
rect 15896 21088 15902 21140
rect 17037 21131 17095 21137
rect 17037 21097 17049 21131
rect 17083 21097 17095 21131
rect 17037 21091 17095 21097
rect 21085 21131 21143 21137
rect 21085 21097 21097 21131
rect 21131 21128 21143 21131
rect 21910 21128 21916 21140
rect 21131 21100 21916 21128
rect 21131 21097 21143 21100
rect 21085 21091 21143 21097
rect 5160 21063 5218 21069
rect 5160 21029 5172 21063
rect 5206 21060 5218 21063
rect 5258 21060 5264 21072
rect 5206 21032 5264 21060
rect 5206 21029 5218 21032
rect 5160 21023 5218 21029
rect 5258 21020 5264 21032
rect 5316 21020 5322 21072
rect 7742 21060 7748 21072
rect 7703 21032 7748 21060
rect 7742 21020 7748 21032
rect 7800 21020 7806 21072
rect 7929 21063 7987 21069
rect 7929 21029 7941 21063
rect 7975 21029 7987 21063
rect 10686 21060 10692 21072
rect 7929 21023 7987 21029
rect 9692 21032 10692 21060
rect 3510 20952 3516 21004
rect 3568 20992 3574 21004
rect 4893 20995 4951 21001
rect 4893 20992 4905 20995
rect 3568 20964 4905 20992
rect 3568 20952 3574 20964
rect 4893 20961 4905 20964
rect 4939 20992 4951 20995
rect 4982 20992 4988 21004
rect 4939 20964 4988 20992
rect 4939 20961 4951 20964
rect 4893 20955 4951 20961
rect 4982 20952 4988 20964
rect 5040 20952 5046 21004
rect 6730 20952 6736 21004
rect 6788 20992 6794 21004
rect 7944 20992 7972 21023
rect 9692 21001 9720 21032
rect 10686 21020 10692 21032
rect 10744 21020 10750 21072
rect 14182 21060 14188 21072
rect 14143 21032 14188 21060
rect 14182 21020 14188 21032
rect 14240 21020 14246 21072
rect 14274 21020 14280 21072
rect 14332 21060 14338 21072
rect 14332 21032 14377 21060
rect 14332 21020 14338 21032
rect 15654 21020 15660 21072
rect 15712 21060 15718 21072
rect 16482 21060 16488 21072
rect 15712 21032 16488 21060
rect 15712 21020 15718 21032
rect 16482 21020 16488 21032
rect 16540 21060 16546 21072
rect 17052 21060 17080 21091
rect 21910 21088 21916 21100
rect 21968 21088 21974 21140
rect 16540 21032 17080 21060
rect 16540 21020 16546 21032
rect 9950 21001 9956 21004
rect 6788 20964 7972 20992
rect 9677 20995 9735 21001
rect 6788 20952 6794 20964
rect 9677 20961 9689 20995
rect 9723 20961 9735 20995
rect 9944 20992 9956 21001
rect 9911 20964 9956 20992
rect 9677 20955 9735 20961
rect 9944 20955 9956 20964
rect 9950 20952 9956 20955
rect 10008 20952 10014 21004
rect 14001 20995 14059 21001
rect 14001 20961 14013 20995
rect 14047 20992 14059 20995
rect 14090 20992 14096 21004
rect 14047 20964 14096 20992
rect 14047 20961 14059 20964
rect 14001 20955 14059 20961
rect 14090 20952 14096 20964
rect 14148 20992 14154 21004
rect 15746 20992 15752 21004
rect 14148 20964 15752 20992
rect 14148 20952 14154 20964
rect 15746 20952 15752 20964
rect 15804 20952 15810 21004
rect 15930 21001 15936 21004
rect 15924 20992 15936 21001
rect 15891 20964 15936 20992
rect 15924 20955 15936 20964
rect 15930 20952 15936 20955
rect 15988 20952 15994 21004
rect 20898 20992 20904 21004
rect 20859 20964 20904 20992
rect 20898 20952 20904 20964
rect 20956 20952 20962 21004
rect 2314 20924 2320 20936
rect 2275 20896 2320 20924
rect 2314 20884 2320 20896
rect 2372 20884 2378 20936
rect 2501 20927 2559 20933
rect 2501 20893 2513 20927
rect 2547 20924 2559 20927
rect 2682 20924 2688 20936
rect 2547 20896 2688 20924
rect 2547 20893 2559 20896
rect 2501 20887 2559 20893
rect 2682 20884 2688 20896
rect 2740 20884 2746 20936
rect 8021 20927 8079 20933
rect 8021 20893 8033 20927
rect 8067 20924 8079 20927
rect 8294 20924 8300 20936
rect 8067 20896 8300 20924
rect 8067 20893 8079 20896
rect 8021 20887 8079 20893
rect 8294 20884 8300 20896
rect 8352 20884 8358 20936
rect 15654 20924 15660 20936
rect 15615 20896 15660 20924
rect 15654 20884 15660 20896
rect 15712 20884 15718 20936
rect 7469 20859 7527 20865
rect 7469 20825 7481 20859
rect 7515 20856 7527 20859
rect 9030 20856 9036 20868
rect 7515 20828 9036 20856
rect 7515 20825 7527 20828
rect 7469 20819 7527 20825
rect 9030 20816 9036 20828
rect 9088 20816 9094 20868
rect 1673 20791 1731 20797
rect 1673 20757 1685 20791
rect 1719 20788 1731 20791
rect 1854 20788 1860 20800
rect 1719 20760 1860 20788
rect 1719 20757 1731 20760
rect 1673 20751 1731 20757
rect 1854 20748 1860 20760
rect 1912 20748 1918 20800
rect 1949 20791 2007 20797
rect 1949 20757 1961 20791
rect 1995 20788 2007 20791
rect 2498 20788 2504 20800
rect 1995 20760 2504 20788
rect 1995 20757 2007 20760
rect 1949 20751 2007 20757
rect 2498 20748 2504 20760
rect 2556 20748 2562 20800
rect 3145 20791 3203 20797
rect 3145 20757 3157 20791
rect 3191 20788 3203 20791
rect 3694 20788 3700 20800
rect 3191 20760 3700 20788
rect 3191 20757 3203 20760
rect 3145 20751 3203 20757
rect 3694 20748 3700 20760
rect 3752 20748 3758 20800
rect 7285 20791 7343 20797
rect 7285 20757 7297 20791
rect 7331 20788 7343 20791
rect 7374 20788 7380 20800
rect 7331 20760 7380 20788
rect 7331 20757 7343 20760
rect 7285 20751 7343 20757
rect 7374 20748 7380 20760
rect 7432 20748 7438 20800
rect 9401 20791 9459 20797
rect 9401 20757 9413 20791
rect 9447 20788 9459 20791
rect 9582 20788 9588 20800
rect 9447 20760 9588 20788
rect 9447 20757 9459 20760
rect 9401 20751 9459 20757
rect 9582 20748 9588 20760
rect 9640 20748 9646 20800
rect 12894 20788 12900 20800
rect 12855 20760 12900 20788
rect 12894 20748 12900 20760
rect 12952 20748 12958 20800
rect 13630 20748 13636 20800
rect 13688 20788 13694 20800
rect 13725 20791 13783 20797
rect 13725 20788 13737 20791
rect 13688 20760 13737 20788
rect 13688 20748 13694 20760
rect 13725 20757 13737 20760
rect 13771 20757 13783 20791
rect 13725 20751 13783 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 2406 20544 2412 20596
rect 2464 20584 2470 20596
rect 2501 20587 2559 20593
rect 2501 20584 2513 20587
rect 2464 20556 2513 20584
rect 2464 20544 2470 20556
rect 2501 20553 2513 20556
rect 2547 20553 2559 20587
rect 2501 20547 2559 20553
rect 2961 20587 3019 20593
rect 2961 20553 2973 20587
rect 3007 20584 3019 20587
rect 3050 20584 3056 20596
rect 3007 20556 3056 20584
rect 3007 20553 3019 20556
rect 2961 20547 3019 20553
rect 3050 20544 3056 20556
rect 3108 20544 3114 20596
rect 4525 20587 4583 20593
rect 4525 20553 4537 20587
rect 4571 20584 4583 20587
rect 4614 20584 4620 20596
rect 4571 20556 4620 20584
rect 4571 20553 4583 20556
rect 4525 20547 4583 20553
rect 4614 20544 4620 20556
rect 4672 20544 4678 20596
rect 6270 20584 6276 20596
rect 6231 20556 6276 20584
rect 6270 20544 6276 20556
rect 6328 20544 6334 20596
rect 6641 20587 6699 20593
rect 6641 20553 6653 20587
rect 6687 20584 6699 20587
rect 7098 20584 7104 20596
rect 6687 20556 7104 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 3145 20519 3203 20525
rect 3145 20485 3157 20519
rect 3191 20516 3203 20519
rect 4430 20516 4436 20528
rect 3191 20488 4436 20516
rect 3191 20485 3203 20488
rect 3145 20479 3203 20485
rect 4430 20476 4436 20488
rect 4488 20476 4494 20528
rect 4706 20516 4712 20528
rect 4667 20488 4712 20516
rect 4706 20476 4712 20488
rect 4764 20476 4770 20528
rect 3602 20448 3608 20460
rect 3563 20420 3608 20448
rect 3602 20408 3608 20420
rect 3660 20408 3666 20460
rect 5169 20451 5227 20457
rect 5169 20417 5181 20451
rect 5215 20448 5227 20451
rect 5442 20448 5448 20460
rect 5215 20420 5448 20448
rect 5215 20417 5227 20420
rect 5169 20411 5227 20417
rect 5442 20408 5448 20420
rect 5500 20408 5506 20460
rect 1854 20380 1860 20392
rect 1815 20352 1860 20380
rect 1854 20340 1860 20352
rect 1912 20340 1918 20392
rect 3694 20380 3700 20392
rect 3655 20352 3700 20380
rect 3694 20340 3700 20352
rect 3752 20340 3758 20392
rect 4982 20340 4988 20392
rect 5040 20380 5046 20392
rect 6840 20389 6868 20556
rect 7098 20544 7104 20556
rect 7156 20544 7162 20596
rect 8294 20544 8300 20596
rect 8352 20584 8358 20596
rect 8757 20587 8815 20593
rect 8757 20584 8769 20587
rect 8352 20556 8769 20584
rect 8352 20544 8358 20556
rect 8757 20553 8769 20556
rect 8803 20584 8815 20587
rect 9125 20587 9183 20593
rect 9125 20584 9137 20587
rect 8803 20556 9137 20584
rect 8803 20553 8815 20556
rect 8757 20547 8815 20553
rect 9125 20553 9137 20556
rect 9171 20553 9183 20587
rect 9398 20584 9404 20596
rect 9359 20556 9404 20584
rect 9125 20547 9183 20553
rect 9140 20448 9168 20547
rect 9398 20544 9404 20556
rect 9456 20544 9462 20596
rect 10781 20587 10839 20593
rect 10781 20553 10793 20587
rect 10827 20584 10839 20587
rect 10962 20584 10968 20596
rect 10827 20556 10968 20584
rect 10827 20553 10839 20556
rect 10781 20547 10839 20553
rect 10962 20544 10968 20556
rect 11020 20544 11026 20596
rect 11149 20587 11207 20593
rect 11149 20553 11161 20587
rect 11195 20584 11207 20587
rect 11238 20584 11244 20596
rect 11195 20556 11244 20584
rect 11195 20553 11207 20556
rect 11149 20547 11207 20553
rect 11238 20544 11244 20556
rect 11296 20544 11302 20596
rect 13446 20544 13452 20596
rect 13504 20584 13510 20596
rect 13633 20587 13691 20593
rect 13633 20584 13645 20587
rect 13504 20556 13645 20584
rect 13504 20544 13510 20556
rect 13633 20553 13645 20556
rect 13679 20553 13691 20587
rect 14090 20584 14096 20596
rect 14051 20556 14096 20584
rect 13633 20547 13691 20553
rect 14090 20544 14096 20556
rect 14148 20544 14154 20596
rect 14274 20544 14280 20596
rect 14332 20584 14338 20596
rect 14369 20587 14427 20593
rect 14369 20584 14381 20587
rect 14332 20556 14381 20584
rect 14332 20544 14338 20556
rect 14369 20553 14381 20556
rect 14415 20553 14427 20587
rect 14369 20547 14427 20553
rect 12526 20516 12532 20528
rect 12487 20488 12532 20516
rect 12526 20476 12532 20488
rect 12584 20476 12590 20528
rect 9950 20448 9956 20460
rect 9140 20420 9956 20448
rect 9950 20408 9956 20420
rect 10008 20408 10014 20460
rect 12894 20408 12900 20460
rect 12952 20448 12958 20460
rect 12989 20451 13047 20457
rect 12989 20448 13001 20451
rect 12952 20420 13001 20448
rect 12952 20408 12958 20420
rect 12989 20417 13001 20420
rect 13035 20448 13047 20451
rect 13722 20448 13728 20460
rect 13035 20420 13728 20448
rect 13035 20417 13047 20420
rect 12989 20411 13047 20417
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 18322 20448 18328 20460
rect 18283 20420 18328 20448
rect 18322 20408 18328 20420
rect 18380 20408 18386 20460
rect 5721 20383 5779 20389
rect 5721 20380 5733 20383
rect 5040 20352 5733 20380
rect 5040 20340 5046 20352
rect 5721 20349 5733 20352
rect 5767 20380 5779 20383
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 5767 20352 6837 20380
rect 5767 20349 5779 20352
rect 5721 20343 5779 20349
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 12069 20383 12127 20389
rect 12069 20349 12081 20383
rect 12115 20380 12127 20383
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 12115 20352 13093 20380
rect 12115 20349 12127 20352
rect 12069 20343 12127 20349
rect 13081 20349 13093 20352
rect 13127 20349 13139 20383
rect 13081 20343 13139 20349
rect 14645 20383 14703 20389
rect 14645 20349 14657 20383
rect 14691 20380 14703 20383
rect 14921 20383 14979 20389
rect 14921 20380 14933 20383
rect 14691 20352 14933 20380
rect 14691 20349 14703 20352
rect 14645 20343 14703 20349
rect 14921 20349 14933 20352
rect 14967 20380 14979 20383
rect 15654 20380 15660 20392
rect 14967 20352 15660 20380
rect 14967 20349 14979 20352
rect 14921 20343 14979 20349
rect 15654 20340 15660 20352
rect 15712 20340 15718 20392
rect 18046 20380 18052 20392
rect 18007 20352 18052 20380
rect 18046 20340 18052 20352
rect 18104 20380 18110 20392
rect 18785 20383 18843 20389
rect 18785 20380 18797 20383
rect 18104 20352 18797 20380
rect 18104 20340 18110 20352
rect 18785 20349 18797 20352
rect 18831 20349 18843 20383
rect 18785 20343 18843 20349
rect 2133 20315 2191 20321
rect 2133 20281 2145 20315
rect 2179 20312 2191 20315
rect 2682 20312 2688 20324
rect 2179 20284 2688 20312
rect 2179 20281 2191 20284
rect 2133 20275 2191 20281
rect 2682 20272 2688 20284
rect 2740 20272 2746 20324
rect 3142 20272 3148 20324
rect 3200 20312 3206 20324
rect 3605 20315 3663 20321
rect 3605 20312 3617 20315
rect 3200 20284 3617 20312
rect 3200 20272 3206 20284
rect 3605 20281 3617 20284
rect 3651 20281 3663 20315
rect 5261 20315 5319 20321
rect 5261 20312 5273 20315
rect 3605 20275 3663 20281
rect 4172 20284 5273 20312
rect 4172 20256 4200 20284
rect 5261 20281 5273 20284
rect 5307 20281 5319 20315
rect 5261 20275 5319 20281
rect 6270 20272 6276 20324
rect 6328 20312 6334 20324
rect 7070 20315 7128 20321
rect 7070 20312 7082 20315
rect 6328 20284 7082 20312
rect 6328 20272 6334 20284
rect 7070 20281 7082 20284
rect 7116 20281 7128 20315
rect 9674 20312 9680 20324
rect 9635 20284 9680 20312
rect 7070 20275 7128 20281
rect 9674 20272 9680 20284
rect 9732 20272 9738 20324
rect 12894 20272 12900 20324
rect 12952 20312 12958 20324
rect 12989 20315 13047 20321
rect 12989 20312 13001 20315
rect 12952 20284 13001 20312
rect 12952 20272 12958 20284
rect 12989 20281 13001 20284
rect 13035 20281 13047 20315
rect 12989 20275 13047 20281
rect 14274 20272 14280 20324
rect 14332 20312 14338 20324
rect 15166 20315 15224 20321
rect 15166 20312 15178 20315
rect 14332 20284 15178 20312
rect 14332 20272 14338 20284
rect 15166 20281 15178 20284
rect 15212 20281 15224 20315
rect 15166 20275 15224 20281
rect 1762 20204 1768 20256
rect 1820 20244 1826 20256
rect 2041 20247 2099 20253
rect 2041 20244 2053 20247
rect 1820 20216 2053 20244
rect 1820 20204 1826 20216
rect 2041 20213 2053 20216
rect 2087 20213 2099 20247
rect 4154 20244 4160 20256
rect 4115 20216 4160 20244
rect 2041 20207 2099 20213
rect 4154 20204 4160 20216
rect 4212 20204 4218 20256
rect 4614 20204 4620 20256
rect 4672 20244 4678 20256
rect 5169 20247 5227 20253
rect 5169 20244 5181 20247
rect 4672 20216 5181 20244
rect 4672 20204 4678 20216
rect 5169 20213 5181 20216
rect 5215 20213 5227 20247
rect 8202 20244 8208 20256
rect 8163 20216 8208 20244
rect 5169 20207 5227 20213
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 9490 20204 9496 20256
rect 9548 20244 9554 20256
rect 9861 20247 9919 20253
rect 9861 20244 9873 20247
rect 9548 20216 9873 20244
rect 9548 20204 9554 20216
rect 9861 20213 9873 20216
rect 9907 20213 9919 20247
rect 9861 20207 9919 20213
rect 10413 20247 10471 20253
rect 10413 20213 10425 20247
rect 10459 20244 10471 20247
rect 10686 20244 10692 20256
rect 10459 20216 10692 20244
rect 10459 20213 10471 20216
rect 10413 20207 10471 20213
rect 10686 20204 10692 20216
rect 10744 20244 10750 20256
rect 11238 20244 11244 20256
rect 10744 20216 11244 20244
rect 10744 20204 10750 20216
rect 11238 20204 11244 20216
rect 11296 20204 11302 20256
rect 11790 20244 11796 20256
rect 11751 20216 11796 20244
rect 11790 20204 11796 20216
rect 11848 20204 11854 20256
rect 11882 20204 11888 20256
rect 11940 20244 11946 20256
rect 12069 20247 12127 20253
rect 12069 20244 12081 20247
rect 11940 20216 12081 20244
rect 11940 20204 11946 20216
rect 12069 20213 12081 20216
rect 12115 20244 12127 20247
rect 12161 20247 12219 20253
rect 12161 20244 12173 20247
rect 12115 20216 12173 20244
rect 12115 20213 12127 20216
rect 12069 20207 12127 20213
rect 12161 20213 12173 20216
rect 12207 20213 12219 20247
rect 12161 20207 12219 20213
rect 13446 20204 13452 20256
rect 13504 20244 13510 20256
rect 14645 20247 14703 20253
rect 14645 20244 14657 20247
rect 13504 20216 14657 20244
rect 13504 20204 13510 20216
rect 14645 20213 14657 20216
rect 14691 20244 14703 20247
rect 14737 20247 14795 20253
rect 14737 20244 14749 20247
rect 14691 20216 14749 20244
rect 14691 20213 14703 20216
rect 14645 20207 14703 20213
rect 14737 20213 14749 20216
rect 14783 20213 14795 20247
rect 14737 20207 14795 20213
rect 16022 20204 16028 20256
rect 16080 20244 16086 20256
rect 16301 20247 16359 20253
rect 16301 20244 16313 20247
rect 16080 20216 16313 20244
rect 16080 20204 16086 20216
rect 16301 20213 16313 20216
rect 16347 20213 16359 20247
rect 20898 20244 20904 20256
rect 20859 20216 20904 20244
rect 16301 20207 16359 20213
rect 20898 20204 20904 20216
rect 20956 20204 20962 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1857 20043 1915 20049
rect 1857 20009 1869 20043
rect 1903 20040 1915 20043
rect 2314 20040 2320 20052
rect 1903 20012 2320 20040
rect 1903 20009 1915 20012
rect 1857 20003 1915 20009
rect 2314 20000 2320 20012
rect 2372 20000 2378 20052
rect 3145 20043 3203 20049
rect 3145 20009 3157 20043
rect 3191 20040 3203 20043
rect 3602 20040 3608 20052
rect 3191 20012 3608 20040
rect 3191 20009 3203 20012
rect 3145 20003 3203 20009
rect 3602 20000 3608 20012
rect 3660 20000 3666 20052
rect 5258 20040 5264 20052
rect 5219 20012 5264 20040
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 6549 20043 6607 20049
rect 6549 20009 6561 20043
rect 6595 20040 6607 20043
rect 6730 20040 6736 20052
rect 6595 20012 6736 20040
rect 6595 20009 6607 20012
rect 6549 20003 6607 20009
rect 6730 20000 6736 20012
rect 6788 20000 6794 20052
rect 6914 20040 6920 20052
rect 6875 20012 6920 20040
rect 6914 20000 6920 20012
rect 6972 20000 6978 20052
rect 8294 20000 8300 20052
rect 8352 20040 8358 20052
rect 8481 20043 8539 20049
rect 8481 20040 8493 20043
rect 8352 20012 8493 20040
rect 8352 20000 8358 20012
rect 8481 20009 8493 20012
rect 8527 20009 8539 20043
rect 8481 20003 8539 20009
rect 9950 20000 9956 20052
rect 10008 20040 10014 20052
rect 10137 20043 10195 20049
rect 10137 20040 10149 20043
rect 10008 20012 10149 20040
rect 10008 20000 10014 20012
rect 10137 20009 10149 20012
rect 10183 20009 10195 20043
rect 10778 20040 10784 20052
rect 10739 20012 10784 20040
rect 10137 20003 10195 20009
rect 10778 20000 10784 20012
rect 10836 20040 10842 20052
rect 11054 20040 11060 20052
rect 10836 20012 11060 20040
rect 10836 20000 10842 20012
rect 11054 20000 11060 20012
rect 11112 20000 11118 20052
rect 11790 20000 11796 20052
rect 11848 20040 11854 20052
rect 12894 20040 12900 20052
rect 11848 20012 12900 20040
rect 11848 20000 11854 20012
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 13541 20043 13599 20049
rect 13541 20009 13553 20043
rect 13587 20040 13599 20043
rect 15654 20040 15660 20052
rect 13587 20012 14320 20040
rect 15615 20012 15660 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 14292 19984 14320 20012
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 2958 19932 2964 19984
rect 3016 19972 3022 19984
rect 3421 19975 3479 19981
rect 3421 19972 3433 19975
rect 3016 19944 3433 19972
rect 3016 19932 3022 19944
rect 3421 19941 3433 19944
rect 3467 19941 3479 19975
rect 4706 19972 4712 19984
rect 4619 19944 4712 19972
rect 3421 19935 3479 19941
rect 4706 19932 4712 19944
rect 4764 19972 4770 19984
rect 5166 19972 5172 19984
rect 4764 19944 5172 19972
rect 4764 19932 4770 19944
rect 5166 19932 5172 19944
rect 5224 19932 5230 19984
rect 10226 19932 10232 19984
rect 10284 19972 10290 19984
rect 12802 19972 12808 19984
rect 10284 19944 12808 19972
rect 10284 19932 10290 19944
rect 12802 19932 12808 19944
rect 12860 19932 12866 19984
rect 14182 19972 14188 19984
rect 14143 19944 14188 19972
rect 14182 19932 14188 19944
rect 14240 19932 14246 19984
rect 14274 19932 14280 19984
rect 14332 19972 14338 19984
rect 14921 19975 14979 19981
rect 14921 19972 14933 19975
rect 14332 19944 14933 19972
rect 14332 19932 14338 19944
rect 14921 19941 14933 19944
rect 14967 19941 14979 19975
rect 14921 19935 14979 19941
rect 7098 19904 7104 19916
rect 7059 19876 7104 19904
rect 7098 19864 7104 19876
rect 7156 19864 7162 19916
rect 7374 19913 7380 19916
rect 7368 19904 7380 19913
rect 7287 19876 7380 19904
rect 7368 19867 7380 19876
rect 7432 19904 7438 19916
rect 8202 19904 8208 19916
rect 7432 19876 8208 19904
rect 7374 19864 7380 19867
rect 7432 19864 7438 19876
rect 8202 19864 8208 19876
rect 8260 19864 8266 19916
rect 11149 19907 11207 19913
rect 11149 19873 11161 19907
rect 11195 19904 11207 19907
rect 11238 19904 11244 19916
rect 11195 19876 11244 19904
rect 11195 19873 11207 19876
rect 11149 19867 11207 19873
rect 11238 19864 11244 19876
rect 11296 19864 11302 19916
rect 11422 19913 11428 19916
rect 11416 19904 11428 19913
rect 11383 19876 11428 19904
rect 11416 19867 11428 19876
rect 11422 19864 11428 19867
rect 11480 19864 11486 19916
rect 13814 19864 13820 19916
rect 13872 19904 13878 19916
rect 14001 19907 14059 19913
rect 14001 19904 14013 19907
rect 13872 19876 14013 19904
rect 13872 19864 13878 19876
rect 14001 19873 14013 19876
rect 14047 19873 14059 19907
rect 15672 19904 15700 20000
rect 16482 19981 16488 19984
rect 16476 19972 16488 19981
rect 16443 19944 16488 19972
rect 16476 19935 16488 19944
rect 16482 19932 16488 19935
rect 16540 19932 16546 19984
rect 19429 19975 19487 19981
rect 19429 19941 19441 19975
rect 19475 19972 19487 19975
rect 20898 19972 20904 19984
rect 19475 19944 20904 19972
rect 19475 19941 19487 19944
rect 19429 19935 19487 19941
rect 20898 19932 20904 19944
rect 20956 19932 20962 19984
rect 16209 19907 16267 19913
rect 16209 19904 16221 19907
rect 15672 19876 16221 19904
rect 14001 19867 14059 19873
rect 16209 19873 16221 19876
rect 16255 19904 16267 19907
rect 16298 19904 16304 19916
rect 16255 19876 16304 19904
rect 16255 19873 16267 19876
rect 16209 19867 16267 19873
rect 16298 19864 16304 19876
rect 16356 19864 16362 19916
rect 19150 19904 19156 19916
rect 19111 19876 19156 19904
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 4798 19836 4804 19848
rect 4759 19808 4804 19836
rect 4617 19799 4675 19805
rect 4632 19768 4660 19799
rect 4798 19796 4804 19808
rect 4856 19796 4862 19848
rect 9677 19839 9735 19845
rect 9677 19805 9689 19839
rect 9723 19836 9735 19839
rect 9766 19836 9772 19848
rect 9723 19808 9772 19836
rect 9723 19805 9735 19808
rect 9677 19799 9735 19805
rect 9766 19796 9772 19808
rect 9824 19796 9830 19848
rect 5442 19768 5448 19780
rect 4632 19740 5448 19768
rect 5442 19728 5448 19740
rect 5500 19728 5506 19780
rect 15838 19728 15844 19780
rect 15896 19768 15902 19780
rect 16114 19768 16120 19780
rect 15896 19740 16120 19768
rect 15896 19728 15902 19740
rect 16114 19728 16120 19740
rect 16172 19728 16178 19780
rect 17586 19768 17592 19780
rect 17547 19740 17592 19768
rect 17586 19728 17592 19740
rect 17644 19728 17650 19780
rect 1673 19703 1731 19709
rect 1673 19669 1685 19703
rect 1719 19700 1731 19703
rect 1762 19700 1768 19712
rect 1719 19672 1768 19700
rect 1719 19669 1731 19672
rect 1673 19663 1731 19669
rect 1762 19660 1768 19672
rect 1820 19660 1826 19712
rect 2682 19700 2688 19712
rect 2643 19672 2688 19700
rect 2682 19660 2688 19672
rect 2740 19660 2746 19712
rect 3786 19700 3792 19712
rect 3747 19672 3792 19700
rect 3786 19660 3792 19672
rect 3844 19660 3850 19712
rect 4246 19700 4252 19712
rect 4207 19672 4252 19700
rect 4246 19660 4252 19672
rect 4304 19660 4310 19712
rect 9401 19703 9459 19709
rect 9401 19669 9413 19703
rect 9447 19700 9459 19703
rect 9490 19700 9496 19712
rect 9447 19672 9496 19700
rect 9447 19669 9459 19672
rect 9401 19663 9459 19669
rect 9490 19660 9496 19672
rect 9548 19700 9554 19712
rect 9858 19700 9864 19712
rect 9548 19672 9864 19700
rect 9548 19660 9554 19672
rect 9858 19660 9864 19672
rect 9916 19660 9922 19712
rect 12529 19703 12587 19709
rect 12529 19669 12541 19703
rect 12575 19700 12587 19703
rect 12894 19700 12900 19712
rect 12575 19672 12900 19700
rect 12575 19669 12587 19672
rect 12529 19663 12587 19669
rect 12894 19660 12900 19672
rect 12952 19660 12958 19712
rect 13722 19700 13728 19712
rect 13683 19672 13728 19700
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 15562 19660 15568 19712
rect 15620 19700 15626 19712
rect 16022 19700 16028 19712
rect 15620 19672 16028 19700
rect 15620 19660 15626 19672
rect 16022 19660 16028 19672
rect 16080 19660 16086 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1673 19499 1731 19505
rect 1673 19465 1685 19499
rect 1719 19496 1731 19499
rect 2682 19496 2688 19508
rect 1719 19468 2688 19496
rect 1719 19465 1731 19468
rect 1673 19459 1731 19465
rect 2682 19456 2688 19468
rect 2740 19456 2746 19508
rect 5166 19496 5172 19508
rect 5127 19468 5172 19496
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 7098 19456 7104 19508
rect 7156 19496 7162 19508
rect 7837 19499 7895 19505
rect 7837 19496 7849 19499
rect 7156 19468 7849 19496
rect 7156 19456 7162 19468
rect 7837 19465 7849 19468
rect 7883 19465 7895 19499
rect 7837 19459 7895 19465
rect 9033 19499 9091 19505
rect 9033 19465 9045 19499
rect 9079 19496 9091 19499
rect 9674 19496 9680 19508
rect 9079 19468 9680 19496
rect 9079 19465 9091 19468
rect 9033 19459 9091 19465
rect 9674 19456 9680 19468
rect 9732 19456 9738 19508
rect 10873 19499 10931 19505
rect 10873 19465 10885 19499
rect 10919 19496 10931 19499
rect 11790 19496 11796 19508
rect 10919 19468 11796 19496
rect 10919 19465 10931 19468
rect 10873 19459 10931 19465
rect 11790 19456 11796 19468
rect 11848 19456 11854 19508
rect 13354 19456 13360 19508
rect 13412 19456 13418 19508
rect 13814 19456 13820 19508
rect 13872 19496 13878 19508
rect 14369 19499 14427 19505
rect 14369 19496 14381 19499
rect 13872 19468 14381 19496
rect 13872 19456 13878 19468
rect 14369 19465 14381 19468
rect 14415 19465 14427 19499
rect 14369 19459 14427 19465
rect 14734 19456 14740 19508
rect 14792 19496 14798 19508
rect 15013 19499 15071 19505
rect 15013 19496 15025 19499
rect 14792 19468 15025 19496
rect 14792 19456 14798 19468
rect 15013 19465 15025 19468
rect 15059 19465 15071 19499
rect 16298 19496 16304 19508
rect 16259 19468 16304 19496
rect 15013 19459 15071 19465
rect 16298 19456 16304 19468
rect 16356 19456 16362 19508
rect 16482 19456 16488 19508
rect 16540 19496 16546 19508
rect 16577 19499 16635 19505
rect 16577 19496 16589 19499
rect 16540 19468 16589 19496
rect 16540 19456 16546 19468
rect 16577 19465 16589 19468
rect 16623 19465 16635 19499
rect 16577 19459 16635 19465
rect 2317 19431 2375 19437
rect 2317 19397 2329 19431
rect 2363 19397 2375 19431
rect 13372 19428 13400 19456
rect 14458 19428 14464 19440
rect 13372 19400 14464 19428
rect 2317 19391 2375 19397
rect 2332 19292 2360 19391
rect 14458 19388 14464 19400
rect 14516 19388 14522 19440
rect 2774 19320 2780 19372
rect 2832 19360 2838 19372
rect 3786 19360 3792 19372
rect 2832 19332 3792 19360
rect 2832 19320 2838 19332
rect 3786 19320 3792 19332
rect 3844 19360 3850 19372
rect 3844 19332 4108 19360
rect 3844 19320 3850 19332
rect 2406 19292 2412 19304
rect 2332 19264 2412 19292
rect 2406 19252 2412 19264
rect 2464 19252 2470 19304
rect 4080 19292 4108 19332
rect 4338 19320 4344 19372
rect 4396 19360 4402 19372
rect 4798 19360 4804 19372
rect 4396 19332 4804 19360
rect 4396 19320 4402 19332
rect 4798 19320 4804 19332
rect 4856 19320 4862 19372
rect 8202 19360 8208 19372
rect 6840 19332 8208 19360
rect 4157 19295 4215 19301
rect 4157 19292 4169 19295
rect 4080 19264 4169 19292
rect 4157 19261 4169 19264
rect 4203 19261 4215 19295
rect 5626 19292 5632 19304
rect 5587 19264 5632 19292
rect 4157 19255 4215 19261
rect 5626 19252 5632 19264
rect 5684 19252 5690 19304
rect 6273 19295 6331 19301
rect 6273 19261 6285 19295
rect 6319 19292 6331 19295
rect 6840 19292 6868 19332
rect 8202 19320 8208 19332
rect 8260 19320 8266 19372
rect 9493 19363 9551 19369
rect 9493 19329 9505 19363
rect 9539 19360 9551 19363
rect 9766 19360 9772 19372
rect 9539 19332 9772 19360
rect 9539 19329 9551 19332
rect 9493 19323 9551 19329
rect 6319 19264 6868 19292
rect 6319 19261 6331 19264
rect 6273 19255 6331 19261
rect 6914 19252 6920 19304
rect 6972 19292 6978 19304
rect 7193 19295 7251 19301
rect 7193 19292 7205 19295
rect 6972 19264 7205 19292
rect 6972 19252 6978 19264
rect 7193 19261 7205 19264
rect 7239 19261 7251 19295
rect 7193 19255 7251 19261
rect 9030 19252 9036 19304
rect 9088 19292 9094 19304
rect 9508 19292 9536 19323
rect 9766 19320 9772 19332
rect 9824 19320 9830 19372
rect 13446 19320 13452 19372
rect 13504 19360 13510 19372
rect 13504 19332 13768 19360
rect 13504 19320 13510 19332
rect 10594 19292 10600 19304
rect 9088 19264 9536 19292
rect 10555 19264 10600 19292
rect 9088 19252 9094 19264
rect 10594 19252 10600 19264
rect 10652 19252 10658 19304
rect 11238 19252 11244 19304
rect 11296 19292 11302 19304
rect 12342 19292 12348 19304
rect 11296 19264 12348 19292
rect 11296 19252 11302 19264
rect 12342 19252 12348 19264
rect 12400 19292 12406 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 12400 19264 12449 19292
rect 12400 19252 12406 19264
rect 12437 19261 12449 19264
rect 12483 19292 12495 19295
rect 13740 19292 13768 19332
rect 15286 19292 15292 19304
rect 12483 19264 13768 19292
rect 15247 19264 15292 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 15286 19252 15292 19264
rect 15344 19292 15350 19304
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 15344 19264 16957 19292
rect 15344 19252 15350 19264
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 16945 19255 17003 19261
rect 21542 19252 21548 19304
rect 21600 19292 21606 19304
rect 22281 19295 22339 19301
rect 22281 19292 22293 19295
rect 21600 19264 22293 19292
rect 21600 19252 21606 19264
rect 22281 19261 22293 19264
rect 22327 19292 22339 19295
rect 22833 19295 22891 19301
rect 22833 19292 22845 19295
rect 22327 19264 22845 19292
rect 22327 19261 22339 19264
rect 22281 19255 22339 19261
rect 22833 19261 22845 19264
rect 22879 19261 22891 19295
rect 22833 19255 22891 19261
rect 2314 19184 2320 19236
rect 2372 19224 2378 19236
rect 2593 19227 2651 19233
rect 2593 19224 2605 19227
rect 2372 19196 2605 19224
rect 2372 19184 2378 19196
rect 2593 19193 2605 19196
rect 2639 19193 2651 19227
rect 2593 19187 2651 19193
rect 2869 19227 2927 19233
rect 2869 19193 2881 19227
rect 2915 19224 2927 19227
rect 3863 19227 3921 19233
rect 2915 19196 3372 19224
rect 2915 19193 2927 19196
rect 2869 19187 2927 19193
rect 3344 19168 3372 19196
rect 3863 19193 3875 19227
rect 3909 19224 3921 19227
rect 4062 19224 4068 19236
rect 3909 19196 4068 19224
rect 3909 19193 3921 19196
rect 3863 19187 3921 19193
rect 4062 19184 4068 19196
rect 4120 19184 4126 19236
rect 4246 19184 4252 19236
rect 4304 19224 4310 19236
rect 4341 19227 4399 19233
rect 4341 19224 4353 19227
rect 4304 19196 4353 19224
rect 4304 19184 4310 19196
rect 4341 19193 4353 19196
rect 4387 19193 4399 19227
rect 4341 19187 4399 19193
rect 4433 19227 4491 19233
rect 4433 19193 4445 19227
rect 4479 19193 4491 19227
rect 4433 19187 4491 19193
rect 2133 19159 2191 19165
rect 2133 19125 2145 19159
rect 2179 19156 2191 19159
rect 2777 19159 2835 19165
rect 2777 19156 2789 19159
rect 2179 19128 2789 19156
rect 2179 19125 2191 19128
rect 2133 19119 2191 19125
rect 2777 19125 2789 19128
rect 2823 19156 2835 19159
rect 2958 19156 2964 19168
rect 2823 19128 2964 19156
rect 2823 19125 2835 19128
rect 2777 19119 2835 19125
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 3326 19156 3332 19168
rect 3287 19128 3332 19156
rect 3326 19116 3332 19128
rect 3384 19116 3390 19168
rect 3697 19159 3755 19165
rect 3697 19125 3709 19159
rect 3743 19156 3755 19159
rect 4448 19156 4476 19187
rect 5994 19184 6000 19236
rect 6052 19224 6058 19236
rect 6641 19227 6699 19233
rect 6641 19224 6653 19227
rect 6052 19196 6653 19224
rect 6052 19184 6058 19196
rect 6641 19193 6653 19196
rect 6687 19224 6699 19227
rect 7377 19227 7435 19233
rect 7377 19224 7389 19227
rect 6687 19196 7389 19224
rect 6687 19193 6699 19196
rect 6641 19187 6699 19193
rect 7377 19193 7389 19196
rect 7423 19193 7435 19227
rect 7377 19187 7435 19193
rect 7469 19227 7527 19233
rect 7469 19193 7481 19227
rect 7515 19224 7527 19227
rect 7558 19224 7564 19236
rect 7515 19196 7564 19224
rect 7515 19193 7527 19196
rect 7469 19187 7527 19193
rect 7558 19184 7564 19196
rect 7616 19184 7622 19236
rect 8202 19184 8208 19236
rect 8260 19224 8266 19236
rect 8481 19227 8539 19233
rect 8481 19224 8493 19227
rect 8260 19196 8493 19224
rect 8260 19184 8266 19196
rect 8481 19193 8493 19196
rect 8527 19224 8539 19227
rect 9585 19227 9643 19233
rect 9585 19224 9597 19227
rect 8527 19196 9597 19224
rect 8527 19193 8539 19196
rect 8481 19187 8539 19193
rect 9585 19193 9597 19196
rect 9631 19224 9643 19227
rect 10042 19224 10048 19236
rect 9631 19196 10048 19224
rect 9631 19193 9643 19196
rect 9585 19187 9643 19193
rect 10042 19184 10048 19196
rect 10100 19184 10106 19236
rect 10226 19184 10232 19236
rect 10284 19184 10290 19236
rect 10321 19227 10379 19233
rect 10321 19193 10333 19227
rect 10367 19224 10379 19227
rect 11146 19224 11152 19236
rect 10367 19196 11152 19224
rect 10367 19193 10379 19196
rect 10321 19187 10379 19193
rect 11146 19184 11152 19196
rect 11204 19184 11210 19236
rect 11422 19224 11428 19236
rect 11383 19196 11428 19224
rect 11422 19184 11428 19196
rect 11480 19224 11486 19236
rect 12704 19227 12762 19233
rect 12704 19224 12716 19227
rect 11480 19196 12716 19224
rect 11480 19184 11486 19196
rect 12704 19193 12716 19196
rect 12750 19224 12762 19227
rect 12894 19224 12900 19236
rect 12750 19196 12900 19224
rect 12750 19193 12762 19196
rect 12704 19187 12762 19193
rect 12894 19184 12900 19196
rect 12952 19184 12958 19236
rect 15470 19224 15476 19236
rect 15431 19196 15476 19224
rect 15470 19184 15476 19196
rect 15528 19184 15534 19236
rect 15562 19184 15568 19236
rect 15620 19224 15626 19236
rect 15620 19196 15713 19224
rect 15620 19184 15626 19196
rect 5442 19156 5448 19168
rect 3743 19128 5448 19156
rect 3743 19125 3755 19128
rect 3697 19119 3755 19125
rect 5442 19116 5448 19128
rect 5500 19116 5506 19168
rect 6907 19159 6965 19165
rect 6907 19125 6919 19159
rect 6953 19156 6965 19159
rect 7098 19156 7104 19168
rect 6953 19128 7104 19156
rect 6953 19125 6965 19128
rect 6907 19119 6965 19125
rect 7098 19116 7104 19128
rect 7156 19116 7162 19168
rect 8754 19156 8760 19168
rect 8715 19128 8760 19156
rect 8754 19116 8760 19128
rect 8812 19156 8818 19168
rect 9493 19159 9551 19165
rect 9493 19156 9505 19159
rect 8812 19128 9505 19156
rect 8812 19116 8818 19128
rect 9493 19125 9505 19128
rect 9539 19125 9551 19159
rect 9493 19119 9551 19125
rect 9766 19116 9772 19168
rect 9824 19156 9830 19168
rect 10244 19156 10272 19184
rect 9824 19128 10272 19156
rect 9824 19116 9830 19128
rect 11054 19116 11060 19168
rect 11112 19156 11118 19168
rect 11333 19159 11391 19165
rect 11333 19156 11345 19159
rect 11112 19128 11345 19156
rect 11112 19116 11118 19128
rect 11333 19125 11345 19128
rect 11379 19125 11391 19159
rect 11333 19119 11391 19125
rect 11885 19159 11943 19165
rect 11885 19125 11897 19159
rect 11931 19156 11943 19159
rect 12253 19159 12311 19165
rect 12253 19156 12265 19159
rect 11931 19128 12265 19156
rect 11931 19125 11943 19128
rect 11885 19119 11943 19125
rect 12253 19125 12265 19128
rect 12299 19156 12311 19159
rect 12342 19156 12348 19168
rect 12299 19128 12348 19156
rect 12299 19125 12311 19128
rect 12253 19119 12311 19125
rect 12342 19116 12348 19128
rect 12400 19156 12406 19168
rect 12618 19156 12624 19168
rect 12400 19128 12624 19156
rect 12400 19116 12406 19128
rect 12618 19116 12624 19128
rect 12676 19116 12682 19168
rect 13814 19156 13820 19168
rect 13775 19128 13820 19156
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 14274 19116 14280 19168
rect 14332 19156 14338 19168
rect 14737 19159 14795 19165
rect 14737 19156 14749 19159
rect 14332 19128 14749 19156
rect 14332 19116 14338 19128
rect 14737 19125 14749 19128
rect 14783 19125 14795 19159
rect 14737 19119 14795 19125
rect 15010 19116 15016 19168
rect 15068 19156 15074 19168
rect 15580 19156 15608 19184
rect 19150 19156 19156 19168
rect 15068 19128 15608 19156
rect 19111 19128 19156 19156
rect 15068 19116 15074 19128
rect 19150 19116 19156 19128
rect 19208 19116 19214 19168
rect 22465 19159 22523 19165
rect 22465 19125 22477 19159
rect 22511 19156 22523 19159
rect 23382 19156 23388 19168
rect 22511 19128 23388 19156
rect 22511 19125 22523 19128
rect 22465 19119 22523 19125
rect 23382 19116 23388 19128
rect 23440 19116 23446 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2314 18952 2320 18964
rect 2275 18924 2320 18952
rect 2314 18912 2320 18924
rect 2372 18912 2378 18964
rect 3881 18955 3939 18961
rect 3881 18921 3893 18955
rect 3927 18952 3939 18955
rect 4246 18952 4252 18964
rect 3927 18924 4252 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 4246 18912 4252 18924
rect 4304 18912 4310 18964
rect 5442 18952 5448 18964
rect 5403 18924 5448 18952
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 7558 18952 7564 18964
rect 7519 18924 7564 18952
rect 7558 18912 7564 18924
rect 7616 18912 7622 18964
rect 9030 18952 9036 18964
rect 8991 18924 9036 18952
rect 9030 18912 9036 18924
rect 9088 18912 9094 18964
rect 10873 18955 10931 18961
rect 10873 18921 10885 18955
rect 10919 18952 10931 18955
rect 11422 18952 11428 18964
rect 10919 18924 11428 18952
rect 10919 18921 10931 18924
rect 10873 18915 10931 18921
rect 11422 18912 11428 18924
rect 11480 18912 11486 18964
rect 15010 18952 15016 18964
rect 14971 18924 15016 18952
rect 15010 18912 15016 18924
rect 15068 18912 15074 18964
rect 15470 18912 15476 18964
rect 15528 18952 15534 18964
rect 16301 18955 16359 18961
rect 16301 18952 16313 18955
rect 15528 18924 16313 18952
rect 15528 18912 15534 18924
rect 16301 18921 16313 18924
rect 16347 18921 16359 18955
rect 16301 18915 16359 18921
rect 2498 18844 2504 18896
rect 2556 18884 2562 18896
rect 2961 18887 3019 18893
rect 2961 18884 2973 18887
rect 2556 18856 2973 18884
rect 2556 18844 2562 18856
rect 2961 18853 2973 18856
rect 3007 18853 3019 18887
rect 2961 18847 3019 18853
rect 3326 18844 3332 18896
rect 3384 18884 3390 18896
rect 4154 18884 4160 18896
rect 3384 18856 4160 18884
rect 3384 18844 3390 18856
rect 4154 18844 4160 18856
rect 4212 18844 4218 18896
rect 7098 18884 7104 18896
rect 7059 18856 7104 18884
rect 7098 18844 7104 18856
rect 7156 18844 7162 18896
rect 10229 18887 10287 18893
rect 10229 18853 10241 18887
rect 10275 18884 10287 18887
rect 10686 18884 10692 18896
rect 10275 18856 10692 18884
rect 10275 18853 10287 18856
rect 10229 18847 10287 18853
rect 10686 18844 10692 18856
rect 10744 18844 10750 18896
rect 11238 18884 11244 18896
rect 11199 18856 11244 18884
rect 11238 18844 11244 18856
rect 11296 18844 11302 18896
rect 14734 18844 14740 18896
rect 14792 18884 14798 18896
rect 15841 18887 15899 18893
rect 15841 18884 15853 18887
rect 14792 18856 15853 18884
rect 14792 18844 14798 18856
rect 15841 18853 15853 18856
rect 15887 18853 15899 18887
rect 15841 18847 15899 18853
rect 15930 18844 15936 18896
rect 15988 18884 15994 18896
rect 15988 18856 16033 18884
rect 15988 18844 15994 18856
rect 2406 18776 2412 18828
rect 2464 18816 2470 18828
rect 4338 18825 4344 18828
rect 2777 18819 2835 18825
rect 2777 18816 2789 18819
rect 2464 18788 2789 18816
rect 2464 18776 2470 18788
rect 2777 18785 2789 18788
rect 2823 18785 2835 18819
rect 4321 18819 4344 18825
rect 4321 18816 4333 18819
rect 2777 18779 2835 18785
rect 3068 18788 4333 18816
rect 3068 18760 3096 18788
rect 4321 18785 4333 18788
rect 4396 18816 4402 18828
rect 6457 18819 6515 18825
rect 4396 18788 4469 18816
rect 4321 18779 4344 18785
rect 4338 18776 4344 18779
rect 4396 18776 4402 18788
rect 6457 18785 6469 18819
rect 6503 18816 6515 18819
rect 6914 18816 6920 18828
rect 6503 18788 6920 18816
rect 6503 18785 6515 18788
rect 6457 18779 6515 18785
rect 6914 18776 6920 18788
rect 6972 18776 6978 18828
rect 10042 18776 10048 18828
rect 10100 18816 10106 18828
rect 10321 18819 10379 18825
rect 10321 18816 10333 18819
rect 10100 18788 10333 18816
rect 10100 18776 10106 18788
rect 10321 18785 10333 18788
rect 10367 18785 10379 18819
rect 10321 18779 10379 18785
rect 11882 18776 11888 18828
rect 11940 18816 11946 18828
rect 12980 18819 13038 18825
rect 12980 18816 12992 18819
rect 11940 18788 12992 18816
rect 11940 18776 11946 18788
rect 12980 18785 12992 18788
rect 13026 18816 13038 18819
rect 13814 18816 13820 18828
rect 13026 18788 13820 18816
rect 13026 18785 13038 18788
rect 12980 18779 13038 18785
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 15654 18816 15660 18828
rect 15615 18788 15660 18816
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 3050 18748 3056 18760
rect 3011 18720 3056 18748
rect 3050 18708 3056 18720
rect 3108 18708 3114 18760
rect 3510 18708 3516 18760
rect 3568 18748 3574 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 3568 18720 4077 18748
rect 3568 18708 3574 18720
rect 4065 18717 4077 18720
rect 4111 18717 4123 18751
rect 4065 18711 4123 18717
rect 7193 18751 7251 18757
rect 7193 18717 7205 18751
rect 7239 18748 7251 18751
rect 7374 18748 7380 18760
rect 7239 18720 7380 18748
rect 7239 18717 7251 18720
rect 7193 18711 7251 18717
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 10226 18748 10232 18760
rect 10187 18720 10232 18748
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 12710 18748 12716 18760
rect 12671 18720 12716 18748
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 2501 18683 2559 18689
rect 2501 18649 2513 18683
rect 2547 18680 2559 18683
rect 2774 18680 2780 18692
rect 2547 18652 2780 18680
rect 2547 18649 2559 18652
rect 2501 18643 2559 18649
rect 2774 18640 2780 18652
rect 2832 18640 2838 18692
rect 9769 18683 9827 18689
rect 9769 18649 9781 18683
rect 9815 18680 9827 18683
rect 9858 18680 9864 18692
rect 9815 18652 9864 18680
rect 9815 18649 9827 18652
rect 9769 18643 9827 18649
rect 9858 18640 9864 18652
rect 9916 18640 9922 18692
rect 2958 18572 2964 18624
rect 3016 18612 3022 18624
rect 4246 18612 4252 18624
rect 3016 18584 4252 18612
rect 3016 18572 3022 18584
rect 4246 18572 4252 18584
rect 4304 18572 4310 18624
rect 6641 18615 6699 18621
rect 6641 18581 6653 18615
rect 6687 18612 6699 18615
rect 6822 18612 6828 18624
rect 6687 18584 6828 18612
rect 6687 18581 6699 18584
rect 6641 18575 6699 18581
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 11330 18572 11336 18624
rect 11388 18612 11394 18624
rect 11701 18615 11759 18621
rect 11701 18612 11713 18615
rect 11388 18584 11713 18612
rect 11388 18572 11394 18584
rect 11701 18581 11713 18584
rect 11747 18581 11759 18615
rect 11701 18575 11759 18581
rect 12529 18615 12587 18621
rect 12529 18581 12541 18615
rect 12575 18612 12587 18615
rect 12894 18612 12900 18624
rect 12575 18584 12900 18612
rect 12575 18581 12587 18584
rect 12529 18575 12587 18581
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 13078 18572 13084 18624
rect 13136 18612 13142 18624
rect 14093 18615 14151 18621
rect 14093 18612 14105 18615
rect 13136 18584 14105 18612
rect 13136 18572 13142 18584
rect 14093 18581 14105 18584
rect 14139 18581 14151 18615
rect 15378 18612 15384 18624
rect 15339 18584 15384 18612
rect 14093 18575 14151 18581
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2041 18411 2099 18417
rect 2041 18377 2053 18411
rect 2087 18408 2099 18411
rect 3050 18408 3056 18420
rect 2087 18380 3056 18408
rect 2087 18377 2099 18380
rect 2041 18371 2099 18377
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 3510 18408 3516 18420
rect 3160 18380 3516 18408
rect 2961 18343 3019 18349
rect 2961 18309 2973 18343
rect 3007 18340 3019 18343
rect 3160 18340 3188 18380
rect 3510 18368 3516 18380
rect 3568 18368 3574 18420
rect 4338 18368 4344 18420
rect 4396 18408 4402 18420
rect 4525 18411 4583 18417
rect 4525 18408 4537 18411
rect 4396 18380 4537 18408
rect 4396 18368 4402 18380
rect 4525 18377 4537 18380
rect 4571 18408 4583 18411
rect 5077 18411 5135 18417
rect 5077 18408 5089 18411
rect 4571 18380 5089 18408
rect 4571 18377 4583 18380
rect 4525 18371 4583 18377
rect 5077 18377 5089 18380
rect 5123 18377 5135 18411
rect 5077 18371 5135 18377
rect 7098 18368 7104 18420
rect 7156 18408 7162 18420
rect 8205 18411 8263 18417
rect 8205 18408 8217 18411
rect 7156 18380 8217 18408
rect 7156 18368 7162 18380
rect 8205 18377 8217 18380
rect 8251 18377 8263 18411
rect 11882 18408 11888 18420
rect 11843 18380 11888 18408
rect 8205 18371 8263 18377
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 12526 18408 12532 18420
rect 12487 18380 12532 18408
rect 12526 18368 12532 18380
rect 12584 18368 12590 18420
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 13446 18408 13452 18420
rect 12768 18380 13452 18408
rect 12768 18368 12774 18380
rect 13446 18368 13452 18380
rect 13504 18368 13510 18420
rect 13906 18368 13912 18420
rect 13964 18408 13970 18420
rect 14093 18411 14151 18417
rect 14093 18408 14105 18411
rect 13964 18380 14105 18408
rect 13964 18368 13970 18380
rect 14093 18377 14105 18380
rect 14139 18377 14151 18411
rect 14093 18371 14151 18377
rect 14734 18368 14740 18420
rect 14792 18408 14798 18420
rect 15013 18411 15071 18417
rect 15013 18408 15025 18411
rect 14792 18380 15025 18408
rect 14792 18368 14798 18380
rect 15013 18377 15025 18380
rect 15059 18377 15071 18411
rect 15013 18371 15071 18377
rect 15746 18368 15752 18420
rect 15804 18408 15810 18420
rect 16945 18411 17003 18417
rect 16945 18408 16957 18411
rect 15804 18380 16957 18408
rect 15804 18368 15810 18380
rect 16945 18377 16957 18380
rect 16991 18377 17003 18411
rect 16945 18371 17003 18377
rect 3007 18312 3188 18340
rect 3007 18309 3019 18312
rect 2961 18303 3019 18309
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18272 2191 18275
rect 2314 18272 2320 18284
rect 2179 18244 2320 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 2314 18232 2320 18244
rect 2372 18232 2378 18284
rect 3160 18281 3188 18312
rect 4154 18300 4160 18352
rect 4212 18340 4218 18352
rect 6362 18340 6368 18352
rect 4212 18312 6368 18340
rect 4212 18300 4218 18312
rect 6362 18300 6368 18312
rect 6420 18300 6426 18352
rect 6917 18343 6975 18349
rect 6917 18309 6929 18343
rect 6963 18340 6975 18343
rect 7926 18340 7932 18352
rect 6963 18312 7932 18340
rect 6963 18309 6975 18312
rect 6917 18303 6975 18309
rect 7926 18300 7932 18312
rect 7984 18300 7990 18352
rect 9309 18343 9367 18349
rect 9309 18309 9321 18343
rect 9355 18340 9367 18343
rect 9582 18340 9588 18352
rect 9355 18312 9588 18340
rect 9355 18309 9367 18312
rect 9309 18303 9367 18309
rect 9582 18300 9588 18312
rect 9640 18300 9646 18352
rect 10870 18340 10876 18352
rect 10831 18312 10876 18340
rect 10870 18300 10876 18312
rect 10928 18300 10934 18352
rect 15657 18343 15715 18349
rect 15657 18309 15669 18343
rect 15703 18309 15715 18343
rect 15657 18303 15715 18309
rect 3145 18275 3203 18281
rect 3145 18241 3157 18275
rect 3191 18272 3203 18275
rect 3191 18244 3225 18272
rect 3191 18241 3203 18244
rect 3145 18235 3203 18241
rect 2685 18207 2743 18213
rect 2685 18173 2697 18207
rect 2731 18204 2743 18207
rect 3050 18204 3056 18216
rect 2731 18176 3056 18204
rect 2731 18173 2743 18176
rect 2685 18167 2743 18173
rect 3050 18164 3056 18176
rect 3108 18204 3114 18216
rect 3412 18207 3470 18213
rect 3412 18204 3424 18207
rect 3108 18176 3424 18204
rect 3108 18164 3114 18176
rect 3412 18173 3424 18176
rect 3458 18204 3470 18207
rect 4172 18204 4200 18300
rect 6273 18275 6331 18281
rect 6273 18241 6285 18275
rect 6319 18272 6331 18275
rect 7374 18272 7380 18284
rect 6319 18244 7380 18272
rect 6319 18241 6331 18244
rect 6273 18235 6331 18241
rect 7374 18232 7380 18244
rect 7432 18272 7438 18284
rect 7469 18275 7527 18281
rect 7469 18272 7481 18275
rect 7432 18244 7481 18272
rect 7432 18232 7438 18244
rect 7469 18241 7481 18244
rect 7515 18272 7527 18275
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 7515 18244 7849 18272
rect 7515 18241 7527 18244
rect 7469 18235 7527 18241
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 9214 18232 9220 18284
rect 9272 18272 9278 18284
rect 9677 18275 9735 18281
rect 9677 18272 9689 18275
rect 9272 18244 9689 18272
rect 9272 18232 9278 18244
rect 9677 18241 9689 18244
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 10962 18232 10968 18284
rect 11020 18272 11026 18284
rect 11330 18272 11336 18284
rect 11020 18244 11336 18272
rect 11020 18232 11026 18244
rect 11330 18232 11336 18244
rect 11388 18232 11394 18284
rect 13078 18272 13084 18284
rect 13039 18244 13084 18272
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 14550 18272 14556 18284
rect 14463 18244 14556 18272
rect 14550 18232 14556 18244
rect 14608 18272 14614 18284
rect 15378 18272 15384 18284
rect 14608 18244 15384 18272
rect 14608 18232 14614 18244
rect 15378 18232 15384 18244
rect 15436 18232 15442 18284
rect 3458 18176 4200 18204
rect 3458 18173 3470 18176
rect 3412 18167 3470 18173
rect 5442 18164 5448 18216
rect 5500 18204 5506 18216
rect 5629 18207 5687 18213
rect 5629 18204 5641 18207
rect 5500 18176 5641 18204
rect 5500 18164 5506 18176
rect 5629 18173 5641 18176
rect 5675 18204 5687 18207
rect 5675 18176 7420 18204
rect 5675 18173 5687 18176
rect 5629 18167 5687 18173
rect 1673 18139 1731 18145
rect 1673 18105 1685 18139
rect 1719 18136 1731 18139
rect 2498 18136 2504 18148
rect 1719 18108 2504 18136
rect 1719 18105 1731 18108
rect 1673 18099 1731 18105
rect 2498 18096 2504 18108
rect 2556 18096 2562 18148
rect 7392 18145 7420 18176
rect 8110 18164 8116 18216
rect 8168 18204 8174 18216
rect 8757 18207 8815 18213
rect 8757 18204 8769 18207
rect 8168 18176 8769 18204
rect 8168 18164 8174 18176
rect 8757 18173 8769 18176
rect 8803 18204 8815 18207
rect 9861 18207 9919 18213
rect 9861 18204 9873 18207
rect 8803 18176 9873 18204
rect 8803 18173 8815 18176
rect 8757 18167 8815 18173
rect 9861 18173 9873 18176
rect 9907 18173 9919 18207
rect 14090 18204 14096 18216
rect 9861 18167 9919 18173
rect 12820 18176 14096 18204
rect 5721 18139 5779 18145
rect 5721 18105 5733 18139
rect 5767 18136 5779 18139
rect 6641 18139 6699 18145
rect 6641 18136 6653 18139
rect 5767 18108 6653 18136
rect 5767 18105 5779 18108
rect 5721 18099 5779 18105
rect 6641 18105 6653 18108
rect 6687 18136 6699 18139
rect 7193 18139 7251 18145
rect 7193 18136 7205 18139
rect 6687 18108 7205 18136
rect 6687 18105 6699 18108
rect 6641 18099 6699 18105
rect 7193 18105 7205 18108
rect 7239 18105 7251 18139
rect 7193 18099 7251 18105
rect 7377 18139 7435 18145
rect 7377 18105 7389 18139
rect 7423 18105 7435 18139
rect 7377 18099 7435 18105
rect 9674 18096 9680 18148
rect 9732 18136 9738 18148
rect 10226 18136 10232 18148
rect 9732 18108 10232 18136
rect 9732 18096 9738 18108
rect 10226 18096 10232 18108
rect 10284 18096 10290 18148
rect 10689 18139 10747 18145
rect 10689 18105 10701 18139
rect 10735 18136 10747 18139
rect 11425 18139 11483 18145
rect 11425 18136 11437 18139
rect 10735 18108 11437 18136
rect 10735 18105 10747 18108
rect 10689 18099 10747 18105
rect 11425 18105 11437 18108
rect 11471 18136 11483 18139
rect 12250 18136 12256 18148
rect 11471 18108 12256 18136
rect 11471 18105 11483 18108
rect 11425 18099 11483 18105
rect 12250 18096 12256 18108
rect 12308 18096 12314 18148
rect 12820 18145 12848 18176
rect 14090 18164 14096 18176
rect 14148 18164 14154 18216
rect 15672 18204 15700 18303
rect 15930 18232 15936 18284
rect 15988 18272 15994 18284
rect 16209 18275 16267 18281
rect 16209 18272 16221 18275
rect 15988 18244 16221 18272
rect 15988 18232 15994 18244
rect 16209 18241 16221 18244
rect 16255 18241 16267 18275
rect 21542 18272 21548 18284
rect 21503 18244 21548 18272
rect 16209 18235 16267 18241
rect 21542 18232 21548 18244
rect 21600 18232 21606 18284
rect 16577 18207 16635 18213
rect 16577 18204 16589 18207
rect 14568 18176 15700 18204
rect 16132 18176 16589 18204
rect 12805 18139 12863 18145
rect 12805 18136 12817 18139
rect 12360 18108 12817 18136
rect 2682 18028 2688 18080
rect 2740 18068 2746 18080
rect 9033 18071 9091 18077
rect 9033 18068 9045 18071
rect 2740 18040 9045 18068
rect 2740 18028 2746 18040
rect 9033 18037 9045 18040
rect 9079 18068 9091 18071
rect 9766 18068 9772 18080
rect 9079 18040 9772 18068
rect 9079 18037 9091 18040
rect 9033 18031 9091 18037
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 11330 18068 11336 18080
rect 11291 18040 11336 18068
rect 11330 18028 11336 18040
rect 11388 18028 11394 18080
rect 12066 18028 12072 18080
rect 12124 18068 12130 18080
rect 12161 18071 12219 18077
rect 12161 18068 12173 18071
rect 12124 18040 12173 18068
rect 12124 18028 12130 18040
rect 12161 18037 12173 18040
rect 12207 18068 12219 18071
rect 12360 18068 12388 18108
rect 12805 18105 12817 18108
rect 12851 18105 12863 18139
rect 12805 18099 12863 18105
rect 12894 18096 12900 18148
rect 12952 18136 12958 18148
rect 12952 18108 13952 18136
rect 12952 18096 12958 18108
rect 12986 18068 12992 18080
rect 12207 18040 12388 18068
rect 12947 18040 12992 18068
rect 12207 18037 12219 18040
rect 12161 18031 12219 18037
rect 12986 18028 12992 18040
rect 13044 18028 13050 18080
rect 13446 18068 13452 18080
rect 13407 18040 13452 18068
rect 13446 18028 13452 18040
rect 13504 18028 13510 18080
rect 13924 18077 13952 18108
rect 14182 18096 14188 18148
rect 14240 18136 14246 18148
rect 14568 18145 14596 18176
rect 16132 18148 16160 18176
rect 16577 18173 16589 18176
rect 16623 18173 16635 18207
rect 21266 18204 21272 18216
rect 21227 18176 21272 18204
rect 16577 18167 16635 18173
rect 21266 18164 21272 18176
rect 21324 18204 21330 18216
rect 22005 18207 22063 18213
rect 22005 18204 22017 18207
rect 21324 18176 22017 18204
rect 21324 18164 21330 18176
rect 22005 18173 22017 18176
rect 22051 18173 22063 18207
rect 22005 18167 22063 18173
rect 14553 18139 14611 18145
rect 14553 18136 14565 18139
rect 14240 18108 14565 18136
rect 14240 18096 14246 18108
rect 14553 18105 14565 18108
rect 14599 18105 14611 18139
rect 14553 18099 14611 18105
rect 14645 18139 14703 18145
rect 14645 18105 14657 18139
rect 14691 18105 14703 18139
rect 15378 18136 15384 18148
rect 15339 18108 15384 18136
rect 14645 18099 14703 18105
rect 13909 18071 13967 18077
rect 13909 18037 13921 18071
rect 13955 18068 13967 18071
rect 14660 18068 14688 18099
rect 15378 18096 15384 18108
rect 15436 18136 15442 18148
rect 15933 18139 15991 18145
rect 15933 18136 15945 18139
rect 15436 18108 15945 18136
rect 15436 18096 15442 18108
rect 15933 18105 15945 18108
rect 15979 18105 15991 18139
rect 16114 18136 16120 18148
rect 16075 18108 16120 18136
rect 15933 18099 15991 18105
rect 16114 18096 16120 18108
rect 16172 18096 16178 18148
rect 13955 18040 14688 18068
rect 13955 18037 13967 18040
rect 13909 18031 13967 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2317 17867 2375 17873
rect 2317 17833 2329 17867
rect 2363 17864 2375 17867
rect 2406 17864 2412 17876
rect 2363 17836 2412 17864
rect 2363 17833 2375 17836
rect 2317 17827 2375 17833
rect 2406 17824 2412 17836
rect 2464 17824 2470 17876
rect 3510 17824 3516 17876
rect 3568 17864 3574 17876
rect 4249 17867 4307 17873
rect 4249 17864 4261 17867
rect 3568 17836 4261 17864
rect 3568 17824 3574 17836
rect 4249 17833 4261 17836
rect 4295 17864 4307 17867
rect 4430 17864 4436 17876
rect 4295 17836 4436 17864
rect 4295 17833 4307 17836
rect 4249 17827 4307 17833
rect 4430 17824 4436 17836
rect 4488 17824 4494 17876
rect 6457 17867 6515 17873
rect 6457 17833 6469 17867
rect 6503 17833 6515 17867
rect 7374 17864 7380 17876
rect 7335 17836 7380 17864
rect 6457 17827 6515 17833
rect 2774 17756 2780 17808
rect 2832 17796 2838 17808
rect 2961 17799 3019 17805
rect 2961 17796 2973 17799
rect 2832 17768 2973 17796
rect 2832 17756 2838 17768
rect 2961 17765 2973 17768
rect 3007 17765 3019 17799
rect 2961 17759 3019 17765
rect 3050 17756 3056 17808
rect 3108 17796 3114 17808
rect 5350 17805 5356 17808
rect 5344 17796 5356 17805
rect 3108 17768 3153 17796
rect 5311 17768 5356 17796
rect 3108 17756 3114 17768
rect 5344 17759 5356 17768
rect 5350 17756 5356 17759
rect 5408 17756 5414 17808
rect 6270 17756 6276 17808
rect 6328 17796 6334 17808
rect 6472 17796 6500 17827
rect 7374 17824 7380 17836
rect 7432 17824 7438 17876
rect 8573 17867 8631 17873
rect 8573 17864 8585 17867
rect 7944 17836 8585 17864
rect 7944 17808 7972 17836
rect 8573 17833 8585 17836
rect 8619 17833 8631 17867
rect 9214 17864 9220 17876
rect 9175 17836 9220 17864
rect 8573 17827 8631 17833
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 10042 17824 10048 17876
rect 10100 17864 10106 17876
rect 10321 17867 10379 17873
rect 10321 17864 10333 17867
rect 10100 17836 10333 17864
rect 10100 17824 10106 17836
rect 10321 17833 10333 17836
rect 10367 17833 10379 17867
rect 10321 17827 10379 17833
rect 10771 17867 10829 17873
rect 10771 17833 10783 17867
rect 10817 17864 10829 17867
rect 11330 17864 11336 17876
rect 10817 17836 11336 17864
rect 10817 17833 10829 17836
rect 10771 17827 10829 17833
rect 11330 17824 11336 17836
rect 11388 17864 11394 17876
rect 11701 17867 11759 17873
rect 11701 17864 11713 17867
rect 11388 17836 11713 17864
rect 11388 17824 11394 17836
rect 11701 17833 11713 17836
rect 11747 17833 11759 17867
rect 11701 17827 11759 17833
rect 11882 17824 11888 17876
rect 11940 17864 11946 17876
rect 12069 17867 12127 17873
rect 12069 17864 12081 17867
rect 11940 17836 12081 17864
rect 11940 17824 11946 17836
rect 12069 17833 12081 17836
rect 12115 17833 12127 17867
rect 12069 17827 12127 17833
rect 12250 17824 12256 17876
rect 12308 17864 12314 17876
rect 13354 17864 13360 17876
rect 12308 17836 13360 17864
rect 12308 17824 12314 17836
rect 13354 17824 13360 17836
rect 13412 17864 13418 17876
rect 13725 17867 13783 17873
rect 13725 17864 13737 17867
rect 13412 17836 13737 17864
rect 13412 17824 13418 17836
rect 13725 17833 13737 17836
rect 13771 17833 13783 17867
rect 14182 17864 14188 17876
rect 14143 17836 14188 17864
rect 13725 17827 13783 17833
rect 14182 17824 14188 17836
rect 14240 17824 14246 17876
rect 14550 17864 14556 17876
rect 14511 17836 14556 17864
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 15105 17867 15163 17873
rect 15105 17833 15117 17867
rect 15151 17864 15163 17867
rect 15151 17836 15976 17864
rect 15151 17833 15163 17836
rect 15105 17827 15163 17833
rect 15948 17808 15976 17836
rect 7101 17799 7159 17805
rect 7101 17796 7113 17799
rect 6328 17768 7113 17796
rect 6328 17756 6334 17768
rect 7101 17765 7113 17768
rect 7147 17796 7159 17799
rect 7558 17796 7564 17808
rect 7147 17768 7564 17796
rect 7147 17765 7159 17768
rect 7101 17759 7159 17765
rect 7558 17756 7564 17768
rect 7616 17756 7622 17808
rect 7926 17796 7932 17808
rect 7887 17768 7932 17796
rect 7926 17756 7932 17768
rect 7984 17756 7990 17808
rect 8113 17799 8171 17805
rect 8113 17765 8125 17799
rect 8159 17765 8171 17799
rect 8113 17759 8171 17765
rect 6822 17688 6828 17740
rect 6880 17728 6886 17740
rect 8128 17728 8156 17759
rect 10226 17756 10232 17808
rect 10284 17796 10290 17808
rect 11241 17799 11299 17805
rect 11241 17796 11253 17799
rect 10284 17768 11253 17796
rect 10284 17756 10290 17768
rect 11241 17765 11253 17768
rect 11287 17796 11299 17799
rect 12434 17796 12440 17808
rect 11287 17768 12440 17796
rect 11287 17765 11299 17768
rect 11241 17759 11299 17765
rect 12434 17756 12440 17768
rect 12492 17756 12498 17808
rect 12529 17799 12587 17805
rect 12529 17765 12541 17799
rect 12575 17796 12587 17799
rect 12986 17796 12992 17808
rect 12575 17768 12992 17796
rect 12575 17765 12587 17768
rect 12529 17759 12587 17765
rect 12986 17756 12992 17768
rect 13044 17756 13050 17808
rect 13262 17796 13268 17808
rect 13223 17768 13268 17796
rect 13262 17756 13268 17768
rect 13320 17756 13326 17808
rect 15838 17796 15844 17808
rect 15799 17768 15844 17796
rect 15838 17756 15844 17768
rect 15896 17756 15902 17808
rect 15930 17756 15936 17808
rect 15988 17796 15994 17808
rect 16301 17799 16359 17805
rect 16301 17796 16313 17799
rect 15988 17768 16313 17796
rect 15988 17756 15994 17768
rect 16301 17765 16313 17768
rect 16347 17796 16359 17799
rect 16390 17796 16396 17808
rect 16347 17768 16396 17796
rect 16347 17765 16359 17768
rect 16301 17759 16359 17765
rect 16390 17756 16396 17768
rect 16448 17756 16454 17808
rect 9122 17728 9128 17740
rect 6880 17700 9128 17728
rect 6880 17688 6886 17700
rect 9122 17688 9128 17700
rect 9180 17688 9186 17740
rect 13078 17688 13084 17740
rect 13136 17728 13142 17740
rect 13357 17731 13415 17737
rect 13357 17728 13369 17731
rect 13136 17700 13369 17728
rect 13136 17688 13142 17700
rect 13357 17697 13369 17700
rect 13403 17697 13415 17731
rect 13357 17691 13415 17697
rect 15378 17688 15384 17740
rect 15436 17728 15442 17740
rect 15657 17731 15715 17737
rect 15657 17728 15669 17731
rect 15436 17700 15669 17728
rect 15436 17688 15442 17700
rect 15657 17697 15669 17700
rect 15703 17728 15715 17731
rect 15746 17728 15752 17740
rect 15703 17700 15752 17728
rect 15703 17697 15715 17700
rect 15657 17691 15715 17697
rect 15746 17688 15752 17700
rect 15804 17688 15810 17740
rect 2866 17660 2872 17672
rect 2827 17632 2872 17660
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 4430 17620 4436 17672
rect 4488 17660 4494 17672
rect 5077 17663 5135 17669
rect 5077 17660 5089 17663
rect 4488 17632 5089 17660
rect 4488 17620 4494 17632
rect 5077 17629 5089 17632
rect 5123 17629 5135 17663
rect 8202 17660 8208 17672
rect 8163 17632 8208 17660
rect 5077 17623 5135 17629
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 11238 17660 11244 17672
rect 11199 17632 11244 17660
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 11333 17663 11391 17669
rect 11333 17629 11345 17663
rect 11379 17660 11391 17663
rect 11422 17660 11428 17672
rect 11379 17632 11428 17660
rect 11379 17629 11391 17632
rect 11333 17623 11391 17629
rect 11422 17620 11428 17632
rect 11480 17620 11486 17672
rect 13170 17660 13176 17672
rect 13131 17632 13176 17660
rect 13170 17620 13176 17632
rect 13228 17620 13234 17672
rect 2498 17592 2504 17604
rect 2459 17564 2504 17592
rect 2498 17552 2504 17564
rect 2556 17552 2562 17604
rect 7650 17592 7656 17604
rect 7611 17564 7656 17592
rect 7650 17552 7656 17564
rect 7708 17552 7714 17604
rect 15286 17552 15292 17604
rect 15344 17592 15350 17604
rect 15381 17595 15439 17601
rect 15381 17592 15393 17595
rect 15344 17564 15393 17592
rect 15344 17552 15350 17564
rect 15381 17561 15393 17564
rect 15427 17561 15439 17595
rect 15381 17555 15439 17561
rect 9953 17527 10011 17533
rect 9953 17493 9965 17527
rect 9999 17524 10011 17527
rect 10686 17524 10692 17536
rect 9999 17496 10692 17524
rect 9999 17493 10011 17496
rect 9953 17487 10011 17493
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 12802 17524 12808 17536
rect 12763 17496 12808 17524
rect 12802 17484 12808 17496
rect 12860 17484 12866 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2501 17323 2559 17329
rect 2501 17289 2513 17323
rect 2547 17320 2559 17323
rect 2774 17320 2780 17332
rect 2547 17292 2780 17320
rect 2547 17289 2559 17292
rect 2501 17283 2559 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 2866 17280 2872 17332
rect 2924 17320 2930 17332
rect 2924 17292 2969 17320
rect 2924 17280 2930 17292
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 3145 17323 3203 17329
rect 3145 17320 3157 17323
rect 3108 17292 3157 17320
rect 3108 17280 3114 17292
rect 3145 17289 3157 17292
rect 3191 17289 3203 17323
rect 3145 17283 3203 17289
rect 3878 17280 3884 17332
rect 3936 17320 3942 17332
rect 4893 17323 4951 17329
rect 4893 17320 4905 17323
rect 3936 17292 4905 17320
rect 3936 17280 3942 17292
rect 4893 17289 4905 17292
rect 4939 17320 4951 17323
rect 4985 17323 5043 17329
rect 4985 17320 4997 17323
rect 4939 17292 4997 17320
rect 4939 17289 4951 17292
rect 4893 17283 4951 17289
rect 4985 17289 4997 17292
rect 5031 17289 5043 17323
rect 4985 17283 5043 17289
rect 5261 17323 5319 17329
rect 5261 17289 5273 17323
rect 5307 17320 5319 17323
rect 5442 17320 5448 17332
rect 5307 17292 5448 17320
rect 5307 17289 5319 17292
rect 5261 17283 5319 17289
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 6270 17320 6276 17332
rect 6231 17292 6276 17320
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 8202 17280 8208 17332
rect 8260 17320 8266 17332
rect 8757 17323 8815 17329
rect 8757 17320 8769 17323
rect 8260 17292 8769 17320
rect 8260 17280 8266 17292
rect 8757 17289 8769 17292
rect 8803 17289 8815 17323
rect 9122 17320 9128 17332
rect 9083 17292 9128 17320
rect 8757 17283 8815 17289
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 10873 17323 10931 17329
rect 10873 17289 10885 17323
rect 10919 17320 10931 17323
rect 10962 17320 10968 17332
rect 10919 17292 10968 17320
rect 10919 17289 10931 17292
rect 10873 17283 10931 17289
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 12253 17323 12311 17329
rect 12253 17289 12265 17323
rect 12299 17320 12311 17323
rect 13078 17320 13084 17332
rect 12299 17292 13084 17320
rect 12299 17289 12311 17292
rect 12253 17283 12311 17289
rect 13078 17280 13084 17292
rect 13136 17320 13142 17332
rect 14461 17323 14519 17329
rect 14461 17320 14473 17323
rect 13136 17292 14473 17320
rect 13136 17280 13142 17292
rect 14461 17289 14473 17292
rect 14507 17289 14519 17323
rect 14461 17283 14519 17289
rect 15838 17280 15844 17332
rect 15896 17320 15902 17332
rect 16025 17323 16083 17329
rect 16025 17320 16037 17323
rect 15896 17292 16037 17320
rect 15896 17280 15902 17292
rect 16025 17289 16037 17292
rect 16071 17289 16083 17323
rect 16390 17320 16396 17332
rect 16351 17292 16396 17320
rect 16025 17283 16083 17289
rect 16390 17280 16396 17292
rect 16448 17280 16454 17332
rect 4341 17255 4399 17261
rect 4341 17221 4353 17255
rect 4387 17252 4399 17255
rect 5350 17252 5356 17264
rect 4387 17224 5356 17252
rect 4387 17221 4399 17224
rect 4341 17215 4399 17221
rect 5350 17212 5356 17224
rect 5408 17212 5414 17264
rect 4430 17144 4436 17196
rect 4488 17184 4494 17196
rect 4617 17187 4675 17193
rect 4617 17184 4629 17187
rect 4488 17156 4629 17184
rect 4488 17144 4494 17156
rect 4617 17153 4629 17156
rect 4663 17184 4675 17187
rect 5442 17184 5448 17196
rect 4663 17156 5448 17184
rect 4663 17153 4675 17156
rect 4617 17147 4675 17153
rect 5442 17144 5448 17156
rect 5500 17184 5506 17196
rect 5813 17187 5871 17193
rect 5500 17156 5672 17184
rect 5500 17144 5506 17156
rect 4893 17119 4951 17125
rect 4893 17085 4905 17119
rect 4939 17116 4951 17119
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 4939 17088 5549 17116
rect 4939 17085 4951 17088
rect 4893 17079 4951 17085
rect 5537 17085 5549 17088
rect 5583 17085 5595 17119
rect 5644 17116 5672 17156
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 6288 17184 6316 17280
rect 10689 17255 10747 17261
rect 10689 17221 10701 17255
rect 10735 17252 10747 17255
rect 11238 17252 11244 17264
rect 10735 17224 11244 17252
rect 10735 17221 10747 17224
rect 10689 17215 10747 17221
rect 11238 17212 11244 17224
rect 11296 17212 11302 17264
rect 5859 17156 6960 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 6549 17119 6607 17125
rect 6549 17116 6561 17119
rect 5644 17088 6561 17116
rect 5537 17079 5595 17085
rect 6549 17085 6561 17088
rect 6595 17116 6607 17119
rect 6822 17116 6828 17128
rect 6595 17088 6828 17116
rect 6595 17085 6607 17088
rect 6549 17079 6607 17085
rect 5552 17048 5580 17079
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 6932 17116 6960 17156
rect 9766 17144 9772 17196
rect 9824 17184 9830 17196
rect 10134 17184 10140 17196
rect 9824 17156 10140 17184
rect 9824 17144 9830 17156
rect 10134 17144 10140 17156
rect 10192 17144 10198 17196
rect 7098 17125 7104 17128
rect 7081 17119 7104 17125
rect 7081 17116 7093 17119
rect 6932 17088 7093 17116
rect 7081 17085 7093 17088
rect 7156 17116 7162 17128
rect 13354 17125 13360 17128
rect 9953 17119 10011 17125
rect 7156 17088 7229 17116
rect 7081 17079 7104 17085
rect 7098 17076 7104 17079
rect 7156 17076 7162 17088
rect 9953 17085 9965 17119
rect 9999 17116 10011 17119
rect 11793 17119 11851 17125
rect 11793 17116 11805 17119
rect 9999 17088 11805 17116
rect 9999 17085 10011 17088
rect 9953 17079 10011 17085
rect 11440 17060 11468 17088
rect 11793 17085 11805 17088
rect 11839 17085 11851 17119
rect 13081 17119 13139 17125
rect 13081 17116 13093 17119
rect 11793 17079 11851 17085
rect 12912 17088 13093 17116
rect 11146 17048 11152 17060
rect 5552 17020 6868 17048
rect 11107 17020 11152 17048
rect 1673 16983 1731 16989
rect 1673 16949 1685 16983
rect 1719 16980 1731 16983
rect 1854 16980 1860 16992
rect 1719 16952 1860 16980
rect 1719 16949 1731 16952
rect 1673 16943 1731 16949
rect 1854 16940 1860 16952
rect 1912 16940 1918 16992
rect 5718 16980 5724 16992
rect 5679 16952 5724 16980
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 6840 16980 6868 17020
rect 11146 17008 11152 17020
rect 11204 17008 11210 17060
rect 11422 17048 11428 17060
rect 11383 17020 11428 17048
rect 11422 17008 11428 17020
rect 11480 17008 11486 17060
rect 12912 17048 12940 17088
rect 13081 17085 13093 17088
rect 13127 17085 13139 17119
rect 13348 17116 13360 17125
rect 13315 17088 13360 17116
rect 13081 17079 13139 17085
rect 13348 17079 13360 17088
rect 13354 17076 13360 17079
rect 13412 17076 13418 17128
rect 13446 17048 13452 17060
rect 12912 17020 13452 17048
rect 12912 16992 12940 17020
rect 13446 17008 13452 17020
rect 13504 17008 13510 17060
rect 7006 16980 7012 16992
rect 6840 16952 7012 16980
rect 7006 16940 7012 16952
rect 7064 16940 7070 16992
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 8205 16983 8263 16989
rect 8205 16980 8217 16983
rect 7432 16952 8217 16980
rect 7432 16940 7438 16952
rect 8205 16949 8217 16952
rect 8251 16949 8263 16983
rect 8205 16943 8263 16949
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 10192 16952 10241 16980
rect 10192 16940 10198 16952
rect 10229 16949 10241 16952
rect 10275 16949 10287 16983
rect 10229 16943 10287 16949
rect 10870 16940 10876 16992
rect 10928 16980 10934 16992
rect 11333 16983 11391 16989
rect 11333 16980 11345 16983
rect 10928 16952 11345 16980
rect 10928 16940 10934 16952
rect 11333 16949 11345 16952
rect 11379 16980 11391 16983
rect 11974 16980 11980 16992
rect 11379 16952 11980 16980
rect 11379 16949 11391 16952
rect 11333 16943 11391 16949
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 12894 16980 12900 16992
rect 12855 16952 12900 16980
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 15286 16980 15292 16992
rect 15247 16952 15292 16980
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 15565 16983 15623 16989
rect 15565 16949 15577 16983
rect 15611 16980 15623 16983
rect 15838 16980 15844 16992
rect 15611 16952 15844 16980
rect 15611 16949 15623 16952
rect 15565 16943 15623 16949
rect 15838 16940 15844 16952
rect 15896 16940 15902 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 4154 16736 4160 16788
rect 4212 16776 4218 16788
rect 4982 16776 4988 16788
rect 4212 16748 4988 16776
rect 4212 16736 4218 16748
rect 4982 16736 4988 16748
rect 5040 16776 5046 16788
rect 5169 16779 5227 16785
rect 5169 16776 5181 16779
rect 5040 16748 5181 16776
rect 5040 16736 5046 16748
rect 5169 16745 5181 16748
rect 5215 16776 5227 16779
rect 5718 16776 5724 16788
rect 5215 16748 5724 16776
rect 5215 16745 5227 16748
rect 5169 16739 5227 16745
rect 5718 16736 5724 16748
rect 5776 16776 5782 16788
rect 5776 16748 5948 16776
rect 5776 16736 5782 16748
rect 5920 16717 5948 16748
rect 8202 16736 8208 16788
rect 8260 16776 8266 16788
rect 8481 16779 8539 16785
rect 8481 16776 8493 16779
rect 8260 16748 8493 16776
rect 8260 16736 8266 16748
rect 8481 16745 8493 16748
rect 8527 16776 8539 16779
rect 8754 16776 8760 16788
rect 8527 16748 8760 16776
rect 8527 16745 8539 16748
rect 8481 16739 8539 16745
rect 8754 16736 8760 16748
rect 8812 16736 8818 16788
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10870 16776 10876 16788
rect 9916 16748 10364 16776
rect 10831 16748 10876 16776
rect 9916 16736 9922 16748
rect 5905 16711 5963 16717
rect 5905 16677 5917 16711
rect 5951 16677 5963 16711
rect 5905 16671 5963 16677
rect 6089 16711 6147 16717
rect 6089 16677 6101 16711
rect 6135 16708 6147 16711
rect 6178 16708 6184 16720
rect 6135 16680 6184 16708
rect 6135 16677 6147 16680
rect 6089 16671 6147 16677
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 7374 16717 7380 16720
rect 7368 16708 7380 16717
rect 7335 16680 7380 16708
rect 7368 16671 7380 16680
rect 7374 16668 7380 16671
rect 7432 16668 7438 16720
rect 10042 16668 10048 16720
rect 10100 16708 10106 16720
rect 10336 16717 10364 16748
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 11146 16776 11152 16788
rect 11107 16748 11152 16776
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 12434 16736 12440 16788
rect 12492 16776 12498 16788
rect 13265 16779 13323 16785
rect 13265 16776 13277 16779
rect 12492 16748 13277 16776
rect 12492 16736 12498 16748
rect 13265 16745 13277 16748
rect 13311 16776 13323 16779
rect 13354 16776 13360 16788
rect 13311 16748 13360 16776
rect 13311 16745 13323 16748
rect 13265 16739 13323 16745
rect 13354 16736 13360 16748
rect 13412 16736 13418 16788
rect 15470 16736 15476 16788
rect 15528 16776 15534 16788
rect 15841 16779 15899 16785
rect 15841 16776 15853 16779
rect 15528 16748 15853 16776
rect 15528 16736 15534 16748
rect 15841 16745 15853 16748
rect 15887 16745 15899 16779
rect 15841 16739 15899 16745
rect 10229 16711 10287 16717
rect 10229 16708 10241 16711
rect 10100 16680 10241 16708
rect 10100 16668 10106 16680
rect 10229 16677 10241 16680
rect 10275 16677 10287 16711
rect 10229 16671 10287 16677
rect 10321 16711 10379 16717
rect 10321 16677 10333 16711
rect 10367 16677 10379 16711
rect 10321 16671 10379 16677
rect 11422 16668 11428 16720
rect 11480 16708 11486 16720
rect 12130 16711 12188 16717
rect 12130 16708 12142 16711
rect 11480 16680 12142 16708
rect 11480 16668 11486 16680
rect 12130 16677 12142 16680
rect 12176 16708 12188 16711
rect 12710 16708 12716 16720
rect 12176 16680 12716 16708
rect 12176 16677 12188 16680
rect 12130 16671 12188 16677
rect 12710 16668 12716 16680
rect 12768 16668 12774 16720
rect 13078 16668 13084 16720
rect 13136 16708 13142 16720
rect 13909 16711 13967 16717
rect 13909 16708 13921 16711
rect 13136 16680 13921 16708
rect 13136 16668 13142 16680
rect 13909 16677 13921 16680
rect 13955 16708 13967 16711
rect 13998 16708 14004 16720
rect 13955 16680 14004 16708
rect 13955 16677 13967 16680
rect 13909 16671 13967 16677
rect 13998 16668 14004 16680
rect 14056 16668 14062 16720
rect 2406 16640 2412 16652
rect 2367 16612 2412 16640
rect 2406 16600 2412 16612
rect 2464 16600 2470 16652
rect 6822 16600 6828 16652
rect 6880 16640 6886 16652
rect 7101 16643 7159 16649
rect 7101 16640 7113 16643
rect 6880 16612 7113 16640
rect 6880 16600 6886 16612
rect 7101 16609 7113 16612
rect 7147 16609 7159 16643
rect 7101 16603 7159 16609
rect 9751 16643 9809 16649
rect 9751 16609 9763 16643
rect 9797 16640 9809 16643
rect 11054 16640 11060 16652
rect 9797 16612 11060 16640
rect 9797 16609 9809 16612
rect 9751 16603 9809 16609
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 15562 16600 15568 16652
rect 15620 16640 15626 16652
rect 15933 16643 15991 16649
rect 15933 16640 15945 16643
rect 15620 16612 15945 16640
rect 15620 16600 15626 16612
rect 15933 16609 15945 16612
rect 15979 16609 15991 16643
rect 15933 16603 15991 16609
rect 6181 16575 6239 16581
rect 6181 16572 6193 16575
rect 5368 16544 6193 16572
rect 1394 16464 1400 16516
rect 1452 16504 1458 16516
rect 1949 16507 2007 16513
rect 1949 16504 1961 16507
rect 1452 16476 1961 16504
rect 1452 16464 1458 16476
rect 1949 16473 1961 16476
rect 1995 16473 2007 16507
rect 1949 16467 2007 16473
rect 5368 16448 5396 16544
rect 6181 16541 6193 16544
rect 6227 16541 6239 16575
rect 6181 16535 6239 16541
rect 9398 16532 9404 16584
rect 9456 16572 9462 16584
rect 10137 16575 10195 16581
rect 10137 16572 10149 16575
rect 9456 16544 10149 16572
rect 9456 16532 9462 16544
rect 10137 16541 10149 16544
rect 10183 16572 10195 16575
rect 10594 16572 10600 16584
rect 10183 16544 10600 16572
rect 10183 16541 10195 16544
rect 10137 16535 10195 16541
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 11882 16572 11888 16584
rect 11843 16544 11888 16572
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 15838 16572 15844 16584
rect 15799 16544 15844 16572
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 1302 16396 1308 16448
rect 1360 16436 1366 16448
rect 1581 16439 1639 16445
rect 1581 16436 1593 16439
rect 1360 16408 1593 16436
rect 1360 16396 1366 16408
rect 1581 16405 1593 16408
rect 1627 16405 1639 16439
rect 1581 16399 1639 16405
rect 4893 16439 4951 16445
rect 4893 16405 4905 16439
rect 4939 16436 4951 16439
rect 5350 16436 5356 16448
rect 4939 16408 5356 16436
rect 4939 16405 4951 16408
rect 4893 16399 4951 16405
rect 5350 16396 5356 16408
rect 5408 16396 5414 16448
rect 5534 16396 5540 16448
rect 5592 16436 5598 16448
rect 5629 16439 5687 16445
rect 5629 16436 5641 16439
rect 5592 16408 5641 16436
rect 5592 16396 5598 16408
rect 5629 16405 5641 16408
rect 5675 16405 5687 16439
rect 5629 16399 5687 16405
rect 6917 16439 6975 16445
rect 6917 16405 6929 16439
rect 6963 16436 6975 16439
rect 7374 16436 7380 16448
rect 6963 16408 7380 16436
rect 6963 16405 6975 16408
rect 6917 16399 6975 16405
rect 7374 16396 7380 16408
rect 7432 16396 7438 16448
rect 15286 16396 15292 16448
rect 15344 16436 15350 16448
rect 15381 16439 15439 16445
rect 15381 16436 15393 16439
rect 15344 16408 15393 16436
rect 15344 16396 15350 16408
rect 15381 16405 15393 16408
rect 15427 16405 15439 16439
rect 15381 16399 15439 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1857 16235 1915 16241
rect 1857 16201 1869 16235
rect 1903 16232 1915 16235
rect 2222 16232 2228 16244
rect 1903 16204 2228 16232
rect 1903 16201 1915 16204
rect 1857 16195 1915 16201
rect 2222 16192 2228 16204
rect 2280 16192 2286 16244
rect 4982 16232 4988 16244
rect 4943 16204 4988 16232
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 6914 16232 6920 16244
rect 6875 16204 6920 16232
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 10042 16192 10048 16244
rect 10100 16232 10106 16244
rect 11057 16235 11115 16241
rect 11057 16232 11069 16235
rect 10100 16204 11069 16232
rect 10100 16192 10106 16204
rect 11057 16201 11069 16204
rect 11103 16201 11115 16235
rect 11057 16195 11115 16201
rect 13081 16235 13139 16241
rect 13081 16201 13093 16235
rect 13127 16232 13139 16235
rect 13262 16232 13268 16244
rect 13127 16204 13268 16232
rect 13127 16201 13139 16204
rect 13081 16195 13139 16201
rect 13262 16192 13268 16204
rect 13320 16192 13326 16244
rect 15838 16192 15844 16244
rect 15896 16232 15902 16244
rect 16209 16235 16267 16241
rect 16209 16232 16221 16235
rect 15896 16204 16221 16232
rect 15896 16192 15902 16204
rect 16209 16201 16221 16204
rect 16255 16201 16267 16235
rect 16209 16195 16267 16201
rect 2041 16167 2099 16173
rect 2041 16133 2053 16167
rect 2087 16164 2099 16167
rect 2498 16164 2504 16176
rect 2087 16136 2504 16164
rect 2087 16133 2099 16136
rect 2041 16127 2099 16133
rect 2498 16124 2504 16136
rect 2556 16124 2562 16176
rect 5258 16164 5264 16176
rect 5219 16136 5264 16164
rect 5258 16124 5264 16136
rect 5316 16124 5322 16176
rect 6362 16124 6368 16176
rect 6420 16164 6426 16176
rect 6638 16164 6644 16176
rect 6420 16136 6644 16164
rect 6420 16124 6426 16136
rect 6638 16124 6644 16136
rect 6696 16124 6702 16176
rect 6822 16124 6828 16176
rect 6880 16164 6886 16176
rect 7837 16167 7895 16173
rect 7837 16164 7849 16167
rect 6880 16136 7849 16164
rect 6880 16124 6886 16136
rect 7837 16133 7849 16136
rect 7883 16164 7895 16167
rect 8481 16167 8539 16173
rect 8481 16164 8493 16167
rect 7883 16136 8493 16164
rect 7883 16133 7895 16136
rect 7837 16127 7895 16133
rect 8481 16133 8493 16136
rect 8527 16164 8539 16167
rect 10594 16164 10600 16176
rect 8527 16136 8708 16164
rect 10555 16136 10600 16164
rect 8527 16133 8539 16136
rect 8481 16127 8539 16133
rect 8680 16108 8708 16136
rect 10594 16124 10600 16136
rect 10652 16124 10658 16176
rect 13170 16124 13176 16176
rect 13228 16164 13234 16176
rect 13357 16167 13415 16173
rect 13357 16164 13369 16167
rect 13228 16136 13369 16164
rect 13228 16124 13234 16136
rect 13357 16133 13369 16136
rect 13403 16133 13415 16167
rect 13357 16127 13415 16133
rect 2222 16056 2228 16108
rect 2280 16096 2286 16108
rect 2409 16099 2467 16105
rect 2409 16096 2421 16099
rect 2280 16068 2421 16096
rect 2280 16056 2286 16068
rect 2409 16065 2421 16068
rect 2455 16065 2467 16099
rect 2409 16059 2467 16065
rect 5721 16099 5779 16105
rect 5721 16065 5733 16099
rect 5767 16096 5779 16099
rect 5994 16096 6000 16108
rect 5767 16068 6000 16096
rect 5767 16065 5779 16068
rect 5721 16059 5779 16065
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 7098 16056 7104 16108
rect 7156 16096 7162 16108
rect 7469 16099 7527 16105
rect 7469 16096 7481 16099
rect 7156 16068 7481 16096
rect 7156 16056 7162 16068
rect 7469 16065 7481 16068
rect 7515 16065 7527 16099
rect 8662 16096 8668 16108
rect 8575 16068 8668 16096
rect 7469 16059 7527 16065
rect 8662 16056 8668 16068
rect 8720 16056 8726 16108
rect 11146 16096 11152 16108
rect 11107 16068 11152 16096
rect 11146 16056 11152 16068
rect 11204 16056 11210 16108
rect 15470 16056 15476 16108
rect 15528 16096 15534 16108
rect 15841 16099 15899 16105
rect 15841 16096 15853 16099
rect 15528 16068 15853 16096
rect 15528 16056 15534 16068
rect 15841 16065 15853 16068
rect 15887 16065 15899 16099
rect 15841 16059 15899 16065
rect 1394 15988 1400 16040
rect 1452 16028 1458 16040
rect 2593 16031 2651 16037
rect 2593 16028 2605 16031
rect 1452 16000 2605 16028
rect 1452 15988 1458 16000
rect 2593 15997 2605 16000
rect 2639 15997 2651 16031
rect 2593 15991 2651 15997
rect 4709 16031 4767 16037
rect 4709 15997 4721 16031
rect 4755 16028 4767 16031
rect 6454 16028 6460 16040
rect 4755 16000 6460 16028
rect 4755 15997 4767 16000
rect 4709 15991 4767 15997
rect 3421 15963 3479 15969
rect 3421 15929 3433 15963
rect 3467 15960 3479 15963
rect 3694 15960 3700 15972
rect 3467 15932 3700 15960
rect 3467 15929 3479 15932
rect 3421 15923 3479 15929
rect 3694 15920 3700 15932
rect 3752 15920 3758 15972
rect 5736 15969 5764 16000
rect 6454 15988 6460 16000
rect 6512 16028 6518 16040
rect 6638 16028 6644 16040
rect 6512 16000 6644 16028
rect 6512 15988 6518 16000
rect 6638 15988 6644 16000
rect 6696 15988 6702 16040
rect 8754 15988 8760 16040
rect 8812 16028 8818 16040
rect 8921 16031 8979 16037
rect 8921 16028 8933 16031
rect 8812 16000 8933 16028
rect 8812 15988 8818 16000
rect 8921 15997 8933 16000
rect 8967 15997 8979 16031
rect 8921 15991 8979 15997
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 15997 13967 16031
rect 13909 15991 13967 15997
rect 5721 15963 5779 15969
rect 5721 15929 5733 15963
rect 5767 15929 5779 15963
rect 5721 15923 5779 15929
rect 5810 15920 5816 15972
rect 5868 15960 5874 15972
rect 7193 15963 7251 15969
rect 7193 15960 7205 15963
rect 5868 15932 5913 15960
rect 6564 15932 7205 15960
rect 5868 15920 5874 15932
rect 1946 15852 1952 15904
rect 2004 15892 2010 15904
rect 2501 15895 2559 15901
rect 2501 15892 2513 15895
rect 2004 15864 2513 15892
rect 2004 15852 2010 15864
rect 2501 15861 2513 15864
rect 2547 15861 2559 15895
rect 2501 15855 2559 15861
rect 3053 15895 3111 15901
rect 3053 15861 3065 15895
rect 3099 15892 3111 15895
rect 3234 15892 3240 15904
rect 3099 15864 3240 15892
rect 3099 15861 3111 15864
rect 3053 15855 3111 15861
rect 3234 15852 3240 15864
rect 3292 15852 3298 15904
rect 3510 15892 3516 15904
rect 3471 15864 3516 15892
rect 3510 15852 3516 15864
rect 3568 15852 3574 15904
rect 3878 15852 3884 15904
rect 3936 15892 3942 15904
rect 4341 15895 4399 15901
rect 4341 15892 4353 15895
rect 3936 15864 4353 15892
rect 3936 15852 3942 15864
rect 4341 15861 4353 15864
rect 4387 15892 4399 15895
rect 5810 15892 5838 15920
rect 6178 15892 6184 15904
rect 4387 15864 5838 15892
rect 6139 15864 6184 15892
rect 4387 15861 4399 15864
rect 4341 15855 4399 15861
rect 6178 15852 6184 15864
rect 6236 15892 6242 15904
rect 6564 15901 6592 15932
rect 7193 15929 7205 15932
rect 7239 15929 7251 15963
rect 7374 15960 7380 15972
rect 7335 15932 7380 15960
rect 7193 15923 7251 15929
rect 7374 15920 7380 15932
rect 7432 15920 7438 15972
rect 11882 15920 11888 15972
rect 11940 15960 11946 15972
rect 11977 15963 12035 15969
rect 11977 15960 11989 15963
rect 11940 15932 11989 15960
rect 11940 15920 11946 15932
rect 11977 15929 11989 15932
rect 12023 15960 12035 15963
rect 12894 15960 12900 15972
rect 12023 15932 12900 15960
rect 12023 15929 12035 15932
rect 11977 15923 12035 15929
rect 12894 15920 12900 15932
rect 12952 15960 12958 15972
rect 13924 15960 13952 15991
rect 13998 15988 14004 16040
rect 14056 16028 14062 16040
rect 14165 16031 14223 16037
rect 14165 16028 14177 16031
rect 14056 16000 14177 16028
rect 14056 15988 14062 16000
rect 14165 15997 14177 16000
rect 14211 15997 14223 16031
rect 16666 16028 16672 16040
rect 16627 16000 16672 16028
rect 14165 15991 14223 15997
rect 16666 15988 16672 16000
rect 16724 16028 16730 16040
rect 17405 16031 17463 16037
rect 17405 16028 17417 16031
rect 16724 16000 17417 16028
rect 16724 15988 16730 16000
rect 17405 15997 17417 16000
rect 17451 15997 17463 16031
rect 17405 15991 17463 15997
rect 12952 15932 13952 15960
rect 12952 15920 12958 15932
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 6236 15864 6561 15892
rect 6236 15852 6242 15864
rect 6549 15861 6561 15864
rect 6595 15861 6607 15895
rect 6549 15855 6607 15861
rect 9950 15852 9956 15904
rect 10008 15892 10014 15904
rect 10045 15895 10103 15901
rect 10045 15892 10057 15895
rect 10008 15864 10057 15892
rect 10008 15852 10014 15864
rect 10045 15861 10057 15864
rect 10091 15861 10103 15895
rect 12710 15892 12716 15904
rect 12671 15864 12716 15892
rect 10045 15855 10103 15861
rect 12710 15852 12716 15864
rect 12768 15852 12774 15904
rect 13817 15895 13875 15901
rect 13817 15861 13829 15895
rect 13863 15892 13875 15895
rect 13924 15892 13952 15932
rect 16945 15963 17003 15969
rect 16945 15929 16957 15963
rect 16991 15960 17003 15963
rect 18414 15960 18420 15972
rect 16991 15932 18420 15960
rect 16991 15929 17003 15932
rect 16945 15923 17003 15929
rect 18414 15920 18420 15932
rect 18472 15920 18478 15972
rect 14550 15892 14556 15904
rect 13863 15864 14556 15892
rect 13863 15861 13875 15864
rect 13817 15855 13875 15861
rect 14550 15852 14556 15864
rect 14608 15852 14614 15904
rect 15289 15895 15347 15901
rect 15289 15861 15301 15895
rect 15335 15892 15347 15895
rect 15470 15892 15476 15904
rect 15335 15864 15476 15892
rect 15335 15861 15347 15864
rect 15289 15855 15347 15861
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 5261 15691 5319 15697
rect 5261 15657 5273 15691
rect 5307 15688 5319 15691
rect 5994 15688 6000 15700
rect 5307 15660 6000 15688
rect 5307 15657 5319 15660
rect 5261 15651 5319 15657
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 7098 15648 7104 15700
rect 7156 15688 7162 15700
rect 7377 15691 7435 15697
rect 7377 15688 7389 15691
rect 7156 15660 7389 15688
rect 7156 15648 7162 15660
rect 7377 15657 7389 15660
rect 7423 15657 7435 15691
rect 7377 15651 7435 15657
rect 8754 15648 8760 15700
rect 8812 15688 8818 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 8812 15660 8953 15688
rect 8812 15648 8818 15660
rect 8941 15657 8953 15660
rect 8987 15657 8999 15691
rect 8941 15651 8999 15657
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 11609 15691 11667 15697
rect 11609 15688 11621 15691
rect 11112 15660 11621 15688
rect 11112 15648 11118 15660
rect 11609 15657 11621 15660
rect 11655 15657 11667 15691
rect 11609 15651 11667 15657
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 13909 15691 13967 15697
rect 13909 15688 13921 15691
rect 13872 15660 13921 15688
rect 13872 15648 13878 15660
rect 13909 15657 13921 15660
rect 13955 15688 13967 15691
rect 13998 15688 14004 15700
rect 13955 15660 14004 15688
rect 13955 15657 13967 15660
rect 13909 15651 13967 15657
rect 13998 15648 14004 15660
rect 14056 15648 14062 15700
rect 5810 15580 5816 15632
rect 5868 15620 5874 15632
rect 7466 15620 7472 15632
rect 5868 15592 7472 15620
rect 5868 15580 5874 15592
rect 7466 15580 7472 15592
rect 7524 15580 7530 15632
rect 8110 15580 8116 15632
rect 8168 15620 8174 15632
rect 8481 15623 8539 15629
rect 8481 15620 8493 15623
rect 8168 15592 8493 15620
rect 8168 15580 8174 15592
rect 8481 15589 8493 15592
rect 8527 15589 8539 15623
rect 8481 15583 8539 15589
rect 8662 15580 8668 15632
rect 8720 15620 8726 15632
rect 10318 15620 10324 15632
rect 8720 15592 10324 15620
rect 8720 15580 8726 15592
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 2038 15552 2044 15564
rect 1443 15524 2044 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 2038 15512 2044 15524
rect 2096 15512 2102 15564
rect 2501 15555 2559 15561
rect 2501 15521 2513 15555
rect 2547 15552 2559 15555
rect 2590 15552 2596 15564
rect 2547 15524 2596 15552
rect 2547 15521 2559 15524
rect 2501 15515 2559 15521
rect 2590 15512 2596 15524
rect 2648 15512 2654 15564
rect 4430 15552 4436 15564
rect 4391 15524 4436 15552
rect 4430 15512 4436 15524
rect 4488 15512 4494 15564
rect 5442 15552 5448 15564
rect 5403 15524 5448 15552
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 5712 15555 5770 15561
rect 5712 15521 5724 15555
rect 5758 15552 5770 15555
rect 5994 15552 6000 15564
rect 5758 15524 6000 15552
rect 5758 15521 5770 15524
rect 5712 15515 5770 15521
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 8018 15552 8024 15564
rect 6840 15524 8024 15552
rect 3145 15419 3203 15425
rect 3145 15385 3157 15419
rect 3191 15416 3203 15419
rect 3326 15416 3332 15428
rect 3191 15388 3332 15416
rect 3191 15385 3203 15388
rect 3145 15379 3203 15385
rect 3326 15376 3332 15388
rect 3384 15376 3390 15428
rect 6840 15425 6868 15524
rect 8018 15512 8024 15524
rect 8076 15512 8082 15564
rect 8294 15552 8300 15564
rect 8255 15524 8300 15552
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 9692 15561 9720 15592
rect 10318 15580 10324 15592
rect 10376 15580 10382 15632
rect 15841 15623 15899 15629
rect 15841 15589 15853 15623
rect 15887 15620 15899 15623
rect 15930 15620 15936 15632
rect 15887 15592 15936 15620
rect 15887 15589 15899 15592
rect 15841 15583 15899 15589
rect 15930 15580 15936 15592
rect 15988 15620 15994 15632
rect 16927 15623 16985 15629
rect 16927 15620 16939 15623
rect 15988 15592 16939 15620
rect 15988 15580 15994 15592
rect 16927 15589 16939 15592
rect 16973 15589 16985 15623
rect 17218 15620 17224 15632
rect 17179 15592 17224 15620
rect 16927 15583 16985 15589
rect 17218 15580 17224 15592
rect 17276 15580 17282 15632
rect 17402 15620 17408 15632
rect 17363 15592 17408 15620
rect 17402 15580 17408 15592
rect 17460 15580 17466 15632
rect 9950 15561 9956 15564
rect 9677 15555 9735 15561
rect 9677 15521 9689 15555
rect 9723 15552 9735 15555
rect 9944 15552 9956 15561
rect 9723 15524 9757 15552
rect 9911 15524 9956 15552
rect 9723 15521 9735 15524
rect 9677 15515 9735 15521
rect 9944 15515 9956 15524
rect 9950 15512 9956 15515
rect 10008 15512 10014 15564
rect 12710 15512 12716 15564
rect 12768 15552 12774 15564
rect 12768 15524 14044 15552
rect 12768 15512 12774 15524
rect 8573 15487 8631 15493
rect 8573 15484 8585 15487
rect 7760 15456 8585 15484
rect 6825 15419 6883 15425
rect 6825 15385 6837 15419
rect 6871 15385 6883 15419
rect 6825 15379 6883 15385
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 2314 15348 2320 15360
rect 2275 15320 2320 15348
rect 2314 15308 2320 15320
rect 2372 15308 2378 15360
rect 2682 15348 2688 15360
rect 2643 15320 2688 15348
rect 2682 15308 2688 15320
rect 2740 15308 2746 15360
rect 3418 15348 3424 15360
rect 3379 15320 3424 15348
rect 3418 15308 3424 15320
rect 3476 15308 3482 15360
rect 3786 15348 3792 15360
rect 3747 15320 3792 15348
rect 3786 15308 3792 15320
rect 3844 15308 3850 15360
rect 7650 15308 7656 15360
rect 7708 15348 7714 15360
rect 7760 15357 7788 15456
rect 8573 15453 8585 15456
rect 8619 15484 8631 15487
rect 8754 15484 8760 15496
rect 8619 15456 8760 15484
rect 8619 15453 8631 15456
rect 8573 15447 8631 15453
rect 8754 15444 8760 15456
rect 8812 15444 8818 15496
rect 13906 15484 13912 15496
rect 13867 15456 13912 15484
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 14016 15493 14044 15524
rect 15286 15512 15292 15564
rect 15344 15552 15350 15564
rect 15657 15555 15715 15561
rect 15657 15552 15669 15555
rect 15344 15524 15669 15552
rect 15344 15512 15350 15524
rect 15657 15521 15669 15524
rect 15703 15521 15715 15555
rect 18414 15552 18420 15564
rect 18375 15524 18420 15552
rect 15657 15515 15715 15521
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 14001 15487 14059 15493
rect 14001 15453 14013 15487
rect 14047 15484 14059 15487
rect 14550 15484 14556 15496
rect 14047 15456 14556 15484
rect 14047 15453 14059 15456
rect 14001 15447 14059 15453
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 15933 15487 15991 15493
rect 15933 15453 15945 15487
rect 15979 15484 15991 15487
rect 16114 15484 16120 15496
rect 15979 15456 16120 15484
rect 15979 15453 15991 15456
rect 15933 15447 15991 15453
rect 16114 15444 16120 15456
rect 16172 15444 16178 15496
rect 17497 15487 17555 15493
rect 17497 15453 17509 15487
rect 17543 15484 17555 15487
rect 18230 15484 18236 15496
rect 17543 15456 18236 15484
rect 17543 15453 17555 15456
rect 17497 15447 17555 15453
rect 13924 15416 13952 15444
rect 14366 15416 14372 15428
rect 13924 15388 14372 15416
rect 14366 15376 14372 15388
rect 14424 15376 14430 15428
rect 15105 15419 15163 15425
rect 15105 15385 15117 15419
rect 15151 15416 15163 15419
rect 15562 15416 15568 15428
rect 15151 15388 15568 15416
rect 15151 15385 15163 15388
rect 15105 15379 15163 15385
rect 15562 15376 15568 15388
rect 15620 15416 15626 15428
rect 17512 15416 17540 15447
rect 18230 15444 18236 15456
rect 18288 15444 18294 15496
rect 15620 15388 17540 15416
rect 15620 15376 15626 15388
rect 7745 15351 7803 15357
rect 7745 15348 7757 15351
rect 7708 15320 7757 15348
rect 7708 15308 7714 15320
rect 7745 15317 7757 15320
rect 7791 15317 7803 15351
rect 8018 15348 8024 15360
rect 7979 15320 8024 15348
rect 7745 15311 7803 15317
rect 8018 15308 8024 15320
rect 8076 15308 8082 15360
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 9858 15348 9864 15360
rect 9539 15320 9864 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 9858 15308 9864 15320
rect 9916 15308 9922 15360
rect 11057 15351 11115 15357
rect 11057 15317 11069 15351
rect 11103 15348 11115 15351
rect 11146 15348 11152 15360
rect 11103 15320 11152 15348
rect 11103 15317 11115 15320
rect 11057 15311 11115 15317
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 12621 15351 12679 15357
rect 12621 15317 12633 15351
rect 12667 15348 12679 15351
rect 13078 15348 13084 15360
rect 12667 15320 13084 15348
rect 12667 15317 12679 15320
rect 12621 15311 12679 15317
rect 13078 15308 13084 15320
rect 13136 15348 13142 15360
rect 13449 15351 13507 15357
rect 13449 15348 13461 15351
rect 13136 15320 13461 15348
rect 13136 15308 13142 15320
rect 13449 15317 13461 15320
rect 13495 15317 13507 15351
rect 15378 15348 15384 15360
rect 15339 15320 15384 15348
rect 13449 15311 13507 15317
rect 15378 15308 15384 15320
rect 15436 15308 15442 15360
rect 18601 15351 18659 15357
rect 18601 15317 18613 15351
rect 18647 15348 18659 15351
rect 20254 15348 20260 15360
rect 18647 15320 20260 15348
rect 18647 15317 18659 15320
rect 18601 15311 18659 15317
rect 20254 15308 20260 15320
rect 20312 15308 20318 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2038 15144 2044 15156
rect 1999 15116 2044 15144
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 2590 15144 2596 15156
rect 2551 15116 2596 15144
rect 2590 15104 2596 15116
rect 2648 15104 2654 15156
rect 3510 15104 3516 15156
rect 3568 15144 3574 15156
rect 3881 15147 3939 15153
rect 3881 15144 3893 15147
rect 3568 15116 3893 15144
rect 3568 15104 3574 15116
rect 3881 15113 3893 15116
rect 3927 15144 3939 15147
rect 5442 15144 5448 15156
rect 3927 15116 4936 15144
rect 5403 15116 5448 15144
rect 3927 15113 3939 15116
rect 3881 15107 3939 15113
rect 2961 15079 3019 15085
rect 2961 15045 2973 15079
rect 3007 15045 3019 15079
rect 2961 15039 3019 15045
rect 2976 15008 3004 15039
rect 3234 15036 3240 15088
rect 3292 15076 3298 15088
rect 4525 15079 4583 15085
rect 4525 15076 4537 15079
rect 3292 15048 4537 15076
rect 3292 15036 3298 15048
rect 4525 15045 4537 15048
rect 4571 15045 4583 15079
rect 4525 15039 4583 15045
rect 4062 15008 4068 15020
rect 2976 14980 4068 15008
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 4246 15008 4252 15020
rect 4207 14980 4252 15008
rect 4246 14968 4252 14980
rect 4304 14968 4310 15020
rect 4908 15017 4936 15116
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 5905 15147 5963 15153
rect 5905 15113 5917 15147
rect 5951 15144 5963 15147
rect 5994 15144 6000 15156
rect 5951 15116 6000 15144
rect 5951 15113 5963 15116
rect 5905 15107 5963 15113
rect 5994 15104 6000 15116
rect 6052 15104 6058 15156
rect 7006 15104 7012 15156
rect 7064 15144 7070 15156
rect 7929 15147 7987 15153
rect 7929 15144 7941 15147
rect 7064 15116 7941 15144
rect 7064 15104 7070 15116
rect 7929 15113 7941 15116
rect 7975 15144 7987 15147
rect 8110 15144 8116 15156
rect 7975 15116 8116 15144
rect 7975 15113 7987 15116
rect 7929 15107 7987 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 8294 15144 8300 15156
rect 8255 15116 8300 15144
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 8757 15147 8815 15153
rect 8757 15113 8769 15147
rect 8803 15144 8815 15147
rect 9950 15144 9956 15156
rect 8803 15116 9956 15144
rect 8803 15113 8815 15116
rect 8757 15107 8815 15113
rect 6914 15076 6920 15088
rect 6875 15048 6920 15076
rect 6914 15036 6920 15048
rect 6972 15036 6978 15088
rect 7466 15036 7472 15088
rect 7524 15076 7530 15088
rect 8772 15076 8800 15107
rect 7524 15048 8800 15076
rect 7524 15036 7530 15048
rect 9122 15036 9128 15088
rect 9180 15076 9186 15088
rect 9309 15079 9367 15085
rect 9309 15076 9321 15079
rect 9180 15048 9321 15076
rect 9180 15036 9186 15048
rect 9309 15045 9321 15048
rect 9355 15045 9367 15079
rect 9309 15039 9367 15045
rect 4893 15011 4951 15017
rect 4893 14977 4905 15011
rect 4939 14977 4951 15011
rect 4893 14971 4951 14977
rect 6178 14968 6184 15020
rect 6236 15008 6242 15020
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 6236 14980 7389 15008
rect 6236 14968 6242 14980
rect 7377 14977 7389 14980
rect 7423 15008 7435 15011
rect 8018 15008 8024 15020
rect 7423 14980 8024 15008
rect 7423 14977 7435 14980
rect 7377 14971 7435 14977
rect 8018 14968 8024 14980
rect 8076 14968 8082 15020
rect 9876 15017 9904 15116
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 10318 15144 10324 15156
rect 10231 15116 10324 15144
rect 10318 15104 10324 15116
rect 10376 15144 10382 15156
rect 11882 15144 11888 15156
rect 10376 15116 11888 15144
rect 10376 15104 10382 15116
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 12621 15147 12679 15153
rect 12621 15113 12633 15147
rect 12667 15144 12679 15147
rect 13262 15144 13268 15156
rect 12667 15116 13268 15144
rect 12667 15113 12679 15116
rect 12621 15107 12679 15113
rect 13262 15104 13268 15116
rect 13320 15104 13326 15156
rect 13633 15147 13691 15153
rect 13633 15113 13645 15147
rect 13679 15144 13691 15147
rect 13722 15144 13728 15156
rect 13679 15116 13728 15144
rect 13679 15113 13691 15116
rect 13633 15107 13691 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 13998 15144 14004 15156
rect 13959 15116 14004 15144
rect 13998 15104 14004 15116
rect 14056 15104 14062 15156
rect 16114 15104 16120 15156
rect 16172 15144 16178 15156
rect 16577 15147 16635 15153
rect 16577 15144 16589 15147
rect 16172 15116 16589 15144
rect 16172 15104 16178 15116
rect 16577 15113 16589 15116
rect 16623 15113 16635 15147
rect 17218 15144 17224 15156
rect 17179 15116 17224 15144
rect 16577 15107 16635 15113
rect 17218 15104 17224 15116
rect 17276 15104 17282 15156
rect 17402 15104 17408 15156
rect 17460 15144 17466 15156
rect 17497 15147 17555 15153
rect 17497 15144 17509 15147
rect 17460 15116 17509 15144
rect 17460 15104 17466 15116
rect 17497 15113 17509 15116
rect 17543 15113 17555 15147
rect 18230 15144 18236 15156
rect 18191 15116 18236 15144
rect 17497 15107 17555 15113
rect 18230 15104 18236 15116
rect 18288 15104 18294 15156
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 18601 15147 18659 15153
rect 18601 15144 18613 15147
rect 18472 15116 18613 15144
rect 18472 15104 18478 15116
rect 18601 15113 18613 15116
rect 18647 15113 18659 15147
rect 18601 15107 18659 15113
rect 10873 15079 10931 15085
rect 10873 15045 10885 15079
rect 10919 15076 10931 15079
rect 11146 15076 11152 15088
rect 10919 15048 11152 15076
rect 10919 15045 10931 15048
rect 10873 15039 10931 15045
rect 11146 15036 11152 15048
rect 11204 15036 11210 15088
rect 12253 15079 12311 15085
rect 12253 15045 12265 15079
rect 12299 15076 12311 15079
rect 12434 15076 12440 15088
rect 12299 15048 12440 15076
rect 12299 15045 12311 15048
rect 12253 15039 12311 15045
rect 12434 15036 12440 15048
rect 12492 15036 12498 15088
rect 9861 15011 9919 15017
rect 9861 14977 9873 15011
rect 9907 14977 9919 15011
rect 9861 14971 9919 14977
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 1670 14940 1676 14952
rect 1443 14912 1676 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 1670 14900 1676 14912
rect 1728 14940 1734 14952
rect 1946 14940 1952 14952
rect 1728 14912 1952 14940
rect 1728 14900 1734 14912
rect 1946 14900 1952 14912
rect 2004 14900 2010 14952
rect 3234 14940 3240 14952
rect 3195 14912 3240 14940
rect 3234 14900 3240 14912
rect 3292 14900 3298 14952
rect 3326 14900 3332 14952
rect 3384 14940 3390 14952
rect 3513 14943 3571 14949
rect 3513 14940 3525 14943
rect 3384 14912 3525 14940
rect 3384 14900 3390 14912
rect 3513 14909 3525 14912
rect 3559 14909 3571 14943
rect 3513 14903 3571 14909
rect 14642 14900 14648 14952
rect 14700 14940 14706 14952
rect 15197 14943 15255 14949
rect 15197 14940 15209 14943
rect 14700 14912 15209 14940
rect 14700 14900 14706 14912
rect 15197 14909 15209 14912
rect 15243 14940 15255 14943
rect 15243 14912 15700 14940
rect 15243 14909 15255 14912
rect 15197 14903 15255 14909
rect 3418 14872 3424 14884
rect 3379 14844 3424 14872
rect 3418 14832 3424 14844
rect 3476 14832 3482 14884
rect 3602 14832 3608 14884
rect 3660 14872 3666 14884
rect 5077 14875 5135 14881
rect 5077 14872 5089 14875
rect 3660 14844 5089 14872
rect 3660 14832 3666 14844
rect 5077 14841 5089 14844
rect 5123 14872 5135 14875
rect 6181 14875 6239 14881
rect 6181 14872 6193 14875
rect 5123 14844 6193 14872
rect 5123 14841 5135 14844
rect 5077 14835 5135 14841
rect 6181 14841 6193 14844
rect 6227 14841 6239 14875
rect 7469 14875 7527 14881
rect 7469 14872 7481 14875
rect 6181 14835 6239 14841
rect 6748 14844 7481 14872
rect 6748 14816 6776 14844
rect 7469 14841 7481 14844
rect 7515 14872 7527 14875
rect 8386 14872 8392 14884
rect 7515 14844 8392 14872
rect 7515 14841 7527 14844
rect 7469 14835 7527 14841
rect 8386 14832 8392 14844
rect 8444 14832 8450 14884
rect 9585 14875 9643 14881
rect 9585 14872 9597 14875
rect 9048 14844 9597 14872
rect 9048 14816 9076 14844
rect 9585 14841 9597 14844
rect 9631 14841 9643 14875
rect 9585 14835 9643 14841
rect 9950 14832 9956 14884
rect 10008 14872 10014 14884
rect 10689 14875 10747 14881
rect 10689 14872 10701 14875
rect 10008 14844 10701 14872
rect 10008 14832 10014 14844
rect 10689 14841 10701 14844
rect 10735 14872 10747 14875
rect 11149 14875 11207 14881
rect 11149 14872 11161 14875
rect 10735 14844 11161 14872
rect 10735 14841 10747 14844
rect 10689 14835 10747 14841
rect 11149 14841 11161 14844
rect 11195 14841 11207 14875
rect 11149 14835 11207 14841
rect 11425 14875 11483 14881
rect 11425 14841 11437 14875
rect 11471 14872 11483 14875
rect 11885 14875 11943 14881
rect 11885 14872 11897 14875
rect 11471 14844 11897 14872
rect 11471 14841 11483 14844
rect 11425 14835 11483 14841
rect 11885 14841 11897 14844
rect 11931 14872 11943 14875
rect 12526 14872 12532 14884
rect 11931 14844 12532 14872
rect 11931 14841 11943 14844
rect 11885 14835 11943 14841
rect 12526 14832 12532 14844
rect 12584 14832 12590 14884
rect 12894 14872 12900 14884
rect 12855 14844 12900 14872
rect 12894 14832 12900 14844
rect 12952 14832 12958 14884
rect 13078 14872 13084 14884
rect 13039 14844 13084 14872
rect 13078 14832 13084 14844
rect 13136 14832 13142 14884
rect 13173 14875 13231 14881
rect 13173 14841 13185 14875
rect 13219 14841 13231 14875
rect 13173 14835 13231 14841
rect 14737 14875 14795 14881
rect 14737 14841 14749 14875
rect 14783 14872 14795 14875
rect 15464 14875 15522 14881
rect 15464 14872 15476 14875
rect 14783 14844 15476 14872
rect 14783 14841 14795 14844
rect 14737 14835 14795 14841
rect 15464 14841 15476 14844
rect 15510 14872 15522 14875
rect 15562 14872 15568 14884
rect 15510 14844 15568 14872
rect 15510 14841 15522 14844
rect 15464 14835 15522 14841
rect 1486 14764 1492 14816
rect 1544 14804 1550 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 1544 14776 1593 14804
rect 1544 14764 1550 14776
rect 1581 14773 1593 14776
rect 1627 14773 1639 14807
rect 1581 14767 1639 14773
rect 2590 14764 2596 14816
rect 2648 14804 2654 14816
rect 2774 14804 2780 14816
rect 2648 14776 2780 14804
rect 2648 14764 2654 14776
rect 2774 14764 2780 14776
rect 2832 14764 2838 14816
rect 4246 14764 4252 14816
rect 4304 14804 4310 14816
rect 4985 14807 5043 14813
rect 4985 14804 4997 14807
rect 4304 14776 4997 14804
rect 4304 14764 4310 14776
rect 4985 14773 4997 14776
rect 5031 14773 5043 14807
rect 4985 14767 5043 14773
rect 6641 14807 6699 14813
rect 6641 14773 6653 14807
rect 6687 14804 6699 14807
rect 6730 14804 6736 14816
rect 6687 14776 6736 14804
rect 6687 14773 6699 14776
rect 6641 14767 6699 14773
rect 6730 14764 6736 14776
rect 6788 14764 6794 14816
rect 7374 14804 7380 14816
rect 7335 14776 7380 14804
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 9030 14804 9036 14816
rect 8991 14776 9036 14804
rect 9030 14764 9036 14776
rect 9088 14764 9094 14816
rect 9398 14764 9404 14816
rect 9456 14804 9462 14816
rect 9769 14807 9827 14813
rect 9769 14804 9781 14807
rect 9456 14776 9781 14804
rect 9456 14764 9462 14776
rect 9769 14773 9781 14776
rect 9815 14773 9827 14807
rect 9769 14767 9827 14773
rect 11054 14764 11060 14816
rect 11112 14804 11118 14816
rect 11333 14807 11391 14813
rect 11333 14804 11345 14807
rect 11112 14776 11345 14804
rect 11112 14764 11118 14776
rect 11333 14773 11345 14776
rect 11379 14773 11391 14807
rect 11333 14767 11391 14773
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 13188 14804 13216 14835
rect 15562 14832 15568 14844
rect 15620 14832 15626 14884
rect 15672 14816 15700 14912
rect 12492 14776 13216 14804
rect 14369 14807 14427 14813
rect 12492 14764 12498 14776
rect 14369 14773 14381 14807
rect 14415 14804 14427 14807
rect 14550 14804 14556 14816
rect 14415 14776 14556 14804
rect 14415 14773 14427 14776
rect 14369 14767 14427 14773
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 15105 14807 15163 14813
rect 15105 14773 15117 14807
rect 15151 14804 15163 14807
rect 15654 14804 15660 14816
rect 15151 14776 15660 14804
rect 15151 14773 15163 14776
rect 15105 14767 15163 14773
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2038 14560 2044 14612
rect 2096 14600 2102 14612
rect 2590 14600 2596 14612
rect 2096 14572 2596 14600
rect 2096 14560 2102 14572
rect 2590 14560 2596 14572
rect 2648 14600 2654 14612
rect 2961 14603 3019 14609
rect 2961 14600 2973 14603
rect 2648 14572 2973 14600
rect 2648 14560 2654 14572
rect 2961 14569 2973 14572
rect 3007 14569 3019 14603
rect 3234 14600 3240 14612
rect 2961 14563 3019 14569
rect 3068 14572 3240 14600
rect 2777 14535 2835 14541
rect 2777 14501 2789 14535
rect 2823 14532 2835 14535
rect 2866 14532 2872 14544
rect 2823 14504 2872 14532
rect 2823 14501 2835 14504
rect 2777 14495 2835 14501
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 3068 14541 3096 14572
rect 3234 14560 3240 14572
rect 3292 14600 3298 14612
rect 3513 14603 3571 14609
rect 3513 14600 3525 14603
rect 3292 14572 3525 14600
rect 3292 14560 3298 14572
rect 3513 14569 3525 14572
rect 3559 14600 3571 14603
rect 3602 14600 3608 14612
rect 3559 14572 3608 14600
rect 3559 14569 3571 14572
rect 3513 14563 3571 14569
rect 3602 14560 3608 14572
rect 3660 14560 3666 14612
rect 4798 14560 4804 14612
rect 4856 14600 4862 14612
rect 5445 14603 5503 14609
rect 5445 14600 5457 14603
rect 4856 14572 5457 14600
rect 4856 14560 4862 14572
rect 5445 14569 5457 14572
rect 5491 14600 5503 14603
rect 5994 14600 6000 14612
rect 5491 14572 6000 14600
rect 5491 14569 5503 14572
rect 5445 14563 5503 14569
rect 5994 14560 6000 14572
rect 6052 14560 6058 14612
rect 6178 14600 6184 14612
rect 6139 14572 6184 14600
rect 6178 14560 6184 14572
rect 6236 14560 6242 14612
rect 8386 14600 8392 14612
rect 8347 14572 8392 14600
rect 8386 14560 8392 14572
rect 8444 14560 8450 14612
rect 9769 14603 9827 14609
rect 9769 14569 9781 14603
rect 9815 14600 9827 14603
rect 9950 14600 9956 14612
rect 9815 14572 9956 14600
rect 9815 14569 9827 14572
rect 9769 14563 9827 14569
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 10042 14560 10048 14612
rect 10100 14600 10106 14612
rect 10229 14603 10287 14609
rect 10229 14600 10241 14603
rect 10100 14572 10241 14600
rect 10100 14560 10106 14572
rect 10229 14569 10241 14572
rect 10275 14569 10287 14603
rect 10229 14563 10287 14569
rect 12805 14603 12863 14609
rect 12805 14569 12817 14603
rect 12851 14600 12863 14603
rect 12894 14600 12900 14612
rect 12851 14572 12900 14600
rect 12851 14569 12863 14572
rect 12805 14563 12863 14569
rect 12894 14560 12900 14572
rect 12952 14560 12958 14612
rect 13173 14603 13231 14609
rect 13173 14569 13185 14603
rect 13219 14600 13231 14603
rect 15102 14600 15108 14612
rect 13219 14572 13952 14600
rect 15063 14572 15108 14600
rect 13219 14569 13231 14572
rect 13173 14563 13231 14569
rect 3053 14535 3111 14541
rect 3053 14501 3065 14535
rect 3099 14501 3111 14535
rect 3053 14495 3111 14501
rect 3326 14492 3332 14544
rect 3384 14532 3390 14544
rect 4310 14535 4368 14541
rect 4310 14532 4322 14535
rect 3384 14504 4322 14532
rect 3384 14492 3390 14504
rect 4310 14501 4322 14504
rect 4356 14532 4368 14535
rect 4522 14532 4528 14544
rect 4356 14504 4528 14532
rect 4356 14501 4368 14504
rect 4310 14495 4368 14501
rect 4522 14492 4528 14504
rect 4580 14492 4586 14544
rect 5534 14492 5540 14544
rect 5592 14532 5598 14544
rect 6457 14535 6515 14541
rect 6457 14532 6469 14535
rect 5592 14504 6469 14532
rect 5592 14492 5598 14504
rect 6457 14501 6469 14504
rect 6503 14532 6515 14535
rect 7374 14532 7380 14544
rect 6503 14504 7380 14532
rect 6503 14501 6515 14504
rect 6457 14495 6515 14501
rect 7374 14492 7380 14504
rect 7432 14492 7438 14544
rect 3510 14424 3516 14476
rect 3568 14464 3574 14476
rect 4065 14467 4123 14473
rect 4065 14464 4077 14467
rect 3568 14436 4077 14464
rect 3568 14424 3574 14436
rect 4065 14433 4077 14436
rect 4111 14464 4123 14467
rect 5442 14464 5448 14476
rect 4111 14436 5448 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14464 6791 14467
rect 7265 14467 7323 14473
rect 7265 14464 7277 14467
rect 6779 14436 7277 14464
rect 6779 14433 6791 14436
rect 6733 14427 6791 14433
rect 7265 14433 7277 14436
rect 7311 14464 7323 14467
rect 7650 14464 7656 14476
rect 7311 14436 7656 14464
rect 7311 14433 7323 14436
rect 7265 14427 7323 14433
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 11048 14467 11106 14473
rect 11048 14464 11060 14467
rect 10008 14436 11060 14464
rect 10008 14424 10014 14436
rect 11048 14433 11060 14436
rect 11094 14464 11106 14467
rect 13188 14464 13216 14563
rect 13924 14541 13952 14572
rect 15102 14560 15108 14572
rect 15160 14560 15166 14612
rect 15930 14600 15936 14612
rect 15891 14572 15936 14600
rect 15930 14560 15936 14572
rect 15988 14560 15994 14612
rect 17494 14600 17500 14612
rect 17455 14572 17500 14600
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 13817 14535 13875 14541
rect 13817 14501 13829 14535
rect 13863 14501 13875 14535
rect 13817 14495 13875 14501
rect 13909 14535 13967 14541
rect 13909 14501 13921 14535
rect 13955 14532 13967 14535
rect 15470 14532 15476 14544
rect 13955 14504 15476 14532
rect 13955 14501 13967 14504
rect 13909 14495 13967 14501
rect 11094 14436 13216 14464
rect 13832 14464 13860 14495
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 15565 14535 15623 14541
rect 15565 14501 15577 14535
rect 15611 14532 15623 14535
rect 16114 14532 16120 14544
rect 15611 14504 16120 14532
rect 15611 14501 15623 14504
rect 15565 14495 15623 14501
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 14642 14464 14648 14476
rect 13832 14436 14648 14464
rect 11094 14433 11106 14436
rect 11048 14427 11106 14433
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 16390 14473 16396 14476
rect 16384 14464 16396 14473
rect 16351 14436 16396 14464
rect 16384 14427 16396 14436
rect 16390 14424 16396 14427
rect 16448 14424 16454 14476
rect 3418 14356 3424 14408
rect 3476 14356 3482 14408
rect 5460 14396 5488 14424
rect 7009 14399 7067 14405
rect 7009 14396 7021 14399
rect 5460 14368 7021 14396
rect 7009 14365 7021 14368
rect 7055 14365 7067 14399
rect 7009 14359 7067 14365
rect 10594 14356 10600 14408
rect 10652 14396 10658 14408
rect 10781 14399 10839 14405
rect 10781 14396 10793 14399
rect 10652 14368 10793 14396
rect 10652 14356 10658 14368
rect 10781 14365 10793 14368
rect 10827 14365 10839 14399
rect 10781 14359 10839 14365
rect 13170 14356 13176 14408
rect 13228 14396 13234 14408
rect 13817 14399 13875 14405
rect 13817 14396 13829 14399
rect 13228 14368 13829 14396
rect 13228 14356 13234 14368
rect 13817 14365 13829 14368
rect 13863 14396 13875 14399
rect 14274 14396 14280 14408
rect 13863 14368 14280 14396
rect 13863 14365 13875 14368
rect 13817 14359 13875 14365
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 15654 14356 15660 14408
rect 15712 14396 15718 14408
rect 16117 14399 16175 14405
rect 16117 14396 16129 14399
rect 15712 14368 16129 14396
rect 15712 14356 15718 14368
rect 16117 14365 16129 14368
rect 16163 14365 16175 14399
rect 16117 14359 16175 14365
rect 2501 14331 2559 14337
rect 2501 14297 2513 14331
rect 2547 14328 2559 14331
rect 3436 14328 3464 14356
rect 2547 14300 3464 14328
rect 2547 14297 2559 14300
rect 2501 14291 2559 14297
rect 11882 14288 11888 14340
rect 11940 14328 11946 14340
rect 13357 14331 13415 14337
rect 13357 14328 13369 14331
rect 11940 14300 13369 14328
rect 11940 14288 11946 14300
rect 13357 14297 13369 14300
rect 13403 14297 13415 14331
rect 13357 14291 13415 14297
rect 1673 14263 1731 14269
rect 1673 14229 1685 14263
rect 1719 14260 1731 14263
rect 1946 14260 1952 14272
rect 1719 14232 1952 14260
rect 1719 14229 1731 14232
rect 1673 14223 1731 14229
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 2041 14263 2099 14269
rect 2041 14229 2053 14263
rect 2087 14260 2099 14263
rect 2130 14260 2136 14272
rect 2087 14232 2136 14260
rect 2087 14229 2099 14232
rect 2041 14223 2099 14229
rect 2130 14220 2136 14232
rect 2188 14220 2194 14272
rect 3881 14263 3939 14269
rect 3881 14229 3893 14263
rect 3927 14260 3939 14263
rect 4062 14260 4068 14272
rect 3927 14232 4068 14260
rect 3927 14229 3939 14232
rect 3881 14223 3939 14229
rect 4062 14220 4068 14232
rect 4120 14220 4126 14272
rect 5350 14220 5356 14272
rect 5408 14260 5414 14272
rect 6733 14263 6791 14269
rect 6733 14260 6745 14263
rect 5408 14232 6745 14260
rect 5408 14220 5414 14232
rect 6733 14229 6745 14232
rect 6779 14260 6791 14263
rect 6825 14263 6883 14269
rect 6825 14260 6837 14263
rect 6779 14232 6837 14260
rect 6779 14229 6791 14232
rect 6733 14223 6791 14229
rect 6825 14229 6837 14232
rect 6871 14229 6883 14263
rect 6825 14223 6883 14229
rect 9309 14263 9367 14269
rect 9309 14229 9321 14263
rect 9355 14260 9367 14263
rect 9398 14260 9404 14272
rect 9355 14232 9404 14260
rect 9355 14229 9367 14232
rect 9309 14223 9367 14229
rect 9398 14220 9404 14232
rect 9456 14220 9462 14272
rect 10689 14263 10747 14269
rect 10689 14229 10701 14263
rect 10735 14260 10747 14263
rect 11146 14260 11152 14272
rect 10735 14232 11152 14260
rect 10735 14229 10747 14232
rect 10689 14223 10747 14229
rect 11146 14220 11152 14232
rect 11204 14220 11210 14272
rect 12161 14263 12219 14269
rect 12161 14229 12173 14263
rect 12207 14260 12219 14263
rect 12526 14260 12532 14272
rect 12207 14232 12532 14260
rect 12207 14229 12219 14232
rect 12161 14223 12219 14229
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14090 14260 14096 14272
rect 13872 14232 14096 14260
rect 13872 14220 13878 14232
rect 14090 14220 14096 14232
rect 14148 14220 14154 14272
rect 14642 14260 14648 14272
rect 14603 14232 14648 14260
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2590 14056 2596 14068
rect 2551 14028 2596 14056
rect 2590 14016 2596 14028
rect 2648 14016 2654 14068
rect 2866 14016 2872 14068
rect 2924 14056 2930 14068
rect 2961 14059 3019 14065
rect 2961 14056 2973 14059
rect 2924 14028 2973 14056
rect 2924 14016 2930 14028
rect 2961 14025 2973 14028
rect 3007 14025 3019 14059
rect 3510 14056 3516 14068
rect 2961 14019 3019 14025
rect 3160 14028 3516 14056
rect 1670 13988 1676 14000
rect 1631 13960 1676 13988
rect 1670 13948 1676 13960
rect 1728 13948 1734 14000
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13920 2191 13923
rect 2314 13920 2320 13932
rect 2179 13892 2320 13920
rect 2179 13889 2191 13892
rect 2133 13883 2191 13889
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 3160 13929 3188 14028
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 4522 14056 4528 14068
rect 4483 14028 4528 14056
rect 4522 14016 4528 14028
rect 4580 14056 4586 14068
rect 5445 14059 5503 14065
rect 5445 14056 5457 14059
rect 4580 14028 5457 14056
rect 4580 14016 4586 14028
rect 5445 14025 5457 14028
rect 5491 14025 5503 14059
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 5445 14019 5503 14025
rect 6840 14028 8769 14056
rect 5534 13948 5540 14000
rect 5592 13988 5598 14000
rect 5813 13991 5871 13997
rect 5813 13988 5825 13991
rect 5592 13960 5825 13988
rect 5592 13948 5598 13960
rect 5813 13957 5825 13960
rect 5859 13957 5871 13991
rect 5813 13951 5871 13957
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13889 3203 13923
rect 3145 13883 3203 13889
rect 5169 13923 5227 13929
rect 5169 13889 5181 13923
rect 5215 13920 5227 13923
rect 5442 13920 5448 13932
rect 5215 13892 5448 13920
rect 5215 13889 5227 13892
rect 5169 13883 5227 13889
rect 5442 13880 5448 13892
rect 5500 13920 5506 13932
rect 5994 13920 6000 13932
rect 5500 13892 6000 13920
rect 5500 13880 5506 13892
rect 5994 13880 6000 13892
rect 6052 13920 6058 13932
rect 6840 13929 6868 14028
rect 8757 14025 8769 14028
rect 8803 14025 8815 14059
rect 9950 14056 9956 14068
rect 9911 14028 9956 14056
rect 8757 14019 8815 14025
rect 8772 13988 8800 14019
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 10594 14056 10600 14068
rect 10555 14028 10600 14056
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 14274 14016 14280 14068
rect 14332 14056 14338 14068
rect 14369 14059 14427 14065
rect 14369 14056 14381 14059
rect 14332 14028 14381 14056
rect 14332 14016 14338 14028
rect 14369 14025 14381 14028
rect 14415 14025 14427 14059
rect 14734 14056 14740 14068
rect 14695 14028 14740 14056
rect 14369 14019 14427 14025
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 10612 13988 10640 14016
rect 10870 13988 10876 14000
rect 8772 13960 10640 13988
rect 10831 13960 10876 13988
rect 10870 13948 10876 13960
rect 10928 13948 10934 14000
rect 14918 13948 14924 14000
rect 14976 13988 14982 14000
rect 15013 13991 15071 13997
rect 15013 13988 15025 13991
rect 14976 13960 15025 13988
rect 14976 13948 14982 13960
rect 15013 13957 15025 13960
rect 15059 13957 15071 13991
rect 15013 13951 15071 13957
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 6052 13892 6561 13920
rect 6052 13880 6058 13892
rect 6549 13889 6561 13892
rect 6595 13920 6607 13923
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6595 13892 6837 13920
rect 6595 13889 6607 13892
rect 6549 13883 6607 13889
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 15378 13920 15384 13932
rect 15160 13892 15384 13920
rect 15160 13880 15166 13892
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 3234 13812 3240 13864
rect 3292 13852 3298 13864
rect 3401 13855 3459 13861
rect 3401 13852 3413 13855
rect 3292 13824 3413 13852
rect 3292 13812 3298 13824
rect 3401 13821 3413 13824
rect 3447 13821 3459 13855
rect 3401 13815 3459 13821
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5132 13824 5641 13852
rect 5132 13812 5138 13824
rect 5629 13821 5641 13824
rect 5675 13852 5687 13855
rect 6181 13855 6239 13861
rect 6181 13852 6193 13855
rect 5675 13824 6193 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 6181 13821 6193 13824
rect 6227 13821 6239 13855
rect 7081 13855 7139 13861
rect 7081 13852 7093 13855
rect 6181 13815 6239 13821
rect 6932 13824 7093 13852
rect 2222 13784 2228 13796
rect 2183 13756 2228 13784
rect 2222 13744 2228 13756
rect 2280 13744 2286 13796
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 6932 13784 6960 13824
rect 7081 13821 7093 13824
rect 7127 13821 7139 13855
rect 11146 13852 11152 13864
rect 11107 13824 11152 13852
rect 7081 13815 7139 13821
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 12253 13855 12311 13861
rect 12253 13821 12265 13855
rect 12299 13852 12311 13855
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12299 13824 12449 13852
rect 12299 13821 12311 13824
rect 12253 13815 12311 13821
rect 12437 13821 12449 13824
rect 12483 13852 12495 13855
rect 15565 13855 15623 13861
rect 15565 13852 15577 13855
rect 12483 13824 12848 13852
rect 12483 13821 12495 13824
rect 12437 13815 12495 13821
rect 12820 13796 12848 13824
rect 15120 13824 15577 13852
rect 6788 13756 6960 13784
rect 10321 13787 10379 13793
rect 6788 13744 6794 13756
rect 10321 13753 10333 13787
rect 10367 13784 10379 13787
rect 11425 13787 11483 13793
rect 11425 13784 11437 13787
rect 10367 13756 11437 13784
rect 10367 13753 10379 13756
rect 10321 13747 10379 13753
rect 11425 13753 11437 13756
rect 11471 13784 11483 13787
rect 12342 13784 12348 13796
rect 11471 13756 12348 13784
rect 11471 13753 11483 13756
rect 11425 13747 11483 13753
rect 12342 13744 12348 13756
rect 12400 13744 12406 13796
rect 12526 13744 12532 13796
rect 12584 13784 12590 13796
rect 12682 13787 12740 13793
rect 12682 13784 12694 13787
rect 12584 13756 12694 13784
rect 12584 13744 12590 13756
rect 12682 13753 12694 13756
rect 12728 13753 12740 13787
rect 12682 13747 12740 13753
rect 12802 13744 12808 13796
rect 12860 13744 12866 13796
rect 14642 13744 14648 13796
rect 14700 13784 14706 13796
rect 14700 13756 14964 13784
rect 14700 13744 14706 13756
rect 2130 13716 2136 13728
rect 2091 13688 2136 13716
rect 2130 13676 2136 13688
rect 2188 13676 2194 13728
rect 8202 13716 8208 13728
rect 8163 13688 8208 13716
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 11330 13716 11336 13728
rect 11243 13688 11336 13716
rect 11330 13676 11336 13688
rect 11388 13716 11394 13728
rect 11793 13719 11851 13725
rect 11793 13716 11805 13719
rect 11388 13688 11805 13716
rect 11388 13676 11394 13688
rect 11793 13685 11805 13688
rect 11839 13685 11851 13719
rect 11793 13679 11851 13685
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 13817 13719 13875 13725
rect 13817 13716 13829 13719
rect 13780 13688 13829 13716
rect 13780 13676 13786 13688
rect 13817 13685 13829 13688
rect 13863 13685 13875 13719
rect 14936 13716 14964 13756
rect 15010 13744 15016 13796
rect 15068 13784 15074 13796
rect 15120 13784 15148 13824
rect 15565 13821 15577 13824
rect 15611 13852 15623 13855
rect 16390 13852 16396 13864
rect 15611 13824 16396 13852
rect 15611 13821 15623 13824
rect 15565 13815 15623 13821
rect 16390 13812 16396 13824
rect 16448 13852 16454 13864
rect 16485 13855 16543 13861
rect 16485 13852 16497 13855
rect 16448 13824 16497 13852
rect 16448 13812 16454 13824
rect 16485 13821 16497 13824
rect 16531 13852 16543 13855
rect 17034 13852 17040 13864
rect 16531 13824 17040 13852
rect 16531 13821 16543 13824
rect 16485 13815 16543 13821
rect 17034 13812 17040 13824
rect 17092 13812 17098 13864
rect 15068 13756 15148 13784
rect 15068 13744 15074 13756
rect 15473 13719 15531 13725
rect 15473 13716 15485 13719
rect 14936 13688 15485 13716
rect 13817 13679 13875 13685
rect 15473 13685 15485 13688
rect 15519 13685 15531 13719
rect 15473 13679 15531 13685
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 16117 13719 16175 13725
rect 16117 13716 16129 13719
rect 15712 13688 16129 13716
rect 15712 13676 15718 13688
rect 16117 13685 16129 13688
rect 16163 13685 16175 13719
rect 16117 13679 16175 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1673 13515 1731 13521
rect 1673 13481 1685 13515
rect 1719 13512 1731 13515
rect 2222 13512 2228 13524
rect 1719 13484 2228 13512
rect 1719 13481 1731 13484
rect 1673 13475 1731 13481
rect 2222 13472 2228 13484
rect 2280 13472 2286 13524
rect 2317 13515 2375 13521
rect 2317 13481 2329 13515
rect 2363 13512 2375 13515
rect 3234 13512 3240 13524
rect 2363 13484 3240 13512
rect 2363 13481 2375 13484
rect 2317 13475 2375 13481
rect 3234 13472 3240 13484
rect 3292 13472 3298 13524
rect 3510 13512 3516 13524
rect 3471 13484 3516 13512
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 6730 13512 6736 13524
rect 6691 13484 6736 13512
rect 6730 13472 6736 13484
rect 6788 13472 6794 13524
rect 7466 13512 7472 13524
rect 7427 13484 7472 13512
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 9217 13515 9275 13521
rect 9217 13481 9229 13515
rect 9263 13512 9275 13515
rect 9950 13512 9956 13524
rect 9263 13484 9956 13512
rect 9263 13481 9275 13484
rect 9217 13475 9275 13481
rect 9950 13472 9956 13484
rect 10008 13472 10014 13524
rect 10870 13472 10876 13524
rect 10928 13512 10934 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 10928 13484 11621 13512
rect 10928 13472 10934 13484
rect 11609 13481 11621 13484
rect 11655 13512 11667 13515
rect 11882 13512 11888 13524
rect 11655 13484 11888 13512
rect 11655 13481 11667 13484
rect 11609 13475 11667 13481
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 14645 13515 14703 13521
rect 14645 13481 14657 13515
rect 14691 13512 14703 13515
rect 15102 13512 15108 13524
rect 14691 13484 15108 13512
rect 14691 13481 14703 13484
rect 14645 13475 14703 13481
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 17034 13512 17040 13524
rect 16995 13484 17040 13512
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 2866 13404 2872 13456
rect 2924 13453 2930 13456
rect 2924 13447 2973 13453
rect 2924 13413 2927 13447
rect 2961 13413 2973 13447
rect 2924 13407 2973 13413
rect 3053 13447 3111 13453
rect 3053 13413 3065 13447
rect 3099 13444 3111 13447
rect 3878 13444 3884 13456
rect 3099 13416 3884 13444
rect 3099 13413 3111 13416
rect 3053 13407 3111 13413
rect 2924 13404 2930 13407
rect 3878 13404 3884 13416
rect 3936 13404 3942 13456
rect 4062 13404 4068 13456
rect 4120 13444 4126 13456
rect 4433 13447 4491 13453
rect 4433 13444 4445 13447
rect 4120 13416 4445 13444
rect 4120 13404 4126 13416
rect 4433 13413 4445 13416
rect 4479 13413 4491 13447
rect 4614 13444 4620 13456
rect 4575 13416 4620 13444
rect 4433 13407 4491 13413
rect 4614 13404 4620 13416
rect 4672 13444 4678 13456
rect 5445 13447 5503 13453
rect 5445 13444 5457 13447
rect 4672 13416 5457 13444
rect 4672 13404 4678 13416
rect 5445 13413 5457 13416
rect 5491 13413 5503 13447
rect 5445 13407 5503 13413
rect 6457 13447 6515 13453
rect 6457 13413 6469 13447
rect 6503 13444 6515 13447
rect 6914 13444 6920 13456
rect 6503 13416 6920 13444
rect 6503 13413 6515 13416
rect 6457 13407 6515 13413
rect 6914 13404 6920 13416
rect 6972 13444 6978 13456
rect 7285 13447 7343 13453
rect 7285 13444 7297 13447
rect 6972 13416 7297 13444
rect 6972 13404 6978 13416
rect 7285 13413 7297 13416
rect 7331 13413 7343 13447
rect 7285 13407 7343 13413
rect 12342 13404 12348 13456
rect 12400 13444 12406 13456
rect 12866 13447 12924 13453
rect 12866 13444 12878 13447
rect 12400 13416 12878 13444
rect 12400 13404 12406 13416
rect 12866 13413 12878 13416
rect 12912 13444 12924 13447
rect 13722 13444 13728 13456
rect 12912 13416 13728 13444
rect 12912 13413 12924 13416
rect 12866 13407 12924 13413
rect 13722 13404 13728 13416
rect 13780 13444 13786 13456
rect 14090 13444 14096 13456
rect 13780 13416 14096 13444
rect 13780 13404 13786 13416
rect 14090 13404 14096 13416
rect 14148 13404 14154 13456
rect 15010 13444 15016 13456
rect 14971 13416 15016 13444
rect 15010 13404 15016 13416
rect 15068 13404 15074 13456
rect 15924 13447 15982 13453
rect 15924 13413 15936 13447
rect 15970 13444 15982 13447
rect 16114 13444 16120 13456
rect 15970 13416 16120 13444
rect 15970 13413 15982 13416
rect 15924 13407 15982 13413
rect 16114 13404 16120 13416
rect 16172 13404 16178 13456
rect 2038 13336 2044 13388
rect 2096 13376 2102 13388
rect 2777 13379 2835 13385
rect 2777 13376 2789 13379
rect 2096 13348 2789 13376
rect 2096 13336 2102 13348
rect 2777 13345 2789 13348
rect 2823 13345 2835 13379
rect 2777 13339 2835 13345
rect 4709 13379 4767 13385
rect 4709 13345 4721 13379
rect 4755 13376 4767 13379
rect 4798 13376 4804 13388
rect 4755 13348 4804 13376
rect 4755 13345 4767 13348
rect 4709 13339 4767 13345
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 5629 13379 5687 13385
rect 5629 13345 5641 13379
rect 5675 13376 5687 13379
rect 6270 13376 6276 13388
rect 5675 13348 6276 13376
rect 5675 13345 5687 13348
rect 5629 13339 5687 13345
rect 6270 13336 6276 13348
rect 6328 13336 6334 13388
rect 11882 13336 11888 13388
rect 11940 13376 11946 13388
rect 12621 13379 12679 13385
rect 12621 13376 12633 13379
rect 11940 13348 12633 13376
rect 11940 13336 11946 13348
rect 12621 13345 12633 13348
rect 12667 13376 12679 13379
rect 12710 13376 12716 13388
rect 12667 13348 12716 13376
rect 12667 13345 12679 13348
rect 12621 13339 12679 13345
rect 12710 13336 12716 13348
rect 12768 13376 12774 13388
rect 18506 13376 18512 13388
rect 12768 13348 15700 13376
rect 18467 13348 18512 13376
rect 12768 13336 12774 13348
rect 15672 13320 15700 13348
rect 18506 13336 18512 13348
rect 18564 13336 18570 13388
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13308 7619 13311
rect 8202 13308 8208 13320
rect 7607 13280 8208 13308
rect 7607 13277 7619 13280
rect 7561 13271 7619 13277
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 10336 13280 11529 13308
rect 4154 13240 4160 13252
rect 4115 13212 4160 13240
rect 4154 13200 4160 13212
rect 4212 13200 4218 13252
rect 10336 13184 10364 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 11698 13308 11704 13320
rect 11659 13280 11704 13308
rect 11517 13271 11575 13277
rect 11698 13268 11704 13280
rect 11756 13308 11762 13320
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 11756 13280 12449 13308
rect 11756 13268 11762 13280
rect 12437 13277 12449 13280
rect 12483 13308 12495 13311
rect 12526 13308 12532 13320
rect 12483 13280 12532 13308
rect 12483 13277 12495 13280
rect 12437 13271 12495 13277
rect 12526 13268 12532 13280
rect 12584 13268 12590 13320
rect 15654 13308 15660 13320
rect 15615 13280 15660 13308
rect 15654 13268 15660 13280
rect 15712 13268 15718 13320
rect 18785 13311 18843 13317
rect 18785 13277 18797 13311
rect 18831 13308 18843 13311
rect 19426 13308 19432 13320
rect 18831 13280 19432 13308
rect 18831 13277 18843 13280
rect 18785 13271 18843 13277
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 11149 13243 11207 13249
rect 11149 13209 11161 13243
rect 11195 13240 11207 13243
rect 11330 13240 11336 13252
rect 11195 13212 11336 13240
rect 11195 13209 11207 13212
rect 11149 13203 11207 13209
rect 11330 13200 11336 13212
rect 11388 13200 11394 13252
rect 2501 13175 2559 13181
rect 2501 13141 2513 13175
rect 2547 13172 2559 13175
rect 3050 13172 3056 13184
rect 2547 13144 3056 13172
rect 2547 13141 2559 13144
rect 2501 13135 2559 13141
rect 3050 13132 3056 13144
rect 3108 13132 3114 13184
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 4062 13172 4068 13184
rect 3927 13144 4068 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 5074 13172 5080 13184
rect 5035 13144 5080 13172
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 5813 13175 5871 13181
rect 5813 13141 5825 13175
rect 5859 13172 5871 13175
rect 6086 13172 6092 13184
rect 5859 13144 6092 13172
rect 5859 13141 5871 13144
rect 5813 13135 5871 13141
rect 6086 13132 6092 13144
rect 6144 13132 6150 13184
rect 7006 13172 7012 13184
rect 6967 13144 7012 13172
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 7558 13132 7564 13184
rect 7616 13172 7622 13184
rect 7929 13175 7987 13181
rect 7929 13172 7941 13175
rect 7616 13144 7941 13172
rect 7616 13132 7622 13144
rect 7929 13141 7941 13144
rect 7975 13141 7987 13175
rect 7929 13135 7987 13141
rect 8389 13175 8447 13181
rect 8389 13141 8401 13175
rect 8435 13172 8447 13175
rect 8478 13172 8484 13184
rect 8435 13144 8484 13172
rect 8435 13141 8447 13144
rect 8389 13135 8447 13141
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 10318 13172 10324 13184
rect 10279 13144 10324 13172
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 10781 13175 10839 13181
rect 10781 13141 10793 13175
rect 10827 13172 10839 13175
rect 11054 13172 11060 13184
rect 10827 13144 11060 13172
rect 10827 13141 10839 13144
rect 10781 13135 10839 13141
rect 11054 13132 11060 13144
rect 11112 13172 11118 13184
rect 11422 13172 11428 13184
rect 11112 13144 11428 13172
rect 11112 13132 11118 13144
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 11514 13132 11520 13184
rect 11572 13172 11578 13184
rect 14001 13175 14059 13181
rect 14001 13172 14013 13175
rect 11572 13144 14013 13172
rect 11572 13132 11578 13144
rect 14001 13141 14013 13144
rect 14047 13141 14059 13175
rect 15470 13172 15476 13184
rect 15431 13144 15476 13172
rect 14001 13135 14059 13141
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2038 12968 2044 12980
rect 1999 12940 2044 12968
rect 2038 12928 2044 12940
rect 2096 12928 2102 12980
rect 2314 12928 2320 12980
rect 2372 12968 2378 12980
rect 2593 12971 2651 12977
rect 2593 12968 2605 12971
rect 2372 12940 2605 12968
rect 2372 12928 2378 12940
rect 2593 12937 2605 12940
rect 2639 12937 2651 12971
rect 2593 12931 2651 12937
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 3878 12968 3884 12980
rect 2832 12940 3096 12968
rect 3839 12940 3884 12968
rect 2832 12928 2838 12940
rect 1670 12860 1676 12912
rect 1728 12900 1734 12912
rect 2409 12903 2467 12909
rect 2409 12900 2421 12903
rect 1728 12872 2421 12900
rect 1728 12860 1734 12872
rect 2409 12869 2421 12872
rect 2455 12900 2467 12903
rect 2866 12900 2872 12912
rect 2455 12872 2872 12900
rect 2455 12869 2467 12872
rect 2409 12863 2467 12869
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 3068 12900 3096 12940
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4614 12968 4620 12980
rect 4203 12940 4620 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 4798 12928 4804 12980
rect 4856 12968 4862 12980
rect 5077 12971 5135 12977
rect 5077 12968 5089 12971
rect 4856 12940 5089 12968
rect 4856 12928 4862 12940
rect 5077 12937 5089 12940
rect 5123 12937 5135 12971
rect 5077 12931 5135 12937
rect 5537 12971 5595 12977
rect 5537 12937 5549 12971
rect 5583 12968 5595 12971
rect 6270 12968 6276 12980
rect 5583 12940 6276 12968
rect 5583 12937 5595 12940
rect 5537 12931 5595 12937
rect 6270 12928 6276 12940
rect 6328 12928 6334 12980
rect 8202 12968 8208 12980
rect 8163 12940 8208 12968
rect 8202 12928 8208 12940
rect 8260 12928 8266 12980
rect 9217 12971 9275 12977
rect 9217 12937 9229 12971
rect 9263 12968 9275 12971
rect 10318 12968 10324 12980
rect 9263 12940 10324 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 10778 12968 10784 12980
rect 10739 12940 10784 12968
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 11882 12968 11888 12980
rect 11843 12940 11888 12968
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 12894 12968 12900 12980
rect 12855 12940 12900 12968
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 14090 12968 14096 12980
rect 14051 12940 14096 12968
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 14642 12928 14648 12980
rect 14700 12968 14706 12980
rect 14737 12971 14795 12977
rect 14737 12968 14749 12971
rect 14700 12940 14749 12968
rect 14700 12928 14706 12940
rect 14737 12937 14749 12940
rect 14783 12937 14795 12971
rect 16114 12968 16120 12980
rect 16075 12940 16120 12968
rect 14737 12931 14795 12937
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 18506 12968 18512 12980
rect 18467 12940 18512 12968
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 5350 12900 5356 12912
rect 3068 12872 5356 12900
rect 3160 12841 3188 12872
rect 5350 12860 5356 12872
rect 5408 12860 5414 12912
rect 6914 12900 6920 12912
rect 6875 12872 6920 12900
rect 6914 12860 6920 12872
rect 6972 12860 6978 12912
rect 10229 12903 10287 12909
rect 10229 12869 10241 12903
rect 10275 12900 10287 12903
rect 10870 12900 10876 12912
rect 10275 12872 10876 12900
rect 10275 12869 10287 12872
rect 10229 12863 10287 12869
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 12710 12860 12716 12912
rect 12768 12900 12774 12912
rect 13078 12900 13084 12912
rect 12768 12872 13084 12900
rect 12768 12860 12774 12872
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 13173 12903 13231 12909
rect 13173 12869 13185 12903
rect 13219 12900 13231 12903
rect 13219 12872 15148 12900
rect 13219 12869 13231 12872
rect 13173 12863 13231 12869
rect 3145 12835 3203 12841
rect 3145 12801 3157 12835
rect 3191 12801 3203 12835
rect 3145 12795 3203 12801
rect 4338 12792 4344 12844
rect 4396 12832 4402 12844
rect 4617 12835 4675 12841
rect 4617 12832 4629 12835
rect 4396 12804 4629 12832
rect 4396 12792 4402 12804
rect 4617 12801 4629 12804
rect 4663 12832 4675 12835
rect 5074 12832 5080 12844
rect 4663 12804 5080 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 6273 12835 6331 12841
rect 6273 12801 6285 12835
rect 6319 12832 6331 12835
rect 6454 12832 6460 12844
rect 6319 12804 6460 12832
rect 6319 12801 6331 12804
rect 6273 12795 6331 12801
rect 1302 12724 1308 12776
rect 1360 12764 1366 12776
rect 1397 12767 1455 12773
rect 1397 12764 1409 12767
rect 1360 12736 1409 12764
rect 1360 12724 1366 12736
rect 1397 12733 1409 12736
rect 1443 12764 1455 12767
rect 1762 12764 1768 12776
rect 1443 12736 1768 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 2869 12767 2927 12773
rect 2869 12733 2881 12767
rect 2915 12764 2927 12767
rect 2915 12736 3648 12764
rect 2915 12733 2927 12736
rect 2869 12727 2927 12733
rect 3620 12705 3648 12736
rect 3878 12724 3884 12776
rect 3936 12764 3942 12776
rect 4430 12764 4436 12776
rect 3936 12736 4436 12764
rect 3936 12724 3942 12736
rect 4430 12724 4436 12736
rect 4488 12764 4494 12776
rect 4709 12767 4767 12773
rect 4709 12764 4721 12767
rect 4488 12736 4721 12764
rect 4488 12724 4494 12736
rect 4709 12733 4721 12736
rect 4755 12733 4767 12767
rect 4709 12727 4767 12733
rect 5629 12767 5687 12773
rect 5629 12733 5641 12767
rect 5675 12764 5687 12767
rect 6288 12764 6316 12795
rect 6454 12792 6460 12804
rect 6512 12792 6518 12844
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 7374 12832 7380 12844
rect 6687 12804 7380 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12832 9827 12835
rect 9950 12832 9956 12844
rect 9815 12804 9956 12832
rect 9815 12801 9827 12804
rect 9769 12795 9827 12801
rect 9950 12792 9956 12804
rect 10008 12792 10014 12844
rect 11054 12792 11060 12844
rect 11112 12832 11118 12844
rect 11333 12835 11391 12841
rect 11333 12832 11345 12835
rect 11112 12804 11345 12832
rect 11112 12792 11118 12804
rect 11333 12801 11345 12804
rect 11379 12801 11391 12835
rect 11333 12795 11391 12801
rect 11422 12792 11428 12844
rect 11480 12832 11486 12844
rect 15120 12841 15148 12872
rect 12253 12835 12311 12841
rect 12253 12832 12265 12835
rect 11480 12804 12265 12832
rect 11480 12792 11486 12804
rect 12253 12801 12265 12804
rect 12299 12832 12311 12835
rect 13541 12835 13599 12841
rect 13541 12832 13553 12835
rect 12299 12804 13553 12832
rect 12299 12801 12311 12804
rect 12253 12795 12311 12801
rect 13541 12801 13553 12804
rect 13587 12801 13599 12835
rect 13541 12795 13599 12801
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12832 15163 12835
rect 16393 12835 16451 12841
rect 16393 12832 16405 12835
rect 15151 12804 16405 12832
rect 15151 12801 15163 12804
rect 15105 12795 15163 12801
rect 16393 12801 16405 12804
rect 16439 12801 16451 12835
rect 16393 12795 16451 12801
rect 5675 12736 6316 12764
rect 5675 12733 5687 12736
rect 5629 12727 5687 12733
rect 6546 12724 6552 12776
rect 6604 12764 6610 12776
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 6604 12736 7849 12764
rect 6604 12724 6610 12736
rect 3605 12699 3663 12705
rect 3605 12665 3617 12699
rect 3651 12696 3663 12699
rect 3970 12696 3976 12708
rect 3651 12668 3976 12696
rect 3651 12665 3663 12668
rect 3605 12659 3663 12665
rect 3970 12656 3976 12668
rect 4028 12656 4034 12708
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 4522 12696 4528 12708
rect 4120 12668 4528 12696
rect 4120 12656 4126 12668
rect 4522 12656 4528 12668
rect 4580 12696 4586 12708
rect 7392 12705 7420 12736
rect 7837 12733 7849 12736
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 12894 12724 12900 12776
rect 12952 12764 12958 12776
rect 14553 12767 14611 12773
rect 12952 12736 13676 12764
rect 12952 12724 12958 12736
rect 4617 12699 4675 12705
rect 4617 12696 4629 12699
rect 4580 12668 4629 12696
rect 4580 12656 4586 12668
rect 4617 12665 4629 12668
rect 4663 12665 4675 12699
rect 4617 12659 4675 12665
rect 7377 12699 7435 12705
rect 7377 12665 7389 12699
rect 7423 12665 7435 12699
rect 7377 12659 7435 12665
rect 7469 12699 7527 12705
rect 7469 12665 7481 12699
rect 7515 12696 7527 12699
rect 8110 12696 8116 12708
rect 7515 12668 8116 12696
rect 7515 12665 7527 12668
rect 7469 12659 7527 12665
rect 8110 12656 8116 12668
rect 8168 12696 8174 12708
rect 8573 12699 8631 12705
rect 8573 12696 8585 12699
rect 8168 12668 8585 12696
rect 8168 12656 8174 12668
rect 8573 12665 8585 12668
rect 8619 12665 8631 12699
rect 8573 12659 8631 12665
rect 9398 12656 9404 12708
rect 9456 12696 9462 12708
rect 9493 12699 9551 12705
rect 9493 12696 9505 12699
rect 9456 12668 9505 12696
rect 9456 12656 9462 12668
rect 9493 12665 9505 12668
rect 9539 12665 9551 12699
rect 11054 12696 11060 12708
rect 11015 12668 11060 12696
rect 9493 12659 9551 12665
rect 11054 12656 11060 12668
rect 11112 12656 11118 12708
rect 13648 12705 13676 12736
rect 14553 12733 14565 12767
rect 14599 12764 14611 12767
rect 15289 12767 15347 12773
rect 15289 12764 15301 12767
rect 14599 12736 15301 12764
rect 14599 12733 14611 12736
rect 14553 12727 14611 12733
rect 15289 12733 15301 12736
rect 15335 12764 15347 12767
rect 16114 12764 16120 12776
rect 15335 12736 16120 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 13633 12699 13691 12705
rect 13633 12665 13645 12699
rect 13679 12665 13691 12699
rect 13633 12659 13691 12665
rect 13725 12699 13783 12705
rect 13725 12665 13737 12699
rect 13771 12696 13783 12699
rect 13998 12696 14004 12708
rect 13771 12668 14004 12696
rect 13771 12665 13783 12668
rect 13725 12659 13783 12665
rect 13998 12656 14004 12668
rect 14056 12656 14062 12708
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 1762 12628 1768 12640
rect 1627 12600 1768 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 1762 12588 1768 12600
rect 1820 12588 1826 12640
rect 3050 12628 3056 12640
rect 3011 12600 3056 12628
rect 3050 12588 3056 12600
rect 3108 12588 3114 12640
rect 4890 12588 4896 12640
rect 4948 12628 4954 12640
rect 5813 12631 5871 12637
rect 5813 12628 5825 12631
rect 4948 12600 5825 12628
rect 4948 12588 4954 12600
rect 5813 12597 5825 12600
rect 5859 12597 5871 12631
rect 5813 12591 5871 12597
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 8941 12631 8999 12637
rect 8941 12628 8953 12631
rect 8076 12600 8953 12628
rect 8076 12588 8082 12600
rect 8941 12597 8953 12600
rect 8987 12628 8999 12631
rect 9030 12628 9036 12640
rect 8987 12600 9036 12628
rect 8987 12597 8999 12600
rect 8941 12591 8999 12597
rect 9030 12588 9036 12600
rect 9088 12628 9094 12640
rect 9677 12631 9735 12637
rect 9677 12628 9689 12631
rect 9088 12600 9689 12628
rect 9088 12588 9094 12600
rect 9677 12597 9689 12600
rect 9723 12597 9735 12631
rect 9677 12591 9735 12597
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10505 12631 10563 12637
rect 10505 12628 10517 12631
rect 10008 12600 10517 12628
rect 10008 12588 10014 12600
rect 10505 12597 10517 12600
rect 10551 12628 10563 12631
rect 11238 12628 11244 12640
rect 10551 12600 11244 12628
rect 10551 12597 10563 12600
rect 10505 12591 10563 12597
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 15197 12631 15255 12637
rect 15197 12597 15209 12631
rect 15243 12628 15255 12631
rect 15470 12628 15476 12640
rect 15243 12600 15476 12628
rect 15243 12597 15255 12600
rect 15197 12591 15255 12597
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 15654 12588 15660 12640
rect 15712 12628 15718 12640
rect 15749 12631 15807 12637
rect 15749 12628 15761 12631
rect 15712 12600 15761 12628
rect 15712 12588 15718 12600
rect 15749 12597 15761 12600
rect 15795 12628 15807 12631
rect 16482 12628 16488 12640
rect 15795 12600 16488 12628
rect 15795 12597 15807 12600
rect 15749 12591 15807 12597
rect 16482 12588 16488 12600
rect 16540 12588 16546 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1394 12384 1400 12436
rect 1452 12424 1458 12436
rect 1857 12427 1915 12433
rect 1857 12424 1869 12427
rect 1452 12396 1869 12424
rect 1452 12384 1458 12396
rect 1857 12393 1869 12396
rect 1903 12393 1915 12427
rect 1857 12387 1915 12393
rect 1872 12288 1900 12387
rect 3050 12384 3056 12436
rect 3108 12424 3114 12436
rect 3421 12427 3479 12433
rect 3421 12424 3433 12427
rect 3108 12396 3433 12424
rect 3108 12384 3114 12396
rect 3421 12393 3433 12396
rect 3467 12393 3479 12427
rect 3878 12424 3884 12436
rect 3839 12396 3884 12424
rect 3421 12387 3479 12393
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 5353 12427 5411 12433
rect 5353 12393 5365 12427
rect 5399 12424 5411 12427
rect 5442 12424 5448 12436
rect 5399 12396 5448 12424
rect 5399 12393 5411 12396
rect 5353 12387 5411 12393
rect 5442 12384 5448 12396
rect 5500 12424 5506 12436
rect 6914 12424 6920 12436
rect 5500 12396 6920 12424
rect 5500 12384 5506 12396
rect 6914 12384 6920 12396
rect 6972 12384 6978 12436
rect 7466 12384 7472 12436
rect 7524 12424 7530 12436
rect 7745 12427 7803 12433
rect 7745 12424 7757 12427
rect 7524 12396 7757 12424
rect 7524 12384 7530 12396
rect 7745 12393 7757 12396
rect 7791 12393 7803 12427
rect 7745 12387 7803 12393
rect 11149 12427 11207 12433
rect 11149 12393 11161 12427
rect 11195 12424 11207 12427
rect 11698 12424 11704 12436
rect 11195 12396 11704 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12802 12424 12808 12436
rect 12492 12396 12808 12424
rect 12492 12384 12498 12396
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 14182 12424 14188 12436
rect 14143 12396 14188 12424
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 1946 12316 1952 12368
rect 2004 12356 2010 12368
rect 2777 12359 2835 12365
rect 2777 12356 2789 12359
rect 2004 12328 2789 12356
rect 2004 12316 2010 12328
rect 2777 12325 2789 12328
rect 2823 12325 2835 12359
rect 2958 12356 2964 12368
rect 2919 12328 2964 12356
rect 2777 12319 2835 12325
rect 2958 12316 2964 12328
rect 3016 12316 3022 12368
rect 4430 12316 4436 12368
rect 4488 12356 4494 12368
rect 4801 12359 4859 12365
rect 4801 12356 4813 12359
rect 4488 12328 4813 12356
rect 4488 12316 4494 12328
rect 4801 12325 4813 12328
rect 4847 12325 4859 12359
rect 5994 12356 6000 12368
rect 4801 12319 4859 12325
rect 5828 12328 6000 12356
rect 2222 12288 2228 12300
rect 1872 12260 2228 12288
rect 2222 12248 2228 12260
rect 2280 12288 2286 12300
rect 3053 12291 3111 12297
rect 3053 12288 3065 12291
rect 2280 12260 3065 12288
rect 2280 12248 2286 12260
rect 3053 12257 3065 12260
rect 3099 12257 3111 12291
rect 3053 12251 3111 12257
rect 3234 12248 3240 12300
rect 3292 12288 3298 12300
rect 5828 12297 5856 12328
rect 5994 12316 6000 12328
rect 6052 12316 6058 12368
rect 7098 12316 7104 12368
rect 7156 12356 7162 12368
rect 7926 12356 7932 12368
rect 7156 12328 7932 12356
rect 7156 12316 7162 12328
rect 7926 12316 7932 12328
rect 7984 12316 7990 12368
rect 9030 12316 9036 12368
rect 9088 12356 9094 12368
rect 10229 12359 10287 12365
rect 10229 12356 10241 12359
rect 9088 12328 10241 12356
rect 9088 12316 9094 12328
rect 10229 12325 10241 12328
rect 10275 12356 10287 12359
rect 11422 12356 11428 12368
rect 10275 12328 11428 12356
rect 10275 12325 10287 12328
rect 10229 12319 10287 12325
rect 11422 12316 11428 12328
rect 11480 12316 11486 12368
rect 11790 12356 11796 12368
rect 11751 12328 11796 12356
rect 11790 12316 11796 12328
rect 11848 12316 11854 12368
rect 13354 12356 13360 12368
rect 13267 12328 13360 12356
rect 13354 12316 13360 12328
rect 13412 12356 13418 12368
rect 13814 12356 13820 12368
rect 13412 12328 13820 12356
rect 13412 12316 13418 12328
rect 13814 12316 13820 12328
rect 13872 12316 13878 12368
rect 14826 12316 14832 12368
rect 14884 12356 14890 12368
rect 15841 12359 15899 12365
rect 15841 12356 15853 12359
rect 14884 12328 15853 12356
rect 14884 12316 14890 12328
rect 15841 12325 15853 12328
rect 15887 12325 15899 12359
rect 15841 12319 15899 12325
rect 4893 12291 4951 12297
rect 4893 12288 4905 12291
rect 3292 12260 4905 12288
rect 3292 12248 3298 12260
rect 4893 12257 4905 12260
rect 4939 12257 4951 12291
rect 4893 12251 4951 12257
rect 5813 12291 5871 12297
rect 5813 12257 5825 12291
rect 5859 12257 5871 12291
rect 6080 12291 6138 12297
rect 6080 12288 6092 12291
rect 5813 12251 5871 12257
rect 5920 12260 6092 12288
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 3016 12192 4721 12220
rect 3016 12180 3022 12192
rect 4709 12189 4721 12192
rect 4755 12220 4767 12223
rect 4798 12220 4804 12232
rect 4755 12192 4804 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12220 5779 12223
rect 5920 12220 5948 12260
rect 6080 12257 6092 12260
rect 6126 12288 6138 12291
rect 6362 12288 6368 12300
rect 6126 12260 6368 12288
rect 6126 12257 6138 12260
rect 6080 12251 6138 12257
rect 6362 12248 6368 12260
rect 6420 12288 6426 12300
rect 8110 12288 8116 12300
rect 6420 12260 8116 12288
rect 6420 12248 6426 12260
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 10042 12288 10048 12300
rect 10003 12260 10048 12288
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 10686 12288 10692 12300
rect 10647 12260 10692 12288
rect 10686 12248 10692 12260
rect 10744 12288 10750 12300
rect 11054 12288 11060 12300
rect 10744 12260 11060 12288
rect 10744 12248 10750 12260
rect 11054 12248 11060 12260
rect 11112 12288 11118 12300
rect 11609 12291 11667 12297
rect 11609 12288 11621 12291
rect 11112 12260 11621 12288
rect 11112 12248 11118 12260
rect 11609 12257 11621 12260
rect 11655 12257 11667 12291
rect 13170 12288 13176 12300
rect 13131 12260 13176 12288
rect 11609 12251 11667 12257
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 13909 12291 13967 12297
rect 13909 12257 13921 12291
rect 13955 12288 13967 12291
rect 13998 12288 14004 12300
rect 13955 12260 14004 12288
rect 13955 12257 13967 12260
rect 13909 12251 13967 12257
rect 13998 12248 14004 12260
rect 14056 12288 14062 12300
rect 15562 12288 15568 12300
rect 14056 12260 15568 12288
rect 14056 12248 14062 12260
rect 15562 12248 15568 12260
rect 15620 12288 15626 12300
rect 15933 12291 15991 12297
rect 15933 12288 15945 12291
rect 15620 12260 15945 12288
rect 15620 12248 15626 12260
rect 15933 12257 15945 12260
rect 15979 12288 15991 12291
rect 16758 12288 16764 12300
rect 15979 12260 16764 12288
rect 15979 12257 15991 12260
rect 15933 12251 15991 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 19521 12291 19579 12297
rect 19521 12288 19533 12291
rect 19484 12260 19533 12288
rect 19484 12248 19490 12260
rect 19521 12257 19533 12260
rect 19567 12257 19579 12291
rect 19521 12251 19579 12257
rect 5767 12192 5948 12220
rect 8389 12223 8447 12229
rect 5767 12189 5779 12192
rect 5721 12183 5779 12189
rect 8389 12189 8401 12223
rect 8435 12220 8447 12223
rect 8662 12220 8668 12232
rect 8435 12192 8668 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 9582 12220 9588 12232
rect 9180 12192 9588 12220
rect 9180 12180 9186 12192
rect 9582 12180 9588 12192
rect 9640 12180 9646 12232
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 11885 12223 11943 12229
rect 11885 12189 11897 12223
rect 11931 12220 11943 12223
rect 13262 12220 13268 12232
rect 11931 12192 13268 12220
rect 11931 12189 11943 12192
rect 11885 12183 11943 12189
rect 2225 12155 2283 12161
rect 2225 12121 2237 12155
rect 2271 12152 2283 12155
rect 2774 12152 2780 12164
rect 2271 12124 2780 12152
rect 2271 12121 2283 12124
rect 2225 12115 2283 12121
rect 2774 12112 2780 12124
rect 2832 12112 2838 12164
rect 4338 12152 4344 12164
rect 4299 12124 4344 12152
rect 4338 12112 4344 12124
rect 4396 12112 4402 12164
rect 8294 12112 8300 12164
rect 8352 12152 8358 12164
rect 9214 12152 9220 12164
rect 8352 12124 9220 12152
rect 8352 12112 8358 12124
rect 9214 12112 9220 12124
rect 9272 12152 9278 12164
rect 10336 12152 10364 12183
rect 10778 12152 10784 12164
rect 9272 12124 10784 12152
rect 9272 12112 9278 12124
rect 10778 12112 10784 12124
rect 10836 12152 10842 12164
rect 11900 12152 11928 12183
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 13446 12220 13452 12232
rect 13407 12192 13452 12220
rect 13446 12180 13452 12192
rect 13504 12180 13510 12232
rect 15838 12220 15844 12232
rect 15799 12192 15844 12220
rect 15838 12180 15844 12192
rect 15896 12180 15902 12232
rect 12894 12152 12900 12164
rect 10836 12124 11928 12152
rect 12855 12124 12900 12152
rect 10836 12112 10842 12124
rect 12894 12112 12900 12124
rect 12952 12112 12958 12164
rect 13354 12112 13360 12164
rect 13412 12152 13418 12164
rect 15010 12152 15016 12164
rect 13412 12124 15016 12152
rect 13412 12112 13418 12124
rect 15010 12112 15016 12124
rect 15068 12112 15074 12164
rect 15381 12155 15439 12161
rect 15381 12121 15393 12155
rect 15427 12152 15439 12155
rect 15470 12152 15476 12164
rect 15427 12124 15476 12152
rect 15427 12121 15439 12124
rect 15381 12115 15439 12121
rect 15470 12112 15476 12124
rect 15528 12112 15534 12164
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 2501 12087 2559 12093
rect 2501 12084 2513 12087
rect 2096 12056 2513 12084
rect 2096 12044 2102 12056
rect 2501 12053 2513 12056
rect 2547 12053 2559 12087
rect 2501 12047 2559 12053
rect 2866 12044 2872 12096
rect 2924 12084 2930 12096
rect 3142 12084 3148 12096
rect 2924 12056 3148 12084
rect 2924 12044 2930 12056
rect 3142 12044 3148 12056
rect 3200 12044 3206 12096
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 7193 12087 7251 12093
rect 7193 12084 7205 12087
rect 6972 12056 7205 12084
rect 6972 12044 6978 12056
rect 7193 12053 7205 12056
rect 7239 12053 7251 12087
rect 7193 12047 7251 12053
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 8113 12087 8171 12093
rect 8113 12084 8125 12087
rect 8076 12056 8125 12084
rect 8076 12044 8082 12056
rect 8113 12053 8125 12056
rect 8159 12053 8171 12087
rect 8113 12047 8171 12053
rect 8570 12044 8576 12096
rect 8628 12084 8634 12096
rect 9125 12087 9183 12093
rect 9125 12084 9137 12087
rect 8628 12056 9137 12084
rect 8628 12044 8634 12056
rect 9125 12053 9137 12056
rect 9171 12084 9183 12087
rect 9398 12084 9404 12096
rect 9171 12056 9404 12084
rect 9171 12053 9183 12056
rect 9125 12047 9183 12053
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 9582 12044 9588 12096
rect 9640 12084 9646 12096
rect 9769 12087 9827 12093
rect 9769 12084 9781 12087
rect 9640 12056 9781 12084
rect 9640 12044 9646 12056
rect 9769 12053 9781 12056
rect 9815 12053 9827 12087
rect 9769 12047 9827 12053
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 11333 12087 11391 12093
rect 11333 12084 11345 12087
rect 11204 12056 11345 12084
rect 11204 12044 11210 12056
rect 11333 12053 11345 12056
rect 11379 12053 11391 12087
rect 11333 12047 11391 12053
rect 12529 12087 12587 12093
rect 12529 12053 12541 12087
rect 12575 12084 12587 12087
rect 12618 12084 12624 12096
rect 12575 12056 12624 12084
rect 12575 12053 12587 12056
rect 12529 12047 12587 12053
rect 12618 12044 12624 12056
rect 12676 12084 12682 12096
rect 12986 12084 12992 12096
rect 12676 12056 12992 12084
rect 12676 12044 12682 12056
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 14737 12087 14795 12093
rect 14737 12053 14749 12087
rect 14783 12084 14795 12087
rect 14826 12084 14832 12096
rect 14783 12056 14832 12084
rect 14783 12053 14795 12056
rect 14737 12047 14795 12053
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 15105 12087 15163 12093
rect 15105 12053 15117 12087
rect 15151 12084 15163 12087
rect 15286 12084 15292 12096
rect 15151 12056 15292 12084
rect 15151 12053 15163 12056
rect 15105 12047 15163 12053
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 19705 12087 19763 12093
rect 19705 12053 19717 12087
rect 19751 12084 19763 12087
rect 20622 12084 20628 12096
rect 19751 12056 20628 12084
rect 19751 12053 19763 12056
rect 19705 12047 19763 12053
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1946 11880 1952 11892
rect 1907 11852 1952 11880
rect 1946 11840 1952 11852
rect 2004 11840 2010 11892
rect 4522 11840 4528 11892
rect 4580 11880 4586 11892
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 4580 11852 5273 11880
rect 4580 11840 4586 11852
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 5261 11843 5319 11849
rect 5994 11840 6000 11892
rect 6052 11880 6058 11892
rect 6181 11883 6239 11889
rect 6181 11880 6193 11883
rect 6052 11852 6193 11880
rect 6052 11840 6058 11852
rect 6181 11849 6193 11852
rect 6227 11880 6239 11883
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 6227 11852 6561 11880
rect 6227 11849 6239 11852
rect 6181 11843 6239 11849
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 6549 11843 6607 11849
rect 4798 11812 4804 11824
rect 4759 11784 4804 11812
rect 4798 11772 4804 11784
rect 4856 11772 4862 11824
rect 6564 11744 6592 11843
rect 8110 11840 8116 11892
rect 8168 11880 8174 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 8168 11852 8217 11880
rect 8168 11840 8174 11852
rect 8205 11849 8217 11852
rect 8251 11849 8263 11883
rect 8205 11843 8263 11849
rect 9125 11883 9183 11889
rect 9125 11849 9137 11883
rect 9171 11880 9183 11883
rect 9490 11880 9496 11892
rect 9171 11852 9496 11880
rect 9171 11849 9183 11852
rect 9125 11843 9183 11849
rect 9490 11840 9496 11852
rect 9548 11880 9554 11892
rect 10042 11880 10048 11892
rect 9548 11852 10048 11880
rect 9548 11840 9554 11852
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10686 11840 10692 11892
rect 10744 11880 10750 11892
rect 10965 11883 11023 11889
rect 10965 11880 10977 11883
rect 10744 11852 10977 11880
rect 10744 11840 10750 11852
rect 10965 11849 10977 11852
rect 11011 11849 11023 11883
rect 10965 11843 11023 11849
rect 11701 11883 11759 11889
rect 11701 11849 11713 11883
rect 11747 11880 11759 11883
rect 11790 11880 11796 11892
rect 11747 11852 11796 11880
rect 11747 11849 11759 11852
rect 11701 11843 11759 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 13446 11880 13452 11892
rect 13407 11852 13452 11880
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 13814 11880 13820 11892
rect 13775 11852 13820 11880
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 15289 11883 15347 11889
rect 15289 11849 15301 11883
rect 15335 11880 15347 11883
rect 15746 11880 15752 11892
rect 15335 11852 15752 11880
rect 15335 11849 15347 11852
rect 15289 11843 15347 11849
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 16758 11880 16764 11892
rect 16719 11852 16764 11880
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 19426 11840 19432 11892
rect 19484 11880 19490 11892
rect 19521 11883 19579 11889
rect 19521 11880 19533 11883
rect 19484 11852 19533 11880
rect 19484 11840 19490 11852
rect 19521 11849 19533 11852
rect 19567 11849 19579 11883
rect 19521 11843 19579 11849
rect 9030 11772 9036 11824
rect 9088 11812 9094 11824
rect 9401 11815 9459 11821
rect 9401 11812 9413 11815
rect 9088 11784 9413 11812
rect 9088 11772 9094 11784
rect 9401 11781 9413 11784
rect 9447 11781 9459 11815
rect 9674 11812 9680 11824
rect 9635 11784 9680 11812
rect 9401 11775 9459 11781
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 12526 11812 12532 11824
rect 12487 11784 12532 11812
rect 12526 11772 12532 11784
rect 12584 11772 12590 11824
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6564 11716 6837 11744
rect 6825 11713 6837 11716
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10229 11747 10287 11753
rect 10229 11744 10241 11747
rect 10100 11716 10241 11744
rect 10100 11704 10106 11716
rect 10229 11713 10241 11716
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 11296 11716 12173 11744
rect 11296 11704 11302 11716
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 2409 11679 2467 11685
rect 2409 11645 2421 11679
rect 2455 11676 2467 11679
rect 3418 11676 3424 11688
rect 2455 11648 3424 11676
rect 2455 11645 2467 11648
rect 2409 11639 2467 11645
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 3602 11636 3608 11688
rect 3660 11676 3666 11688
rect 3786 11676 3792 11688
rect 3660 11648 3792 11676
rect 3660 11636 3666 11648
rect 3786 11636 3792 11648
rect 3844 11636 3850 11688
rect 5166 11636 5172 11688
rect 5224 11676 5230 11688
rect 5813 11679 5871 11685
rect 5813 11676 5825 11679
rect 5224 11648 5825 11676
rect 5224 11636 5230 11648
rect 5813 11645 5825 11648
rect 5859 11676 5871 11679
rect 6914 11676 6920 11688
rect 5859 11648 6920 11676
rect 5859 11645 5871 11648
rect 5813 11639 5871 11645
rect 6914 11636 6920 11648
rect 6972 11636 6978 11688
rect 7092 11679 7150 11685
rect 7092 11645 7104 11679
rect 7138 11676 7150 11679
rect 8202 11676 8208 11688
rect 7138 11648 8208 11676
rect 7138 11645 7150 11648
rect 7092 11639 7150 11645
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 9953 11679 10011 11685
rect 9953 11645 9965 11679
rect 9999 11676 10011 11679
rect 12176 11676 12204 11707
rect 12805 11679 12863 11685
rect 12805 11676 12817 11679
rect 9999 11648 10732 11676
rect 12176 11648 12817 11676
rect 9999 11645 10011 11648
rect 9953 11639 10011 11645
rect 2222 11568 2228 11620
rect 2280 11608 2286 11620
rect 2654 11611 2712 11617
rect 2654 11608 2666 11611
rect 2280 11580 2666 11608
rect 2280 11568 2286 11580
rect 2654 11577 2666 11580
rect 2700 11577 2712 11611
rect 5534 11608 5540 11620
rect 5495 11580 5540 11608
rect 2654 11571 2712 11577
rect 5534 11568 5540 11580
rect 5592 11568 5598 11620
rect 10134 11608 10140 11620
rect 10095 11580 10140 11608
rect 10134 11568 10140 11580
rect 10192 11568 10198 11620
rect 10704 11617 10732 11648
rect 12805 11645 12817 11648
rect 12851 11645 12863 11679
rect 12805 11639 12863 11645
rect 14001 11679 14059 11685
rect 14001 11645 14013 11679
rect 14047 11676 14059 11679
rect 14182 11676 14188 11688
rect 14047 11648 14188 11676
rect 14047 11645 14059 11648
rect 14001 11639 14059 11645
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11676 14979 11679
rect 15194 11676 15200 11688
rect 14967 11648 15200 11676
rect 14967 11645 14979 11648
rect 14921 11639 14979 11645
rect 15194 11636 15200 11648
rect 15252 11676 15258 11688
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 15252 11648 15393 11676
rect 15252 11636 15258 11648
rect 15381 11645 15393 11648
rect 15427 11645 15439 11679
rect 15381 11639 15439 11645
rect 10689 11611 10747 11617
rect 10689 11577 10701 11611
rect 10735 11608 10747 11611
rect 11149 11611 11207 11617
rect 11149 11608 11161 11611
rect 10735 11580 11161 11608
rect 10735 11577 10747 11580
rect 10689 11571 10747 11577
rect 11149 11577 11161 11580
rect 11195 11577 11207 11611
rect 12986 11608 12992 11620
rect 12947 11580 12992 11608
rect 11149 11571 11207 11577
rect 12986 11568 12992 11580
rect 13044 11568 13050 11620
rect 13081 11611 13139 11617
rect 13081 11577 13093 11611
rect 13127 11608 13139 11611
rect 13262 11608 13268 11620
rect 13127 11580 13268 11608
rect 13127 11577 13139 11580
rect 13081 11571 13139 11577
rect 13262 11568 13268 11580
rect 13320 11568 13326 11620
rect 14274 11608 14280 11620
rect 14235 11580 14280 11608
rect 14274 11568 14280 11580
rect 14332 11568 14338 11620
rect 15286 11568 15292 11620
rect 15344 11608 15350 11620
rect 15626 11611 15684 11617
rect 15626 11608 15638 11611
rect 15344 11580 15638 11608
rect 15344 11568 15350 11580
rect 15626 11577 15638 11580
rect 15672 11577 15684 11611
rect 15626 11571 15684 11577
rect 1394 11540 1400 11552
rect 1355 11512 1400 11540
rect 1394 11500 1400 11512
rect 1452 11500 1458 11552
rect 2317 11543 2375 11549
rect 2317 11509 2329 11543
rect 2363 11540 2375 11543
rect 3050 11540 3056 11552
rect 2363 11512 3056 11540
rect 2363 11509 2375 11512
rect 2317 11503 2375 11509
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 3786 11540 3792 11552
rect 3747 11512 3792 11540
rect 3786 11500 3792 11512
rect 3844 11500 3850 11552
rect 4338 11540 4344 11552
rect 4299 11512 4344 11540
rect 4338 11500 4344 11512
rect 4396 11500 4402 11552
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 5721 11543 5779 11549
rect 5721 11540 5733 11543
rect 5500 11512 5733 11540
rect 5500 11500 5506 11512
rect 5721 11509 5733 11512
rect 5767 11509 5779 11543
rect 5721 11503 5779 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 2222 11336 2228 11348
rect 2179 11308 2228 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 3510 11336 3516 11348
rect 2832 11308 3516 11336
rect 2832 11296 2838 11308
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 5534 11336 5540 11348
rect 5495 11308 5540 11336
rect 5534 11296 5540 11308
rect 5592 11336 5598 11348
rect 5795 11339 5853 11345
rect 5795 11336 5807 11339
rect 5592 11308 5807 11336
rect 5592 11296 5598 11308
rect 5795 11305 5807 11308
rect 5841 11305 5853 11339
rect 5795 11299 5853 11305
rect 6273 11339 6331 11345
rect 6273 11305 6285 11339
rect 6319 11336 6331 11339
rect 6454 11336 6460 11348
rect 6319 11308 6460 11336
rect 6319 11305 6331 11308
rect 6273 11299 6331 11305
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 7837 11339 7895 11345
rect 7837 11305 7849 11339
rect 7883 11336 7895 11339
rect 8202 11336 8208 11348
rect 7883 11308 8208 11336
rect 7883 11305 7895 11308
rect 7837 11299 7895 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 9214 11296 9220 11348
rect 9272 11336 9278 11348
rect 9401 11339 9459 11345
rect 9401 11336 9413 11339
rect 9272 11308 9413 11336
rect 9272 11296 9278 11308
rect 9401 11305 9413 11308
rect 9447 11305 9459 11339
rect 9401 11299 9459 11305
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10689 11339 10747 11345
rect 10689 11336 10701 11339
rect 10192 11308 10701 11336
rect 10192 11296 10198 11308
rect 10689 11305 10701 11308
rect 10735 11305 10747 11339
rect 10689 11299 10747 11305
rect 10778 11296 10784 11348
rect 10836 11336 10842 11348
rect 11057 11339 11115 11345
rect 11057 11336 11069 11339
rect 10836 11308 11069 11336
rect 10836 11296 10842 11308
rect 11057 11305 11069 11308
rect 11103 11305 11115 11339
rect 11057 11299 11115 11305
rect 13170 11296 13176 11348
rect 13228 11336 13234 11348
rect 13541 11339 13599 11345
rect 13541 11336 13553 11339
rect 13228 11308 13553 11336
rect 13228 11296 13234 11308
rect 13541 11305 13553 11308
rect 13587 11305 13599 11339
rect 13541 11299 13599 11305
rect 15105 11339 15163 11345
rect 15105 11305 15117 11339
rect 15151 11336 15163 11339
rect 15286 11336 15292 11348
rect 15151 11308 15292 11336
rect 15151 11305 15163 11308
rect 15105 11299 15163 11305
rect 15286 11296 15292 11308
rect 15344 11336 15350 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 15344 11308 16681 11336
rect 15344 11296 15350 11308
rect 16669 11305 16681 11308
rect 16715 11305 16727 11339
rect 16669 11299 16727 11305
rect 1394 11228 1400 11280
rect 1452 11268 1458 11280
rect 2498 11268 2504 11280
rect 1452 11240 2504 11268
rect 1452 11228 1458 11240
rect 2498 11228 2504 11240
rect 2556 11268 2562 11280
rect 2593 11271 2651 11277
rect 2593 11268 2605 11271
rect 2556 11240 2605 11268
rect 2556 11228 2562 11240
rect 2593 11237 2605 11240
rect 2639 11237 2651 11271
rect 2593 11231 2651 11237
rect 2869 11271 2927 11277
rect 2869 11237 2881 11271
rect 2915 11268 2927 11271
rect 3326 11268 3332 11280
rect 2915 11240 3332 11268
rect 2915 11237 2927 11240
rect 2869 11231 2927 11237
rect 3326 11228 3332 11240
rect 3384 11268 3390 11280
rect 3786 11268 3792 11280
rect 3384 11240 3792 11268
rect 3384 11228 3390 11240
rect 3786 11228 3792 11240
rect 3844 11228 3850 11280
rect 4614 11228 4620 11280
rect 4672 11268 4678 11280
rect 4709 11271 4767 11277
rect 4709 11268 4721 11271
rect 4672 11240 4721 11268
rect 4672 11228 4678 11240
rect 4709 11237 4721 11240
rect 4755 11237 4767 11271
rect 4709 11231 4767 11237
rect 4798 11228 4804 11280
rect 4856 11268 4862 11280
rect 4856 11240 4901 11268
rect 4856 11228 4862 11240
rect 6362 11228 6368 11280
rect 6420 11268 6426 11280
rect 8573 11271 8631 11277
rect 6420 11240 6465 11268
rect 6420 11228 6426 11240
rect 8573 11237 8585 11271
rect 8619 11268 8631 11271
rect 9030 11268 9036 11280
rect 8619 11240 9036 11268
rect 8619 11237 8631 11240
rect 8573 11231 8631 11237
rect 9030 11228 9036 11240
rect 9088 11228 9094 11280
rect 9674 11228 9680 11280
rect 9732 11268 9738 11280
rect 10045 11271 10103 11277
rect 10045 11268 10057 11271
rect 9732 11240 10057 11268
rect 9732 11228 9738 11240
rect 10045 11237 10057 11240
rect 10091 11237 10103 11271
rect 10045 11231 10103 11237
rect 10229 11271 10287 11277
rect 10229 11237 10241 11271
rect 10275 11237 10287 11271
rect 10229 11231 10287 11237
rect 14737 11271 14795 11277
rect 14737 11237 14749 11271
rect 14783 11268 14795 11271
rect 15654 11268 15660 11280
rect 14783 11240 15660 11268
rect 14783 11237 14795 11240
rect 14737 11231 14795 11237
rect 2222 11160 2228 11212
rect 2280 11200 2286 11212
rect 3142 11200 3148 11212
rect 2280 11172 3148 11200
rect 2280 11160 2286 11172
rect 3142 11160 3148 11172
rect 3200 11160 3206 11212
rect 3234 11160 3240 11212
rect 3292 11200 3298 11212
rect 3881 11203 3939 11209
rect 3881 11200 3893 11203
rect 3292 11172 3893 11200
rect 3292 11160 3298 11172
rect 3881 11169 3893 11172
rect 3927 11200 3939 11203
rect 5166 11200 5172 11212
rect 3927 11172 5172 11200
rect 3927 11169 3939 11172
rect 3881 11163 3939 11169
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 5442 11160 5448 11212
rect 5500 11200 5506 11212
rect 6380 11200 6408 11228
rect 5500 11172 6408 11200
rect 8389 11203 8447 11209
rect 5500 11160 5506 11172
rect 8389 11169 8401 11203
rect 8435 11200 8447 11203
rect 9582 11200 9588 11212
rect 8435 11172 9588 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 9582 11160 9588 11172
rect 9640 11160 9646 11212
rect 10244 11200 10272 11231
rect 15654 11228 15660 11240
rect 15712 11228 15718 11280
rect 11054 11200 11060 11212
rect 10244 11172 11060 11200
rect 3329 11135 3387 11141
rect 1964 11104 2636 11132
rect 1964 11008 1992 11104
rect 2317 11067 2375 11073
rect 2317 11033 2329 11067
rect 2363 11064 2375 11067
rect 2608 11064 2636 11104
rect 3329 11101 3341 11135
rect 3375 11132 3387 11135
rect 3418 11132 3424 11144
rect 3375 11104 3424 11132
rect 3375 11101 3387 11104
rect 3329 11095 3387 11101
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 4709 11095 4767 11101
rect 5092 11104 6193 11132
rect 4249 11067 4307 11073
rect 4249 11064 4261 11067
rect 2363 11036 2544 11064
rect 2608 11036 4261 11064
rect 2363 11033 2375 11036
rect 2317 11027 2375 11033
rect 1673 10999 1731 11005
rect 1673 10965 1685 10999
rect 1719 10996 1731 10999
rect 1946 10996 1952 11008
rect 1719 10968 1952 10996
rect 1719 10965 1731 10968
rect 1673 10959 1731 10965
rect 1946 10956 1952 10968
rect 2004 10956 2010 11008
rect 2516 10996 2544 11036
rect 4249 11033 4261 11036
rect 4295 11033 4307 11067
rect 4724 11064 4752 11095
rect 5092 11076 5120 11104
rect 6181 11101 6193 11104
rect 6227 11101 6239 11135
rect 8570 11132 8576 11144
rect 6181 11095 6239 11101
rect 7024 11104 8576 11132
rect 5074 11064 5080 11076
rect 4724 11036 5080 11064
rect 4249 11027 4307 11033
rect 5074 11024 5080 11036
rect 5132 11024 5138 11076
rect 5350 11024 5356 11076
rect 5408 11064 5414 11076
rect 6914 11064 6920 11076
rect 5408 11036 6920 11064
rect 5408 11024 5414 11036
rect 6914 11024 6920 11036
rect 6972 11064 6978 11076
rect 7024 11073 7052 11104
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 8665 11135 8723 11141
rect 8665 11101 8677 11135
rect 8711 11132 8723 11135
rect 8849 11135 8907 11141
rect 8849 11132 8861 11135
rect 8711 11104 8861 11132
rect 8711 11101 8723 11104
rect 8665 11095 8723 11101
rect 8849 11101 8861 11104
rect 8895 11101 8907 11135
rect 10244 11132 10272 11172
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 11330 11160 11336 11212
rect 11388 11200 11394 11212
rect 11497 11203 11555 11209
rect 11497 11200 11509 11203
rect 11388 11172 11509 11200
rect 11388 11160 11394 11172
rect 11497 11169 11509 11172
rect 11543 11169 11555 11203
rect 13722 11200 13728 11212
rect 13683 11172 13728 11200
rect 11497 11163 11555 11169
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 15545 11203 15603 11209
rect 15545 11200 15557 11203
rect 14700 11172 15557 11200
rect 14700 11160 14706 11172
rect 15545 11169 15557 11172
rect 15591 11169 15603 11203
rect 15545 11163 15603 11169
rect 8849 11095 8907 11101
rect 9048 11104 10272 11132
rect 10321 11135 10379 11141
rect 7009 11067 7067 11073
rect 7009 11064 7021 11067
rect 6972 11036 7021 11064
rect 6972 11024 6978 11036
rect 7009 11033 7021 11036
rect 7055 11033 7067 11067
rect 7009 11027 7067 11033
rect 8113 11067 8171 11073
rect 8113 11033 8125 11067
rect 8159 11064 8171 11067
rect 9048 11064 9076 11104
rect 10321 11101 10333 11135
rect 10367 11132 10379 11135
rect 10778 11132 10784 11144
rect 10367 11104 10784 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 11238 11132 11244 11144
rect 11199 11104 11244 11132
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 13998 11132 14004 11144
rect 13959 11104 14004 11132
rect 13998 11092 14004 11104
rect 14056 11092 14062 11144
rect 15194 11092 15200 11144
rect 15252 11132 15258 11144
rect 15289 11135 15347 11141
rect 15289 11132 15301 11135
rect 15252 11104 15301 11132
rect 15252 11092 15258 11104
rect 15289 11101 15301 11104
rect 15335 11101 15347 11135
rect 15289 11095 15347 11101
rect 9766 11064 9772 11076
rect 8159 11036 9076 11064
rect 9727 11036 9772 11064
rect 8159 11033 8171 11036
rect 8113 11027 8171 11033
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 13262 11064 13268 11076
rect 13223 11036 13268 11064
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 2866 10996 2872 11008
rect 2516 10968 2872 10996
rect 2866 10956 2872 10968
rect 2924 10956 2930 11008
rect 4614 10956 4620 11008
rect 4672 10996 4678 11008
rect 5994 10996 6000 11008
rect 4672 10968 6000 10996
rect 4672 10956 4678 10968
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 7374 10996 7380 11008
rect 7335 10968 7380 10996
rect 7374 10956 7380 10968
rect 7432 10956 7438 11008
rect 8754 10956 8760 11008
rect 8812 10996 8818 11008
rect 8849 10999 8907 11005
rect 8849 10996 8861 10999
rect 8812 10968 8861 10996
rect 8812 10956 8818 10968
rect 8849 10965 8861 10968
rect 8895 10996 8907 10999
rect 9125 10999 9183 11005
rect 9125 10996 9137 10999
rect 8895 10968 9137 10996
rect 8895 10965 8907 10968
rect 8849 10959 8907 10965
rect 9125 10965 9137 10968
rect 9171 10996 9183 10999
rect 10042 10996 10048 11008
rect 9171 10968 10048 10996
rect 9171 10965 9183 10968
rect 9125 10959 9183 10965
rect 10042 10956 10048 10968
rect 10100 10956 10106 11008
rect 12618 10996 12624 11008
rect 12579 10968 12624 10996
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 15304 10996 15332 11095
rect 16482 10996 16488 11008
rect 15304 10968 16488 10996
rect 16482 10956 16488 10968
rect 16540 10956 16546 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2498 10792 2504 10804
rect 2459 10764 2504 10792
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 3418 10792 3424 10804
rect 2915 10764 3424 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 1581 10727 1639 10733
rect 1581 10693 1593 10727
rect 1627 10724 1639 10727
rect 2958 10724 2964 10736
rect 1627 10696 2964 10724
rect 1627 10693 1639 10696
rect 1581 10687 1639 10693
rect 2958 10684 2964 10696
rect 3016 10684 3022 10736
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 3068 10665 3096 10764
rect 3418 10752 3424 10764
rect 3476 10752 3482 10804
rect 5442 10792 5448 10804
rect 5403 10764 5448 10792
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 6181 10795 6239 10801
rect 6181 10761 6193 10795
rect 6227 10792 6239 10795
rect 6454 10792 6460 10804
rect 6227 10764 6460 10792
rect 6227 10761 6239 10764
rect 6181 10755 6239 10761
rect 6454 10752 6460 10764
rect 6512 10752 6518 10804
rect 7101 10795 7159 10801
rect 7101 10761 7113 10795
rect 7147 10792 7159 10795
rect 8938 10792 8944 10804
rect 7147 10764 8944 10792
rect 7147 10761 7159 10764
rect 7101 10755 7159 10761
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 9953 10795 10011 10801
rect 9953 10761 9965 10795
rect 9999 10792 10011 10795
rect 10042 10792 10048 10804
rect 9999 10764 10048 10792
rect 9999 10761 10011 10764
rect 9953 10755 10011 10761
rect 10042 10752 10048 10764
rect 10100 10792 10106 10804
rect 11057 10795 11115 10801
rect 11057 10792 11069 10795
rect 10100 10764 11069 10792
rect 10100 10752 10106 10764
rect 11057 10761 11069 10764
rect 11103 10792 11115 10795
rect 11330 10792 11336 10804
rect 11103 10764 11336 10792
rect 11103 10761 11115 10764
rect 11057 10755 11115 10761
rect 11330 10752 11336 10764
rect 11388 10752 11394 10804
rect 13170 10752 13176 10804
rect 13228 10792 13234 10804
rect 13909 10795 13967 10801
rect 13909 10792 13921 10795
rect 13228 10764 13921 10792
rect 13228 10752 13234 10764
rect 13909 10761 13921 10764
rect 13955 10792 13967 10795
rect 14553 10795 14611 10801
rect 14553 10792 14565 10795
rect 13955 10764 14565 10792
rect 13955 10761 13967 10764
rect 13909 10755 13967 10761
rect 14553 10761 14565 10764
rect 14599 10792 14611 10795
rect 14642 10792 14648 10804
rect 14599 10764 14648 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 14826 10752 14832 10804
rect 14884 10792 14890 10804
rect 15105 10795 15163 10801
rect 15105 10792 15117 10795
rect 14884 10764 15117 10792
rect 14884 10752 14890 10764
rect 15105 10761 15117 10764
rect 15151 10761 15163 10795
rect 15105 10755 15163 10761
rect 8113 10727 8171 10733
rect 8113 10693 8125 10727
rect 8159 10724 8171 10727
rect 8294 10724 8300 10736
rect 8159 10696 8300 10724
rect 8159 10693 8171 10696
rect 8113 10687 8171 10693
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10625 3111 10659
rect 7650 10656 7656 10668
rect 7563 10628 7656 10656
rect 3053 10619 3111 10625
rect 7650 10616 7656 10628
rect 7708 10656 7714 10668
rect 8128 10656 8156 10687
rect 8294 10684 8300 10696
rect 8352 10684 8358 10736
rect 12437 10659 12495 10665
rect 7708 10628 8708 10656
rect 7708 10616 7714 10628
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10588 2191 10591
rect 2222 10588 2228 10600
rect 2179 10560 2228 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 2222 10548 2228 10560
rect 2280 10588 2286 10600
rect 3326 10597 3332 10600
rect 3320 10588 3332 10597
rect 2280 10560 3332 10588
rect 2280 10548 2286 10560
rect 3320 10551 3332 10560
rect 3326 10548 3332 10551
rect 3384 10548 3390 10600
rect 5350 10588 5356 10600
rect 3436 10560 5356 10588
rect 1946 10480 1952 10532
rect 2004 10520 2010 10532
rect 2041 10523 2099 10529
rect 2041 10520 2053 10523
rect 2004 10492 2053 10520
rect 2004 10480 2010 10492
rect 2041 10489 2053 10492
rect 2087 10489 2099 10523
rect 2041 10483 2099 10489
rect 3436 10464 3464 10560
rect 5350 10548 5356 10560
rect 5408 10548 5414 10600
rect 5534 10588 5540 10600
rect 5495 10560 5540 10588
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 7282 10548 7288 10600
rect 7340 10588 7346 10600
rect 7377 10591 7435 10597
rect 7377 10588 7389 10591
rect 7340 10560 7389 10588
rect 7340 10548 7346 10560
rect 7377 10557 7389 10560
rect 7423 10557 7435 10591
rect 7377 10551 7435 10557
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8352 10560 8585 10588
rect 8352 10548 8358 10560
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 8680 10588 8708 10628
rect 12437 10625 12449 10659
rect 12483 10656 12495 10659
rect 12529 10659 12587 10665
rect 12529 10656 12541 10659
rect 12483 10628 12541 10656
rect 12483 10625 12495 10628
rect 12437 10619 12495 10625
rect 12529 10625 12541 10628
rect 12575 10625 12587 10659
rect 12529 10619 12587 10625
rect 15286 10616 15292 10668
rect 15344 10656 15350 10668
rect 15657 10659 15715 10665
rect 15657 10656 15669 10659
rect 15344 10628 15669 10656
rect 15344 10616 15350 10628
rect 15657 10625 15669 10628
rect 15703 10625 15715 10659
rect 15657 10619 15715 10625
rect 8829 10591 8887 10597
rect 8829 10588 8841 10591
rect 8680 10560 8841 10588
rect 8573 10551 8631 10557
rect 8829 10557 8841 10560
rect 8875 10557 8887 10591
rect 8829 10551 8887 10557
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 12785 10591 12843 10597
rect 12785 10588 12797 10591
rect 12676 10560 12797 10588
rect 12676 10548 12682 10560
rect 12785 10557 12797 10560
rect 12831 10557 12843 10591
rect 16574 10588 16580 10600
rect 16535 10560 16580 10588
rect 12785 10551 12843 10557
rect 16574 10548 16580 10560
rect 16632 10588 16638 10600
rect 17313 10591 17371 10597
rect 17313 10588 17325 10591
rect 16632 10560 17325 10588
rect 16632 10548 16638 10560
rect 17313 10557 17325 10560
rect 17359 10557 17371 10591
rect 17313 10551 17371 10557
rect 6457 10523 6515 10529
rect 6457 10520 6469 10523
rect 5092 10492 6469 10520
rect 5092 10464 5120 10492
rect 6457 10489 6469 10492
rect 6503 10489 6515 10523
rect 6457 10483 6515 10489
rect 11238 10480 11244 10532
rect 11296 10520 11302 10532
rect 11296 10492 11744 10520
rect 11296 10480 11302 10492
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 3418 10452 3424 10464
rect 2188 10424 3424 10452
rect 2188 10412 2194 10424
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 4522 10452 4528 10464
rect 4479 10424 4528 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 4522 10412 4528 10424
rect 4580 10412 4586 10464
rect 5074 10452 5080 10464
rect 5035 10424 5080 10452
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 5718 10452 5724 10464
rect 5679 10424 5724 10452
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7561 10455 7619 10461
rect 7561 10452 7573 10455
rect 6972 10424 7573 10452
rect 6972 10412 6978 10424
rect 7561 10421 7573 10424
rect 7607 10421 7619 10455
rect 7561 10415 7619 10421
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 8389 10455 8447 10461
rect 8389 10452 8401 10455
rect 8352 10424 8401 10452
rect 8352 10412 8358 10424
rect 8389 10421 8401 10424
rect 8435 10421 8447 10455
rect 8389 10415 8447 10421
rect 10597 10455 10655 10461
rect 10597 10421 10609 10455
rect 10643 10452 10655 10455
rect 10778 10452 10784 10464
rect 10643 10424 10784 10452
rect 10643 10421 10655 10424
rect 10597 10415 10655 10421
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 11149 10455 11207 10461
rect 11149 10421 11161 10455
rect 11195 10452 11207 10455
rect 11422 10452 11428 10464
rect 11195 10424 11428 10452
rect 11195 10421 11207 10424
rect 11149 10415 11207 10421
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 11716 10461 11744 10492
rect 13538 10480 13544 10532
rect 13596 10520 13602 10532
rect 14921 10523 14979 10529
rect 14921 10520 14933 10523
rect 13596 10492 14933 10520
rect 13596 10480 13602 10492
rect 14921 10489 14933 10492
rect 14967 10520 14979 10523
rect 15381 10523 15439 10529
rect 15381 10520 15393 10523
rect 14967 10492 15393 10520
rect 14967 10489 14979 10492
rect 14921 10483 14979 10489
rect 15381 10489 15393 10492
rect 15427 10520 15439 10523
rect 15654 10520 15660 10532
rect 15427 10492 15660 10520
rect 15427 10489 15439 10492
rect 15381 10483 15439 10489
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 16850 10520 16856 10532
rect 16811 10492 16856 10520
rect 16850 10480 16856 10492
rect 16908 10480 16914 10532
rect 11701 10455 11759 10461
rect 11701 10421 11713 10455
rect 11747 10452 11759 10455
rect 12253 10455 12311 10461
rect 12253 10452 12265 10455
rect 11747 10424 12265 10452
rect 11747 10421 11759 10424
rect 11701 10415 11759 10421
rect 12253 10421 12265 10424
rect 12299 10452 12311 10455
rect 12437 10455 12495 10461
rect 12437 10452 12449 10455
rect 12299 10424 12449 10452
rect 12299 10421 12311 10424
rect 12253 10415 12311 10421
rect 12437 10421 12449 10424
rect 12483 10452 12495 10455
rect 13630 10452 13636 10464
rect 12483 10424 13636 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 15562 10452 15568 10464
rect 15523 10424 15568 10452
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 16117 10455 16175 10461
rect 16117 10421 16129 10455
rect 16163 10452 16175 10455
rect 16482 10452 16488 10464
rect 16163 10424 16488 10452
rect 16163 10421 16175 10424
rect 16117 10415 16175 10421
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1673 10251 1731 10257
rect 1673 10217 1685 10251
rect 1719 10248 1731 10251
rect 2222 10248 2228 10260
rect 1719 10220 2228 10248
rect 1719 10217 1731 10220
rect 1673 10211 1731 10217
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 2406 10208 2412 10260
rect 2464 10248 2470 10260
rect 2682 10248 2688 10260
rect 2464 10220 2688 10248
rect 2464 10208 2470 10220
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 3421 10251 3479 10257
rect 3421 10248 3433 10251
rect 3384 10220 3433 10248
rect 3384 10208 3390 10220
rect 3421 10217 3433 10220
rect 3467 10217 3479 10251
rect 3421 10211 3479 10217
rect 3510 10208 3516 10260
rect 3568 10248 3574 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3568 10220 3801 10248
rect 3568 10208 3574 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 4614 10248 4620 10260
rect 4575 10220 4620 10248
rect 3789 10211 3847 10217
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 4798 10208 4804 10260
rect 4856 10248 4862 10260
rect 4985 10251 5043 10257
rect 4985 10248 4997 10251
rect 4856 10220 4997 10248
rect 4856 10208 4862 10220
rect 4985 10217 4997 10220
rect 5031 10217 5043 10251
rect 4985 10211 5043 10217
rect 7466 10208 7472 10260
rect 7524 10248 7530 10260
rect 7561 10251 7619 10257
rect 7561 10248 7573 10251
rect 7524 10220 7573 10248
rect 7524 10208 7530 10220
rect 7561 10217 7573 10220
rect 7607 10248 7619 10251
rect 7650 10248 7656 10260
rect 7607 10220 7656 10248
rect 7607 10217 7619 10220
rect 7561 10211 7619 10217
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 9030 10248 9036 10260
rect 8991 10220 9036 10248
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 9582 10248 9588 10260
rect 9539 10220 9588 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 9582 10208 9588 10220
rect 9640 10208 9646 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 9732 10220 9873 10248
rect 9732 10208 9738 10220
rect 9861 10217 9873 10220
rect 9907 10217 9919 10251
rect 9861 10211 9919 10217
rect 11054 10208 11060 10260
rect 11112 10248 11118 10260
rect 11517 10251 11575 10257
rect 11517 10248 11529 10251
rect 11112 10220 11529 10248
rect 11112 10208 11118 10220
rect 11517 10217 11529 10220
rect 11563 10217 11575 10251
rect 11517 10211 11575 10217
rect 12611 10251 12669 10257
rect 12611 10217 12623 10251
rect 12657 10248 12669 10251
rect 13722 10248 13728 10260
rect 12657 10220 13728 10248
rect 12657 10217 12669 10220
rect 12611 10211 12669 10217
rect 13722 10208 13728 10220
rect 13780 10248 13786 10260
rect 14645 10251 14703 10257
rect 14645 10248 14657 10251
rect 13780 10220 14657 10248
rect 13780 10208 13786 10220
rect 14645 10217 14657 10220
rect 14691 10217 14703 10251
rect 14645 10211 14703 10217
rect 2958 10180 2964 10192
rect 2919 10152 2964 10180
rect 2958 10140 2964 10152
rect 3016 10140 3022 10192
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 5721 10183 5779 10189
rect 5721 10180 5733 10183
rect 5592 10152 5733 10180
rect 5592 10140 5598 10152
rect 5721 10149 5733 10152
rect 5767 10149 5779 10183
rect 5721 10143 5779 10149
rect 8573 10183 8631 10189
rect 8573 10149 8585 10183
rect 8619 10180 8631 10183
rect 8849 10183 8907 10189
rect 8849 10180 8861 10183
rect 8619 10152 8861 10180
rect 8619 10149 8631 10152
rect 8573 10143 8631 10149
rect 8849 10149 8861 10152
rect 8895 10149 8907 10183
rect 10686 10180 10692 10192
rect 8849 10143 8907 10149
rect 9784 10152 10692 10180
rect 2682 10072 2688 10124
rect 2740 10112 2746 10124
rect 4065 10115 4123 10121
rect 2740 10084 3096 10112
rect 2740 10072 2746 10084
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3068 10053 3096 10084
rect 4065 10081 4077 10115
rect 4111 10112 4123 10115
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 4111 10084 6561 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 6549 10081 6561 10084
rect 6595 10081 6607 10115
rect 6549 10075 6607 10081
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 4522 10044 4528 10056
rect 3099 10016 4528 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10044 5871 10047
rect 6086 10044 6092 10056
rect 5859 10016 6092 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 2501 9979 2559 9985
rect 2501 9945 2513 9979
rect 2547 9976 2559 9979
rect 5626 9976 5632 9988
rect 2547 9948 5632 9976
rect 2547 9945 2559 9948
rect 2501 9939 2559 9945
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 5736 9976 5764 10007
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 6564 10044 6592 10075
rect 6638 10072 6644 10124
rect 6696 10112 6702 10124
rect 6733 10115 6791 10121
rect 6733 10112 6745 10115
rect 6696 10084 6745 10112
rect 6696 10072 6702 10084
rect 6733 10081 6745 10084
rect 6779 10081 6791 10115
rect 9784 10112 9812 10152
rect 10686 10140 10692 10152
rect 10744 10140 10750 10192
rect 12434 10140 12440 10192
rect 12492 10180 12498 10192
rect 13081 10183 13139 10189
rect 13081 10180 13093 10183
rect 12492 10152 13093 10180
rect 12492 10140 12498 10152
rect 13081 10149 13093 10152
rect 13127 10149 13139 10183
rect 13081 10143 13139 10149
rect 13170 10140 13176 10192
rect 13228 10180 13234 10192
rect 13228 10152 13273 10180
rect 13228 10140 13234 10152
rect 15470 10140 15476 10192
rect 15528 10180 15534 10192
rect 15657 10183 15715 10189
rect 15657 10180 15669 10183
rect 15528 10152 15669 10180
rect 15528 10140 15534 10152
rect 15657 10149 15669 10152
rect 15703 10149 15715 10183
rect 15657 10143 15715 10149
rect 15841 10183 15899 10189
rect 15841 10149 15853 10183
rect 15887 10180 15899 10183
rect 16114 10180 16120 10192
rect 15887 10152 16120 10180
rect 15887 10149 15899 10152
rect 15841 10143 15899 10149
rect 16114 10140 16120 10152
rect 16172 10140 16178 10192
rect 10502 10112 10508 10124
rect 6733 10075 6791 10081
rect 8128 10084 9812 10112
rect 10463 10084 10508 10112
rect 6917 10047 6975 10053
rect 6917 10044 6929 10047
rect 6564 10016 6929 10044
rect 6917 10013 6929 10016
rect 6963 10013 6975 10047
rect 6917 10007 6975 10013
rect 6273 9979 6331 9985
rect 6273 9976 6285 9979
rect 5736 9948 6285 9976
rect 6273 9945 6285 9948
rect 6319 9976 6331 9979
rect 6822 9976 6828 9988
rect 6319 9948 6828 9976
rect 6319 9945 6331 9948
rect 6273 9939 6331 9945
rect 6822 9936 6828 9948
rect 6880 9936 6886 9988
rect 8128 9985 8156 10084
rect 10502 10072 10508 10084
rect 10560 10112 10566 10124
rect 11149 10115 11207 10121
rect 11149 10112 11161 10115
rect 10560 10084 11161 10112
rect 10560 10072 10566 10084
rect 11149 10081 11161 10084
rect 11195 10081 11207 10115
rect 11149 10075 11207 10081
rect 12710 10072 12716 10124
rect 12768 10112 12774 10124
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 12768 10084 12909 10112
rect 12768 10072 12774 10084
rect 12897 10081 12909 10084
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 14093 10115 14151 10121
rect 14093 10081 14105 10115
rect 14139 10112 14151 10115
rect 14274 10112 14280 10124
rect 14139 10084 14280 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 14274 10072 14280 10084
rect 14332 10112 14338 10124
rect 14642 10112 14648 10124
rect 14332 10084 14648 10112
rect 14332 10072 14338 10084
rect 14642 10072 14648 10084
rect 14700 10072 14706 10124
rect 8570 10044 8576 10056
rect 8531 10016 8576 10044
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 8665 10047 8723 10053
rect 8665 10013 8677 10047
rect 8711 10044 8723 10047
rect 8754 10044 8760 10056
rect 8711 10016 8760 10044
rect 8711 10013 8723 10016
rect 8665 10007 8723 10013
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 8849 10047 8907 10053
rect 8849 10013 8861 10047
rect 8895 10044 8907 10047
rect 9030 10044 9036 10056
rect 8895 10016 9036 10044
rect 8895 10013 8907 10016
rect 8849 10007 8907 10013
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 10778 10044 10784 10056
rect 10691 10016 10784 10044
rect 10778 10004 10784 10016
rect 10836 10044 10842 10056
rect 12437 10047 12495 10053
rect 12437 10044 12449 10047
rect 10836 10016 12449 10044
rect 10836 10004 10842 10016
rect 12437 10013 12449 10016
rect 12483 10044 12495 10047
rect 12618 10044 12624 10056
rect 12483 10016 12624 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 15930 10044 15936 10056
rect 15891 10016 15936 10044
rect 15930 10004 15936 10016
rect 15988 10004 15994 10056
rect 8113 9979 8171 9985
rect 8113 9945 8125 9979
rect 8159 9945 8171 9979
rect 8113 9939 8171 9945
rect 14182 9936 14188 9988
rect 14240 9976 14246 9988
rect 15378 9976 15384 9988
rect 14240 9948 15148 9976
rect 15339 9948 15384 9976
rect 14240 9936 14246 9948
rect 3878 9868 3884 9920
rect 3936 9908 3942 9920
rect 4249 9911 4307 9917
rect 4249 9908 4261 9911
rect 3936 9880 4261 9908
rect 3936 9868 3942 9880
rect 4249 9877 4261 9880
rect 4295 9877 4307 9911
rect 5258 9908 5264 9920
rect 5219 9880 5264 9908
rect 4249 9871 4307 9877
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 7929 9911 7987 9917
rect 7929 9877 7941 9911
rect 7975 9908 7987 9911
rect 8754 9908 8760 9920
rect 7975 9880 8760 9908
rect 7975 9877 7987 9880
rect 7929 9871 7987 9877
rect 8754 9868 8760 9880
rect 8812 9868 8818 9920
rect 10229 9911 10287 9917
rect 10229 9877 10241 9911
rect 10275 9908 10287 9911
rect 11054 9908 11060 9920
rect 10275 9880 11060 9908
rect 10275 9877 10287 9880
rect 10229 9871 10287 9877
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11882 9908 11888 9920
rect 11843 9880 11888 9908
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 13906 9908 13912 9920
rect 13867 9880 13912 9908
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 14274 9908 14280 9920
rect 14235 9880 14280 9908
rect 14274 9868 14280 9880
rect 14332 9868 14338 9920
rect 15120 9917 15148 9948
rect 15378 9936 15384 9948
rect 15436 9936 15442 9988
rect 15105 9911 15163 9917
rect 15105 9877 15117 9911
rect 15151 9908 15163 9911
rect 15562 9908 15568 9920
rect 15151 9880 15568 9908
rect 15151 9877 15163 9880
rect 15105 9871 15163 9877
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3605 9707 3663 9713
rect 3605 9704 3617 9707
rect 3016 9676 3617 9704
rect 3016 9664 3022 9676
rect 3605 9673 3617 9676
rect 3651 9673 3663 9707
rect 9030 9704 9036 9716
rect 8991 9676 9036 9704
rect 3605 9667 3663 9673
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 9677 9707 9735 9713
rect 9677 9673 9689 9707
rect 9723 9704 9735 9707
rect 10502 9704 10508 9716
rect 9723 9676 10508 9704
rect 9723 9673 9735 9676
rect 9677 9667 9735 9673
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 10689 9707 10747 9713
rect 10689 9673 10701 9707
rect 10735 9704 10747 9707
rect 10778 9704 10784 9716
rect 10735 9676 10784 9704
rect 10735 9673 10747 9676
rect 10689 9667 10747 9673
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 13170 9704 13176 9716
rect 12544 9676 13176 9704
rect 2501 9639 2559 9645
rect 2501 9605 2513 9639
rect 2547 9636 2559 9639
rect 2682 9636 2688 9648
rect 2547 9608 2688 9636
rect 2547 9605 2559 9608
rect 2501 9599 2559 9605
rect 2682 9596 2688 9608
rect 2740 9596 2746 9648
rect 6270 9596 6276 9648
rect 6328 9636 6334 9648
rect 6457 9639 6515 9645
rect 6457 9636 6469 9639
rect 6328 9608 6469 9636
rect 6328 9596 6334 9608
rect 6457 9605 6469 9608
rect 6503 9636 6515 9639
rect 6549 9639 6607 9645
rect 6549 9636 6561 9639
rect 6503 9608 6561 9636
rect 6503 9605 6515 9608
rect 6457 9599 6515 9605
rect 6549 9605 6561 9608
rect 6595 9605 6607 9639
rect 6549 9599 6607 9605
rect 6822 9596 6828 9648
rect 6880 9636 6886 9648
rect 6917 9639 6975 9645
rect 6917 9636 6929 9639
rect 6880 9608 6929 9636
rect 6880 9596 6886 9608
rect 6917 9605 6929 9608
rect 6963 9605 6975 9639
rect 6917 9599 6975 9605
rect 11054 9596 11060 9648
rect 11112 9636 11118 9648
rect 11790 9636 11796 9648
rect 11112 9608 11796 9636
rect 11112 9596 11118 9608
rect 11790 9596 11796 9608
rect 11848 9596 11854 9648
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 2648 9540 3065 9568
rect 2648 9528 2654 9540
rect 3053 9537 3065 9540
rect 3099 9537 3111 9571
rect 3053 9531 3111 9537
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9568 8171 9571
rect 8754 9568 8760 9580
rect 8159 9540 8760 9568
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 8754 9528 8760 9540
rect 8812 9568 8818 9580
rect 9401 9571 9459 9577
rect 9401 9568 9413 9571
rect 8812 9540 9413 9568
rect 8812 9528 8818 9540
rect 9401 9537 9413 9540
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 1578 9500 1584 9512
rect 1539 9472 1584 9500
rect 1578 9460 1584 9472
rect 1636 9460 1642 9512
rect 2869 9503 2927 9509
rect 2869 9469 2881 9503
rect 2915 9469 2927 9503
rect 2869 9463 2927 9469
rect 1854 9432 1860 9444
rect 1815 9404 1860 9432
rect 1854 9392 1860 9404
rect 1912 9392 1918 9444
rect 2884 9432 2912 9463
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4522 9509 4528 9512
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 4212 9472 4261 9500
rect 4212 9460 4218 9472
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4516 9500 4528 9509
rect 4483 9472 4528 9500
rect 4249 9463 4307 9469
rect 4516 9463 4528 9472
rect 4522 9460 4528 9463
rect 4580 9460 4586 9512
rect 6273 9503 6331 9509
rect 6273 9469 6285 9503
rect 6319 9500 6331 9503
rect 8386 9500 8392 9512
rect 6319 9472 7512 9500
rect 8347 9472 8392 9500
rect 6319 9469 6331 9472
rect 6273 9463 6331 9469
rect 3694 9432 3700 9444
rect 2884 9404 3700 9432
rect 3694 9392 3700 9404
rect 3752 9432 3758 9444
rect 4338 9432 4344 9444
rect 3752 9404 4344 9432
rect 3752 9392 3758 9404
rect 4338 9392 4344 9404
rect 4396 9392 4402 9444
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 3234 9364 3240 9376
rect 2832 9336 3240 9364
rect 2832 9324 2838 9336
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 4154 9364 4160 9376
rect 4067 9336 4160 9364
rect 4154 9324 4160 9336
rect 4212 9364 4218 9376
rect 4890 9364 4896 9376
rect 4212 9336 4896 9364
rect 4212 9324 4218 9336
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5629 9367 5687 9373
rect 5629 9333 5641 9367
rect 5675 9364 5687 9367
rect 6288 9364 6316 9463
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 7484 9441 7512 9472
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 9416 9500 9444 9531
rect 9490 9528 9496 9580
rect 9548 9568 9554 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 9548 9540 10149 9568
rect 9548 9528 9554 9540
rect 10137 9537 10149 9540
rect 10183 9568 10195 9571
rect 11146 9568 11152 9580
rect 10183 9540 11152 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 11146 9528 11152 9540
rect 11204 9528 11210 9580
rect 10229 9503 10287 9509
rect 10229 9500 10241 9503
rect 9416 9472 10241 9500
rect 10229 9469 10241 9472
rect 10275 9469 10287 9503
rect 10229 9463 10287 9469
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 12544 9500 12572 9676
rect 13170 9664 13176 9676
rect 13228 9664 13234 9716
rect 15470 9664 15476 9716
rect 15528 9704 15534 9716
rect 15749 9707 15807 9713
rect 15749 9704 15761 9707
rect 15528 9676 15761 9704
rect 15528 9664 15534 9676
rect 15749 9673 15761 9676
rect 15795 9673 15807 9707
rect 16850 9704 16856 9716
rect 16811 9676 16856 9704
rect 15749 9667 15807 9673
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 12894 9636 12900 9648
rect 12855 9608 12900 9636
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 13354 9636 13360 9648
rect 13315 9608 13360 9636
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 12299 9472 12572 9500
rect 12713 9503 12771 9509
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 12713 9469 12725 9503
rect 12759 9500 12771 9503
rect 13372 9500 13400 9596
rect 18046 9568 18052 9580
rect 15304 9540 18052 9568
rect 12759 9472 13400 9500
rect 12759 9469 12771 9472
rect 12713 9463 12771 9469
rect 13630 9460 13636 9512
rect 13688 9500 13694 9512
rect 13817 9503 13875 9509
rect 13817 9500 13829 9503
rect 13688 9472 13829 9500
rect 13688 9460 13694 9472
rect 13817 9469 13829 9472
rect 13863 9469 13875 9503
rect 13817 9463 13875 9469
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 14073 9503 14131 9509
rect 14073 9500 14085 9503
rect 13964 9472 14085 9500
rect 13964 9460 13970 9472
rect 14073 9469 14085 9472
rect 14119 9469 14131 9503
rect 14073 9463 14131 9469
rect 14366 9460 14372 9512
rect 14424 9500 14430 9512
rect 14458 9500 14464 9512
rect 14424 9472 14464 9500
rect 14424 9460 14430 9472
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 7193 9435 7251 9441
rect 7193 9432 7205 9435
rect 6972 9404 7205 9432
rect 6972 9392 6978 9404
rect 7193 9401 7205 9404
rect 7239 9401 7251 9435
rect 7193 9395 7251 9401
rect 7469 9435 7527 9441
rect 7469 9401 7481 9435
rect 7515 9432 7527 9435
rect 7558 9432 7564 9444
rect 7515 9404 7564 9432
rect 7515 9401 7527 9404
rect 7469 9395 7527 9401
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 10870 9392 10876 9444
rect 10928 9432 10934 9444
rect 15304 9432 15332 9540
rect 18046 9528 18052 9540
rect 18104 9528 18110 9580
rect 16301 9503 16359 9509
rect 16301 9469 16313 9503
rect 16347 9500 16359 9503
rect 16850 9500 16856 9512
rect 16347 9472 16856 9500
rect 16347 9469 16359 9472
rect 16301 9463 16359 9469
rect 16850 9460 16856 9472
rect 16908 9460 16914 9512
rect 16114 9432 16120 9444
rect 10928 9404 15332 9432
rect 16075 9404 16120 9432
rect 10928 9392 10934 9404
rect 16114 9392 16120 9404
rect 16172 9392 16178 9444
rect 5675 9336 6316 9364
rect 6457 9367 6515 9373
rect 5675 9333 5687 9336
rect 5629 9327 5687 9333
rect 6457 9333 6469 9367
rect 6503 9364 6515 9367
rect 7377 9367 7435 9373
rect 7377 9364 7389 9367
rect 6503 9336 7389 9364
rect 6503 9333 6515 9336
rect 6457 9327 6515 9333
rect 7377 9333 7389 9336
rect 7423 9333 7435 9367
rect 7377 9327 7435 9333
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 8573 9367 8631 9373
rect 8573 9364 8585 9367
rect 8444 9336 8585 9364
rect 8444 9324 8450 9336
rect 8573 9333 8585 9336
rect 8619 9333 8631 9367
rect 10134 9364 10140 9376
rect 10095 9336 10140 9364
rect 8573 9327 8631 9333
rect 10134 9324 10140 9336
rect 10192 9364 10198 9376
rect 10965 9367 11023 9373
rect 10965 9364 10977 9367
rect 10192 9336 10977 9364
rect 10192 9324 10198 9336
rect 10965 9333 10977 9336
rect 11011 9333 11023 9367
rect 11146 9364 11152 9376
rect 11107 9336 11152 9364
rect 10965 9327 11023 9333
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 13630 9364 13636 9376
rect 11296 9336 13636 9364
rect 11296 9324 11302 9336
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 15194 9364 15200 9376
rect 15155 9336 15200 9364
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 16485 9367 16543 9373
rect 16485 9333 16497 9367
rect 16531 9364 16543 9367
rect 17494 9364 17500 9376
rect 16531 9336 17500 9364
rect 16531 9333 16543 9336
rect 16485 9327 16543 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1673 9163 1731 9169
rect 1673 9129 1685 9163
rect 1719 9160 1731 9163
rect 2038 9160 2044 9172
rect 1719 9132 2044 9160
rect 1719 9129 1731 9132
rect 1673 9123 1731 9129
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 3789 9163 3847 9169
rect 3789 9160 3801 9163
rect 2924 9132 3801 9160
rect 2924 9120 2930 9132
rect 3789 9129 3801 9132
rect 3835 9129 3847 9163
rect 3789 9123 3847 9129
rect 4341 9163 4399 9169
rect 4341 9129 4353 9163
rect 4387 9160 4399 9163
rect 4522 9160 4528 9172
rect 4387 9132 4528 9160
rect 4387 9129 4399 9132
rect 4341 9123 4399 9129
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 8294 9120 8300 9172
rect 8352 9120 8358 9172
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 8628 9132 8953 9160
rect 8628 9120 8634 9132
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 9490 9160 9496 9172
rect 9451 9132 9496 9160
rect 8941 9123 8999 9129
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 9858 9160 9864 9172
rect 9819 9132 9864 9160
rect 9858 9120 9864 9132
rect 9916 9120 9922 9172
rect 10686 9160 10692 9172
rect 10647 9132 10692 9160
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 12492 9132 12537 9160
rect 12492 9120 12498 9132
rect 12710 9120 12716 9172
rect 12768 9160 12774 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12768 9132 13001 9160
rect 12768 9120 12774 9132
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 14642 9160 14648 9172
rect 14603 9132 14648 9160
rect 12989 9123 13047 9129
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 15930 9160 15936 9172
rect 15891 9132 15936 9160
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 2774 9052 2780 9104
rect 2832 9092 2838 9104
rect 2961 9095 3019 9101
rect 2961 9092 2973 9095
rect 2832 9064 2973 9092
rect 2832 9052 2838 9064
rect 2961 9061 2973 9064
rect 3007 9092 3019 9095
rect 3970 9092 3976 9104
rect 3007 9064 3976 9092
rect 3007 9061 3019 9064
rect 2961 9055 3019 9061
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 5169 9095 5227 9101
rect 5169 9092 5181 9095
rect 4212 9064 5181 9092
rect 4212 9052 4218 9064
rect 5169 9061 5181 9064
rect 5215 9092 5227 9095
rect 5258 9092 5264 9104
rect 5215 9064 5264 9092
rect 5215 9061 5227 9064
rect 5169 9055 5227 9061
rect 5258 9052 5264 9064
rect 5316 9052 5322 9104
rect 6362 9052 6368 9104
rect 6420 9092 6426 9104
rect 6730 9092 6736 9104
rect 6420 9064 6736 9092
rect 6420 9052 6426 9064
rect 6730 9052 6736 9064
rect 6788 9052 6794 9104
rect 8312 9092 8340 9120
rect 7024 9064 8340 9092
rect 2317 9027 2375 9033
rect 2317 8993 2329 9027
rect 2363 9024 2375 9027
rect 3050 9024 3056 9036
rect 2363 8996 3056 9024
rect 2363 8993 2375 8996
rect 2317 8987 2375 8993
rect 3050 8984 3056 8996
rect 3108 8984 3114 9036
rect 3510 9024 3516 9036
rect 3471 8996 3516 9024
rect 3510 8984 3516 8996
rect 3568 8984 3574 9036
rect 4985 9027 5043 9033
rect 4985 8993 4997 9027
rect 5031 9024 5043 9027
rect 5031 8996 6500 9024
rect 5031 8993 5043 8996
rect 4985 8987 5043 8993
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 5258 8956 5264 8968
rect 5219 8928 5264 8956
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5500 8928 6009 8956
rect 5500 8916 5506 8928
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 5166 8848 5172 8900
rect 5224 8888 5230 8900
rect 5224 8860 5488 8888
rect 5224 8848 5230 8860
rect 2501 8823 2559 8829
rect 2501 8789 2513 8823
rect 2547 8820 2559 8823
rect 2682 8820 2688 8832
rect 2547 8792 2688 8820
rect 2547 8789 2559 8792
rect 2501 8783 2559 8789
rect 2682 8780 2688 8792
rect 2740 8780 2746 8832
rect 4709 8823 4767 8829
rect 4709 8789 4721 8823
rect 4755 8820 4767 8823
rect 5350 8820 5356 8832
rect 4755 8792 5356 8820
rect 4755 8789 4767 8792
rect 4709 8783 4767 8789
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 5460 8820 5488 8860
rect 5629 8823 5687 8829
rect 5629 8820 5641 8823
rect 5460 8792 5641 8820
rect 5629 8789 5641 8792
rect 5675 8820 5687 8823
rect 6086 8820 6092 8832
rect 5675 8792 6092 8820
rect 5675 8789 5687 8792
rect 5629 8783 5687 8789
rect 6086 8780 6092 8792
rect 6144 8780 6150 8832
rect 6472 8829 6500 8996
rect 6822 8984 6828 9036
rect 6880 9024 6886 9036
rect 7024 9033 7052 9064
rect 13538 9052 13544 9104
rect 13596 9092 13602 9104
rect 13814 9092 13820 9104
rect 13596 9064 13820 9092
rect 13596 9052 13602 9064
rect 13814 9052 13820 9064
rect 13872 9092 13878 9104
rect 14185 9095 14243 9101
rect 14185 9092 14197 9095
rect 13872 9064 14197 9092
rect 13872 9052 13878 9064
rect 14185 9061 14197 9064
rect 14231 9061 14243 9095
rect 14185 9055 14243 9061
rect 7009 9027 7067 9033
rect 7009 9024 7021 9027
rect 6880 8996 7021 9024
rect 6880 8984 6886 8996
rect 7009 8993 7021 8996
rect 7055 8993 7067 9027
rect 7009 8987 7067 8993
rect 7276 9027 7334 9033
rect 7276 8993 7288 9027
rect 7322 9024 7334 9027
rect 7558 9024 7564 9036
rect 7322 8996 7564 9024
rect 7322 8993 7334 8996
rect 7276 8987 7334 8993
rect 7558 8984 7564 8996
rect 7616 9024 7622 9036
rect 8938 9024 8944 9036
rect 7616 8996 8944 9024
rect 7616 8984 7622 8996
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 9674 8984 9680 8996
rect 9732 9024 9738 9036
rect 10042 9024 10048 9036
rect 9732 8996 10048 9024
rect 9732 8984 9738 8996
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 11330 9033 11336 9036
rect 11324 8987 11336 9033
rect 11388 9024 11394 9036
rect 11388 8996 11424 9024
rect 11330 8984 11336 8987
rect 11388 8984 11394 8996
rect 12342 8984 12348 9036
rect 12400 9024 12406 9036
rect 15013 9027 15071 9033
rect 15013 9024 15025 9027
rect 12400 8996 15025 9024
rect 12400 8984 12406 8996
rect 15013 8993 15025 8996
rect 15059 8993 15071 9027
rect 15013 8987 15071 8993
rect 15289 9027 15347 9033
rect 15289 8993 15301 9027
rect 15335 9024 15347 9027
rect 15378 9024 15384 9036
rect 15335 8996 15384 9024
rect 15335 8993 15347 8996
rect 15289 8987 15347 8993
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 16390 9024 16396 9036
rect 16351 8996 16396 9024
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 11054 8956 11060 8968
rect 11015 8928 11060 8956
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 14182 8956 14188 8968
rect 14143 8928 14188 8956
rect 14182 8916 14188 8928
rect 14240 8916 14246 8968
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8956 14335 8959
rect 14642 8956 14648 8968
rect 14323 8928 14648 8956
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 13541 8891 13599 8897
rect 13541 8857 13553 8891
rect 13587 8888 13599 8891
rect 14292 8888 14320 8919
rect 14642 8916 14648 8928
rect 14700 8916 14706 8968
rect 13587 8860 14320 8888
rect 13587 8857 13599 8860
rect 13541 8851 13599 8857
rect 6457 8823 6515 8829
rect 6457 8789 6469 8823
rect 6503 8820 6515 8823
rect 6730 8820 6736 8832
rect 6503 8792 6736 8820
rect 6503 8789 6515 8792
rect 6457 8783 6515 8789
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 6914 8820 6920 8832
rect 6875 8792 6920 8820
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 8168 8792 8401 8820
rect 8168 8780 8174 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 8389 8783 8447 8789
rect 10321 8823 10379 8829
rect 10321 8789 10333 8823
rect 10367 8820 10379 8823
rect 10502 8820 10508 8832
rect 10367 8792 10508 8820
rect 10367 8789 10379 8792
rect 10321 8783 10379 8789
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 13630 8780 13636 8832
rect 13688 8820 13694 8832
rect 13725 8823 13783 8829
rect 13725 8820 13737 8823
rect 13688 8792 13737 8820
rect 13688 8780 13694 8792
rect 13725 8789 13737 8792
rect 13771 8789 13783 8823
rect 13725 8783 13783 8789
rect 15286 8780 15292 8832
rect 15344 8820 15350 8832
rect 15473 8823 15531 8829
rect 15473 8820 15485 8823
rect 15344 8792 15485 8820
rect 15344 8780 15350 8792
rect 15473 8789 15485 8792
rect 15519 8789 15531 8823
rect 15473 8783 15531 8789
rect 16298 8780 16304 8832
rect 16356 8820 16362 8832
rect 16577 8823 16635 8829
rect 16577 8820 16589 8823
rect 16356 8792 16589 8820
rect 16356 8780 16362 8792
rect 16577 8789 16589 8792
rect 16623 8789 16635 8823
rect 16577 8783 16635 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2501 8619 2559 8625
rect 2501 8585 2513 8619
rect 2547 8616 2559 8619
rect 2547 8588 2820 8616
rect 2547 8585 2559 8588
rect 2501 8579 2559 8585
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 1854 8480 1860 8492
rect 1719 8452 1860 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 2792 8424 2820 8588
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3694 8616 3700 8628
rect 2924 8588 3700 8616
rect 2924 8576 2930 8588
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 3970 8576 3976 8628
rect 4028 8616 4034 8628
rect 6638 8616 6644 8628
rect 4028 8588 5764 8616
rect 6551 8588 6644 8616
rect 4028 8576 4034 8588
rect 3510 8548 3516 8560
rect 3471 8520 3516 8548
rect 3510 8508 3516 8520
rect 3568 8508 3574 8560
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 5629 8551 5687 8557
rect 5629 8548 5641 8551
rect 5592 8520 5641 8548
rect 5592 8508 5598 8520
rect 5629 8517 5641 8520
rect 5675 8517 5687 8551
rect 5736 8548 5764 8588
rect 6638 8576 6644 8588
rect 6696 8616 6702 8628
rect 7558 8616 7564 8628
rect 6696 8588 7564 8616
rect 6696 8576 6702 8588
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 8202 8616 8208 8628
rect 7883 8588 8208 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 8202 8576 8208 8588
rect 8260 8616 8266 8628
rect 8570 8616 8576 8628
rect 8260 8588 8576 8616
rect 8260 8576 8266 8588
rect 8570 8576 8576 8588
rect 8628 8616 8634 8628
rect 10870 8616 10876 8628
rect 8628 8588 10876 8616
rect 8628 8576 8634 8588
rect 10870 8576 10876 8588
rect 10928 8616 10934 8628
rect 11054 8616 11060 8628
rect 10928 8588 11060 8616
rect 10928 8576 10934 8588
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11330 8576 11336 8628
rect 11388 8616 11394 8628
rect 11425 8619 11483 8625
rect 11425 8616 11437 8619
rect 11388 8588 11437 8616
rect 11388 8576 11394 8588
rect 11425 8585 11437 8588
rect 11471 8616 11483 8619
rect 11698 8616 11704 8628
rect 11471 8588 11704 8616
rect 11471 8585 11483 8588
rect 11425 8579 11483 8585
rect 11698 8576 11704 8588
rect 11756 8616 11762 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 11756 8588 11805 8616
rect 11756 8576 11762 8588
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 11793 8579 11851 8585
rect 7929 8551 7987 8557
rect 7929 8548 7941 8551
rect 5736 8520 7941 8548
rect 5629 8511 5687 8517
rect 7929 8517 7941 8520
rect 7975 8517 7987 8551
rect 7929 8511 7987 8517
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 8389 8551 8447 8557
rect 8389 8548 8401 8551
rect 8352 8520 8401 8548
rect 8352 8508 8358 8520
rect 8389 8517 8401 8520
rect 8435 8517 8447 8551
rect 8389 8511 8447 8517
rect 9674 8508 9680 8560
rect 9732 8548 9738 8560
rect 9953 8551 10011 8557
rect 9953 8548 9965 8551
rect 9732 8520 9965 8548
rect 9732 8508 9738 8520
rect 9953 8517 9965 8520
rect 9999 8517 10011 8551
rect 9953 8511 10011 8517
rect 3050 8440 3056 8492
rect 3108 8480 3114 8492
rect 3329 8483 3387 8489
rect 3329 8480 3341 8483
rect 3108 8452 3341 8480
rect 3108 8440 3114 8452
rect 3329 8449 3341 8452
rect 3375 8449 3387 8483
rect 3329 8443 3387 8449
rect 6086 8440 6092 8492
rect 6144 8480 6150 8492
rect 7098 8480 7104 8492
rect 6144 8452 7104 8480
rect 6144 8440 6150 8452
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7282 8480 7288 8492
rect 7243 8452 7288 8480
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 8846 8480 8852 8492
rect 8536 8452 8852 8480
rect 8536 8440 8542 8452
rect 8846 8440 8852 8452
rect 8904 8440 8910 8492
rect 9306 8480 9312 8492
rect 9267 8452 9312 8480
rect 9306 8440 9312 8452
rect 9364 8480 9370 8492
rect 10318 8480 10324 8492
rect 9364 8452 10324 8480
rect 9364 8440 9370 8452
rect 10318 8440 10324 8452
rect 10376 8440 10382 8492
rect 10502 8480 10508 8492
rect 10463 8452 10508 8480
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 11808 8480 11836 8579
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 13964 8588 15240 8616
rect 13964 8576 13970 8588
rect 12434 8508 12440 8560
rect 12492 8548 12498 8560
rect 12529 8551 12587 8557
rect 12529 8548 12541 8551
rect 12492 8520 12541 8548
rect 12492 8508 12498 8520
rect 12529 8517 12541 8520
rect 12575 8517 12587 8551
rect 12529 8511 12587 8517
rect 13722 8508 13728 8560
rect 13780 8548 13786 8560
rect 14093 8551 14151 8557
rect 14093 8548 14105 8551
rect 13780 8520 14105 8548
rect 13780 8508 13786 8520
rect 14093 8517 14105 8520
rect 14139 8548 14151 8551
rect 15212 8548 15240 8588
rect 15378 8576 15384 8628
rect 15436 8616 15442 8628
rect 16209 8619 16267 8625
rect 16209 8616 16221 8619
rect 15436 8588 16221 8616
rect 15436 8576 15442 8588
rect 16209 8585 16221 8588
rect 16255 8585 16267 8619
rect 16209 8579 16267 8585
rect 16390 8576 16396 8628
rect 16448 8616 16454 8628
rect 16577 8619 16635 8625
rect 16577 8616 16589 8619
rect 16448 8588 16589 8616
rect 16448 8576 16454 8588
rect 16577 8585 16589 8588
rect 16623 8585 16635 8619
rect 16577 8579 16635 8585
rect 15657 8551 15715 8557
rect 15657 8548 15669 8551
rect 14139 8520 14320 8548
rect 15212 8520 15669 8548
rect 14139 8517 14151 8520
rect 14093 8511 14151 8517
rect 13078 8480 13084 8492
rect 11808 8452 13084 8480
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 14292 8489 14320 8520
rect 15657 8517 15669 8520
rect 15703 8517 15715 8551
rect 15657 8511 15715 8517
rect 14277 8483 14335 8489
rect 14277 8449 14289 8483
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8412 1458 8424
rect 1946 8412 1952 8424
rect 1452 8384 1952 8412
rect 1452 8372 1458 8384
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2774 8372 2780 8424
rect 2832 8372 2838 8424
rect 3142 8412 3148 8424
rect 2976 8384 3148 8412
rect 2976 8344 3004 8384
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 3234 8372 3240 8424
rect 3292 8412 3298 8424
rect 3694 8412 3700 8424
rect 3292 8384 3700 8412
rect 3292 8372 3298 8384
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 4157 8415 4215 8421
rect 4157 8381 4169 8415
rect 4203 8412 4215 8415
rect 4249 8415 4307 8421
rect 4249 8412 4261 8415
rect 4203 8384 4261 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 4249 8381 4261 8384
rect 4295 8412 4307 8415
rect 4890 8412 4896 8424
rect 4295 8384 4896 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 6273 8415 6331 8421
rect 6273 8381 6285 8415
rect 6319 8412 6331 8415
rect 7006 8412 7012 8424
rect 6319 8384 7012 8412
rect 6319 8381 6331 8384
rect 6273 8375 6331 8381
rect 7006 8372 7012 8384
rect 7064 8372 7070 8424
rect 8662 8412 8668 8424
rect 8623 8384 8668 8412
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 9490 8412 9496 8424
rect 8864 8384 9496 8412
rect 4522 8353 4528 8356
rect 2792 8316 3004 8344
rect 3053 8347 3111 8353
rect 2792 8285 2820 8316
rect 3053 8313 3065 8347
rect 3099 8344 3111 8347
rect 3513 8347 3571 8353
rect 3513 8344 3525 8347
rect 3099 8316 3525 8344
rect 3099 8313 3111 8316
rect 3053 8307 3111 8313
rect 3513 8313 3525 8316
rect 3559 8313 3571 8347
rect 4516 8344 4528 8353
rect 3513 8307 3571 8313
rect 3620 8316 4200 8344
rect 4483 8316 4528 8344
rect 2767 8279 2825 8285
rect 2767 8245 2779 8279
rect 2813 8245 2825 8279
rect 2767 8239 2825 8245
rect 3237 8279 3295 8285
rect 3237 8245 3249 8279
rect 3283 8276 3295 8279
rect 3418 8276 3424 8288
rect 3283 8248 3424 8276
rect 3283 8245 3295 8248
rect 3237 8239 3295 8245
rect 3418 8236 3424 8248
rect 3476 8276 3482 8288
rect 3620 8276 3648 8316
rect 3476 8248 3648 8276
rect 4172 8276 4200 8316
rect 4516 8307 4528 8316
rect 4522 8304 4528 8307
rect 4580 8304 4586 8356
rect 8864 8353 8892 8384
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 8205 8347 8263 8353
rect 8205 8344 8217 8347
rect 4632 8316 8217 8344
rect 4632 8276 4660 8316
rect 8205 8313 8217 8316
rect 8251 8344 8263 8347
rect 8849 8347 8907 8353
rect 8849 8344 8861 8347
rect 8251 8316 8861 8344
rect 8251 8313 8263 8316
rect 8205 8307 8263 8313
rect 8849 8313 8861 8316
rect 8895 8313 8907 8347
rect 8849 8307 8907 8313
rect 8938 8304 8944 8356
rect 8996 8344 9002 8356
rect 10520 8344 10548 8440
rect 12066 8372 12072 8424
rect 12124 8412 12130 8424
rect 12253 8415 12311 8421
rect 12253 8412 12265 8415
rect 12124 8384 12265 8412
rect 12124 8372 12130 8384
rect 12253 8381 12265 8384
rect 12299 8412 12311 8415
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12299 8384 12817 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12805 8381 12817 8384
rect 12851 8412 12863 8415
rect 12894 8412 12900 8424
rect 12851 8384 12900 8412
rect 12851 8381 12863 8384
rect 12805 8375 12863 8381
rect 12894 8372 12900 8384
rect 12952 8372 12958 8424
rect 14292 8412 14320 8443
rect 16114 8412 16120 8424
rect 14292 8384 16120 8412
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 8996 8316 10548 8344
rect 8996 8304 9002 8316
rect 13538 8304 13544 8356
rect 13596 8344 13602 8356
rect 13633 8347 13691 8353
rect 13633 8344 13645 8347
rect 13596 8316 13645 8344
rect 13596 8304 13602 8316
rect 13633 8313 13645 8316
rect 13679 8313 13691 8347
rect 13633 8307 13691 8313
rect 14544 8347 14602 8353
rect 14544 8313 14556 8347
rect 14590 8344 14602 8347
rect 14642 8344 14648 8356
rect 14590 8316 14648 8344
rect 14590 8313 14602 8316
rect 14544 8307 14602 8313
rect 14642 8304 14648 8316
rect 14700 8304 14706 8356
rect 16482 8304 16488 8356
rect 16540 8344 16546 8356
rect 16761 8347 16819 8353
rect 16761 8344 16773 8347
rect 16540 8316 16773 8344
rect 16540 8304 16546 8316
rect 16761 8313 16773 8316
rect 16807 8313 16819 8347
rect 16761 8307 16819 8313
rect 4172 8248 4660 8276
rect 7929 8279 7987 8285
rect 3476 8236 3482 8248
rect 7929 8245 7941 8279
rect 7975 8276 7987 8279
rect 9769 8279 9827 8285
rect 9769 8276 9781 8279
rect 7975 8248 9781 8276
rect 7975 8245 7987 8248
rect 7929 8239 7987 8245
rect 9769 8245 9781 8248
rect 9815 8276 9827 8279
rect 9858 8276 9864 8288
rect 9815 8248 9864 8276
rect 9815 8245 9827 8248
rect 9769 8239 9827 8245
rect 9858 8236 9864 8248
rect 9916 8276 9922 8288
rect 10413 8279 10471 8285
rect 10413 8276 10425 8279
rect 9916 8248 10425 8276
rect 9916 8236 9922 8248
rect 10413 8245 10425 8248
rect 10459 8276 10471 8279
rect 10962 8276 10968 8288
rect 10459 8248 10968 8276
rect 10459 8245 10471 8248
rect 10413 8239 10471 8245
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 12989 8279 13047 8285
rect 12989 8245 13001 8279
rect 13035 8276 13047 8279
rect 13446 8276 13452 8288
rect 13035 8248 13452 8276
rect 13035 8245 13047 8248
rect 12989 8239 13047 8245
rect 13446 8236 13452 8248
rect 13504 8236 13510 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2314 8072 2320 8084
rect 2227 8044 2320 8072
rect 2314 8032 2320 8044
rect 2372 8072 2378 8084
rect 3050 8072 3056 8084
rect 2372 8044 3056 8072
rect 2372 8032 2378 8044
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 3418 8072 3424 8084
rect 3379 8044 3424 8072
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 4154 8072 4160 8084
rect 3927 8044 4160 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 4341 8075 4399 8081
rect 4341 8041 4353 8075
rect 4387 8072 4399 8075
rect 4522 8072 4528 8084
rect 4387 8044 4528 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 4522 8032 4528 8044
rect 4580 8072 4586 8084
rect 4709 8075 4767 8081
rect 4709 8072 4721 8075
rect 4580 8044 4721 8072
rect 4580 8032 4586 8044
rect 4709 8041 4721 8044
rect 4755 8072 4767 8075
rect 5258 8072 5264 8084
rect 4755 8044 5264 8072
rect 4755 8041 4767 8044
rect 4709 8035 4767 8041
rect 5258 8032 5264 8044
rect 5316 8072 5322 8084
rect 6273 8075 6331 8081
rect 6273 8072 6285 8075
rect 5316 8044 6285 8072
rect 5316 8032 5322 8044
rect 6273 8041 6285 8044
rect 6319 8041 6331 8075
rect 6273 8035 6331 8041
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 8662 8072 8668 8084
rect 8619 8044 8668 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 8938 8072 8944 8084
rect 8899 8044 8944 8072
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10413 8075 10471 8081
rect 10413 8072 10425 8075
rect 10100 8044 10425 8072
rect 10100 8032 10106 8044
rect 10413 8041 10425 8044
rect 10459 8041 10471 8075
rect 10413 8035 10471 8041
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 11146 8072 11152 8084
rect 10919 8044 11152 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 11146 8032 11152 8044
rect 11204 8072 11210 8084
rect 12342 8072 12348 8084
rect 11204 8044 12348 8072
rect 11204 8032 11210 8044
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 14182 8072 14188 8084
rect 14143 8044 14188 8072
rect 14182 8032 14188 8044
rect 14240 8072 14246 8084
rect 15289 8075 15347 8081
rect 15289 8072 15301 8075
rect 14240 8044 15301 8072
rect 14240 8032 14246 8044
rect 15289 8041 15301 8044
rect 15335 8041 15347 8075
rect 15289 8035 15347 8041
rect 17681 8075 17739 8081
rect 17681 8041 17693 8075
rect 17727 8041 17739 8075
rect 17681 8035 17739 8041
rect 2961 8007 3019 8013
rect 2961 7973 2973 8007
rect 3007 8004 3019 8007
rect 3234 8004 3240 8016
rect 3007 7976 3240 8004
rect 3007 7973 3019 7976
rect 2961 7967 3019 7973
rect 3234 7964 3240 7976
rect 3292 8004 3298 8016
rect 3602 8004 3608 8016
rect 3292 7976 3608 8004
rect 3292 7964 3298 7976
rect 3602 7964 3608 7976
rect 3660 7964 3666 8016
rect 8021 8007 8079 8013
rect 8021 7973 8033 8007
rect 8067 8004 8079 8007
rect 8294 8004 8300 8016
rect 8067 7976 8300 8004
rect 8067 7973 8079 7976
rect 8021 7967 8079 7973
rect 8294 7964 8300 7976
rect 8352 8004 8358 8016
rect 9582 8004 9588 8016
rect 8352 7976 9588 8004
rect 8352 7964 8358 7976
rect 9582 7964 9588 7976
rect 9640 7964 9646 8016
rect 11422 8004 11428 8016
rect 11383 7976 11428 8004
rect 11422 7964 11428 7976
rect 11480 7964 11486 8016
rect 11606 8004 11612 8016
rect 11567 7976 11612 8004
rect 11606 7964 11612 7976
rect 11664 7964 11670 8016
rect 11698 7964 11704 8016
rect 11756 8004 11762 8016
rect 13081 8007 13139 8013
rect 11756 7976 11801 8004
rect 11756 7964 11762 7976
rect 13081 7973 13093 8007
rect 13127 8004 13139 8007
rect 13722 8004 13728 8016
rect 13127 7976 13728 8004
rect 13127 7973 13139 7976
rect 13081 7967 13139 7973
rect 13722 7964 13728 7976
rect 13780 7964 13786 8016
rect 13817 8007 13875 8013
rect 13817 7973 13829 8007
rect 13863 8004 13875 8007
rect 13906 8004 13912 8016
rect 13863 7976 13912 8004
rect 13863 7973 13875 7976
rect 13817 7967 13875 7973
rect 13906 7964 13912 7976
rect 13964 7964 13970 8016
rect 14642 8004 14648 8016
rect 14555 7976 14648 8004
rect 14642 7964 14648 7976
rect 14700 8004 14706 8016
rect 17696 8004 17724 8035
rect 14700 7976 17724 8004
rect 14700 7964 14706 7976
rect 4614 7896 4620 7948
rect 4672 7936 4678 7948
rect 5166 7945 5172 7948
rect 5149 7939 5172 7945
rect 5149 7936 5161 7939
rect 4672 7908 5161 7936
rect 4672 7896 4678 7908
rect 5149 7905 5161 7908
rect 5224 7936 5230 7948
rect 7837 7939 7895 7945
rect 5224 7908 5297 7936
rect 5149 7899 5172 7905
rect 5166 7896 5172 7899
rect 5224 7896 5230 7908
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 8202 7936 8208 7948
rect 7883 7908 8208 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7936 9735 7939
rect 9766 7936 9772 7948
rect 9723 7908 9772 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 12986 7896 12992 7948
rect 13044 7936 13050 7948
rect 15378 7936 15384 7948
rect 13044 7908 15384 7936
rect 13044 7896 13050 7908
rect 15378 7896 15384 7908
rect 15436 7896 15442 7948
rect 16114 7896 16120 7948
rect 16172 7936 16178 7948
rect 16301 7939 16359 7945
rect 16301 7936 16313 7939
rect 16172 7908 16313 7936
rect 16172 7896 16178 7908
rect 16301 7905 16313 7908
rect 16347 7936 16359 7939
rect 16390 7936 16396 7948
rect 16347 7908 16396 7936
rect 16347 7905 16359 7908
rect 16301 7899 16359 7905
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 16574 7945 16580 7948
rect 16568 7936 16580 7945
rect 16535 7908 16580 7936
rect 16568 7899 16580 7908
rect 16574 7896 16580 7899
rect 16632 7896 16638 7948
rect 2958 7868 2964 7880
rect 2919 7840 2964 7868
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 3050 7828 3056 7880
rect 3108 7868 3114 7880
rect 4890 7868 4896 7880
rect 3108 7840 3153 7868
rect 4851 7840 4896 7868
rect 3108 7828 3114 7840
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 8110 7868 8116 7880
rect 8071 7840 8116 7868
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7868 10011 7871
rect 10042 7868 10048 7880
rect 9999 7840 10048 7868
rect 9999 7837 10011 7840
rect 9953 7831 10011 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 13630 7868 13636 7880
rect 13591 7840 13636 7868
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 14918 7868 14924 7880
rect 14879 7840 14924 7868
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 6730 7760 6736 7812
rect 6788 7800 6794 7812
rect 7561 7803 7619 7809
rect 7561 7800 7573 7803
rect 6788 7772 7573 7800
rect 6788 7760 6794 7772
rect 7561 7769 7573 7772
rect 7607 7769 7619 7803
rect 7561 7763 7619 7769
rect 12529 7803 12587 7809
rect 12529 7769 12541 7803
rect 12575 7800 12587 7803
rect 13446 7800 13452 7812
rect 12575 7772 13452 7800
rect 12575 7769 12587 7772
rect 12529 7763 12587 7769
rect 13446 7760 13452 7772
rect 13504 7760 13510 7812
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7732 1823 7735
rect 2130 7732 2136 7744
rect 1811 7704 2136 7732
rect 1811 7701 1823 7704
rect 1765 7695 1823 7701
rect 2130 7692 2136 7704
rect 2188 7692 2194 7744
rect 2498 7732 2504 7744
rect 2459 7704 2504 7732
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 5258 7692 5264 7744
rect 5316 7732 5322 7744
rect 6917 7735 6975 7741
rect 6917 7732 6929 7735
rect 5316 7704 6929 7732
rect 5316 7692 5322 7704
rect 6917 7701 6929 7704
rect 6963 7732 6975 7735
rect 7006 7732 7012 7744
rect 6963 7704 7012 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7285 7735 7343 7741
rect 7285 7701 7297 7735
rect 7331 7732 7343 7735
rect 7466 7732 7472 7744
rect 7331 7704 7472 7732
rect 7331 7701 7343 7704
rect 7285 7695 7343 7701
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 9306 7732 9312 7744
rect 9267 7704 9312 7732
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 11149 7735 11207 7741
rect 11149 7701 11161 7735
rect 11195 7732 11207 7735
rect 11238 7732 11244 7744
rect 11195 7704 11244 7732
rect 11195 7701 11207 7704
rect 11149 7695 11207 7701
rect 11238 7692 11244 7704
rect 11296 7732 11302 7744
rect 12069 7735 12127 7741
rect 12069 7732 12081 7735
rect 11296 7704 12081 7732
rect 11296 7692 11302 7704
rect 12069 7701 12081 7704
rect 12115 7701 12127 7735
rect 13262 7732 13268 7744
rect 13223 7704 13268 7732
rect 12069 7695 12127 7701
rect 13262 7692 13268 7704
rect 13320 7692 13326 7744
rect 15838 7732 15844 7744
rect 15799 7704 15844 7732
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 16114 7732 16120 7744
rect 16075 7704 16120 7732
rect 16114 7692 16120 7704
rect 16172 7692 16178 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1765 7531 1823 7537
rect 1765 7497 1777 7531
rect 1811 7528 1823 7531
rect 2958 7528 2964 7540
rect 1811 7500 2964 7528
rect 1811 7497 1823 7500
rect 1765 7491 1823 7497
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 4614 7528 4620 7540
rect 3191 7500 4620 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 4706 7488 4712 7540
rect 4764 7528 4770 7540
rect 4801 7531 4859 7537
rect 4801 7528 4813 7531
rect 4764 7500 4813 7528
rect 4764 7488 4770 7500
rect 4801 7497 4813 7500
rect 4847 7497 4859 7531
rect 4801 7491 4859 7497
rect 5077 7531 5135 7537
rect 5077 7497 5089 7531
rect 5123 7528 5135 7531
rect 5442 7528 5448 7540
rect 5123 7500 5448 7528
rect 5123 7497 5135 7500
rect 5077 7491 5135 7497
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 6089 7531 6147 7537
rect 6089 7497 6101 7531
rect 6135 7528 6147 7531
rect 6270 7528 6276 7540
rect 6135 7500 6276 7528
rect 6135 7497 6147 7500
rect 6089 7491 6147 7497
rect 6270 7488 6276 7500
rect 6328 7528 6334 7540
rect 6822 7528 6828 7540
rect 6328 7500 6828 7528
rect 6328 7488 6334 7500
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 7837 7531 7895 7537
rect 7837 7528 7849 7531
rect 7156 7500 7849 7528
rect 7156 7488 7162 7500
rect 7837 7497 7849 7500
rect 7883 7528 7895 7531
rect 8110 7528 8116 7540
rect 7883 7500 8116 7528
rect 7883 7497 7895 7500
rect 7837 7491 7895 7497
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8294 7528 8300 7540
rect 8255 7500 8300 7528
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 10229 7531 10287 7537
rect 10229 7497 10241 7531
rect 10275 7528 10287 7531
rect 11422 7528 11428 7540
rect 10275 7500 11428 7528
rect 10275 7497 10287 7500
rect 10229 7491 10287 7497
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 11698 7488 11704 7540
rect 11756 7528 11762 7540
rect 12069 7531 12127 7537
rect 12069 7528 12081 7531
rect 11756 7500 12081 7528
rect 11756 7488 11762 7500
rect 12069 7497 12081 7500
rect 12115 7497 12127 7531
rect 12069 7491 12127 7497
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 14001 7531 14059 7537
rect 14001 7528 14013 7531
rect 13780 7500 14013 7528
rect 13780 7488 13786 7500
rect 14001 7497 14013 7500
rect 14047 7497 14059 7531
rect 17586 7528 17592 7540
rect 17547 7500 17592 7528
rect 14001 7491 14059 7497
rect 17586 7488 17592 7500
rect 17644 7488 17650 7540
rect 3326 7460 3332 7472
rect 3287 7432 3332 7460
rect 3326 7420 3332 7432
rect 3384 7420 3390 7472
rect 4525 7463 4583 7469
rect 4525 7429 4537 7463
rect 4571 7460 4583 7463
rect 6178 7460 6184 7472
rect 4571 7432 6184 7460
rect 4571 7429 4583 7432
rect 4525 7423 4583 7429
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7392 3847 7395
rect 4062 7392 4068 7404
rect 3835 7364 4068 7392
rect 3835 7361 3847 7364
rect 3789 7355 3847 7361
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 5552 7401 5580 7432
rect 6178 7420 6184 7432
rect 6236 7460 6242 7472
rect 6454 7460 6460 7472
rect 6236 7432 6460 7460
rect 6236 7420 6242 7432
rect 6454 7420 6460 7432
rect 6512 7420 6518 7472
rect 6917 7463 6975 7469
rect 6917 7429 6929 7463
rect 6963 7460 6975 7463
rect 7558 7460 7564 7472
rect 6963 7432 7564 7460
rect 6963 7429 6975 7432
rect 6917 7423 6975 7429
rect 7558 7420 7564 7432
rect 7616 7420 7622 7472
rect 9217 7463 9275 7469
rect 9217 7429 9229 7463
rect 9263 7460 9275 7463
rect 9582 7460 9588 7472
rect 9263 7432 9588 7460
rect 9263 7429 9275 7432
rect 9217 7423 9275 7429
rect 9582 7420 9588 7432
rect 9640 7420 9646 7472
rect 10778 7460 10784 7472
rect 10739 7432 10784 7460
rect 10778 7420 10784 7432
rect 10836 7420 10842 7472
rect 11606 7420 11612 7472
rect 11664 7460 11670 7472
rect 11793 7463 11851 7469
rect 11793 7460 11805 7463
rect 11664 7432 11805 7460
rect 11664 7420 11670 7432
rect 11793 7429 11805 7432
rect 11839 7429 11851 7463
rect 11793 7423 11851 7429
rect 13906 7420 13912 7472
rect 13964 7460 13970 7472
rect 14921 7463 14979 7469
rect 14921 7460 14933 7463
rect 13964 7432 14933 7460
rect 13964 7420 13970 7432
rect 14921 7429 14933 7432
rect 14967 7429 14979 7463
rect 15562 7460 15568 7472
rect 15523 7432 15568 7460
rect 14921 7423 14979 7429
rect 15562 7420 15568 7432
rect 15620 7420 15626 7472
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7392 5687 7395
rect 6086 7392 6092 7404
rect 5675 7364 6092 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 6086 7352 6092 7364
rect 6144 7392 6150 7404
rect 6638 7392 6644 7404
rect 6144 7364 6644 7392
rect 6144 7352 6150 7364
rect 6638 7352 6644 7364
rect 6696 7352 6702 7404
rect 7466 7392 7472 7404
rect 7427 7364 7472 7392
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 11238 7392 11244 7404
rect 11199 7364 11244 7392
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 11333 7395 11391 7401
rect 11333 7361 11345 7395
rect 11379 7392 11391 7395
rect 12250 7392 12256 7404
rect 11379 7364 12256 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 2314 7284 2320 7336
rect 2372 7324 2378 7336
rect 3881 7327 3939 7333
rect 2372 7296 2417 7324
rect 2372 7284 2378 7296
rect 3881 7293 3893 7327
rect 3927 7324 3939 7327
rect 3970 7324 3976 7336
rect 3927 7296 3976 7324
rect 3927 7293 3939 7296
rect 3881 7287 3939 7293
rect 3970 7284 3976 7296
rect 4028 7284 4034 7336
rect 4890 7284 4896 7336
rect 4948 7324 4954 7336
rect 6178 7324 6184 7336
rect 4948 7296 6184 7324
rect 4948 7284 4954 7296
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 7193 7327 7251 7333
rect 7193 7324 7205 7327
rect 7064 7296 7205 7324
rect 7064 7284 7070 7296
rect 7193 7293 7205 7296
rect 7239 7293 7251 7327
rect 7193 7287 7251 7293
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7324 8723 7327
rect 10597 7327 10655 7333
rect 8711 7296 9812 7324
rect 8711 7293 8723 7296
rect 8665 7287 8723 7293
rect 2038 7256 2044 7268
rect 1999 7228 2044 7256
rect 2038 7216 2044 7228
rect 2096 7216 2102 7268
rect 2130 7216 2136 7268
rect 2188 7256 2194 7268
rect 2225 7259 2283 7265
rect 2225 7256 2237 7259
rect 2188 7228 2237 7256
rect 2188 7216 2194 7228
rect 2225 7225 2237 7228
rect 2271 7256 2283 7259
rect 7098 7256 7104 7268
rect 2271 7228 7104 7256
rect 2271 7225 2283 7228
rect 2225 7219 2283 7225
rect 7098 7216 7104 7228
rect 7156 7216 7162 7268
rect 9490 7256 9496 7268
rect 9451 7228 9496 7256
rect 9490 7216 9496 7228
rect 9548 7216 9554 7268
rect 9784 7265 9812 7296
rect 10597 7293 10609 7327
rect 10643 7324 10655 7327
rect 11348 7324 11376 7355
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12526 7352 12532 7404
rect 12584 7392 12590 7404
rect 12621 7395 12679 7401
rect 12621 7392 12633 7395
rect 12584 7364 12633 7392
rect 12584 7352 12590 7364
rect 12621 7361 12633 7364
rect 12667 7361 12679 7395
rect 14458 7392 14464 7404
rect 12621 7355 12679 7361
rect 14292 7364 14464 7392
rect 10643 7296 11376 7324
rect 10643 7293 10655 7296
rect 10597 7287 10655 7293
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12400 7296 12449 7324
rect 12400 7284 12406 7296
rect 12437 7293 12449 7296
rect 12483 7324 12495 7327
rect 13262 7324 13268 7336
rect 12483 7296 13268 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 13262 7284 13268 7296
rect 13320 7284 13326 7336
rect 14292 7333 14320 7364
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 14553 7395 14611 7401
rect 14553 7361 14565 7395
rect 14599 7392 14611 7395
rect 14642 7392 14648 7404
rect 14599 7364 14648 7392
rect 14599 7361 14611 7364
rect 14553 7355 14611 7361
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 16025 7395 16083 7401
rect 16025 7361 16037 7395
rect 16071 7392 16083 7395
rect 16114 7392 16120 7404
rect 16071 7364 16120 7392
rect 16071 7361 16083 7364
rect 16025 7355 16083 7361
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 13633 7327 13691 7333
rect 13633 7293 13645 7327
rect 13679 7324 13691 7327
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 13679 7296 14289 7324
rect 13679 7293 13691 7296
rect 13633 7287 13691 7293
rect 14277 7293 14289 7296
rect 14323 7293 14335 7327
rect 19058 7324 19064 7336
rect 14277 7287 14335 7293
rect 15764 7296 19064 7324
rect 9769 7259 9827 7265
rect 9769 7225 9781 7259
rect 9815 7256 9827 7259
rect 10686 7256 10692 7268
rect 9815 7228 10692 7256
rect 9815 7225 9827 7228
rect 9769 7219 9827 7225
rect 10686 7216 10692 7228
rect 10744 7216 10750 7268
rect 11146 7216 11152 7268
rect 11204 7256 11210 7268
rect 11241 7259 11299 7265
rect 11241 7256 11253 7259
rect 11204 7228 11253 7256
rect 11204 7216 11210 7228
rect 11241 7225 11253 7228
rect 11287 7225 11299 7259
rect 11241 7219 11299 7225
rect 13449 7259 13507 7265
rect 13449 7225 13461 7259
rect 13495 7256 13507 7259
rect 15764 7256 15792 7296
rect 19058 7284 19064 7296
rect 19116 7284 19122 7336
rect 13495 7228 14412 7256
rect 13495 7225 13507 7228
rect 13449 7219 13507 7225
rect 2774 7188 2780 7200
rect 2735 7160 2780 7188
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 3789 7191 3847 7197
rect 3789 7157 3801 7191
rect 3835 7188 3847 7191
rect 4062 7188 4068 7200
rect 3835 7160 4068 7188
rect 3835 7157 3847 7160
rect 3789 7151 3847 7157
rect 4062 7148 4068 7160
rect 4120 7148 4126 7200
rect 4706 7148 4712 7200
rect 4764 7188 4770 7200
rect 5537 7191 5595 7197
rect 5537 7188 5549 7191
rect 4764 7160 5549 7188
rect 4764 7148 4770 7160
rect 5537 7157 5549 7160
rect 5583 7157 5595 7191
rect 5537 7151 5595 7157
rect 6270 7148 6276 7200
rect 6328 7188 6334 7200
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 6328 7160 6561 7188
rect 6328 7148 6334 7160
rect 6549 7157 6561 7160
rect 6595 7188 6607 7191
rect 7377 7191 7435 7197
rect 7377 7188 7389 7191
rect 6595 7160 7389 7188
rect 6595 7157 6607 7160
rect 6549 7151 6607 7157
rect 7377 7157 7389 7160
rect 7423 7188 7435 7191
rect 7926 7188 7932 7200
rect 7423 7160 7932 7188
rect 7423 7157 7435 7160
rect 7377 7151 7435 7157
rect 7926 7148 7932 7160
rect 7984 7148 7990 7200
rect 9033 7191 9091 7197
rect 9033 7157 9045 7191
rect 9079 7188 9091 7191
rect 9677 7191 9735 7197
rect 9677 7188 9689 7191
rect 9079 7160 9689 7188
rect 9079 7157 9091 7160
rect 9033 7151 9091 7157
rect 9677 7157 9689 7160
rect 9723 7188 9735 7191
rect 9858 7188 9864 7200
rect 9723 7160 9864 7188
rect 9723 7157 9735 7160
rect 9677 7151 9735 7157
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 13633 7191 13691 7197
rect 13633 7188 13645 7191
rect 13228 7160 13645 7188
rect 13228 7148 13234 7160
rect 13633 7157 13645 7160
rect 13679 7188 13691 7191
rect 13725 7191 13783 7197
rect 13725 7188 13737 7191
rect 13679 7160 13737 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 13725 7157 13737 7160
rect 13771 7157 13783 7191
rect 14384 7188 14412 7228
rect 15304 7228 15792 7256
rect 14461 7191 14519 7197
rect 14461 7188 14473 7191
rect 14384 7160 14473 7188
rect 13725 7151 13783 7157
rect 14461 7157 14473 7160
rect 14507 7188 14519 7191
rect 14826 7188 14832 7200
rect 14507 7160 14832 7188
rect 14507 7157 14519 7160
rect 14461 7151 14519 7157
rect 14826 7148 14832 7160
rect 14884 7188 14890 7200
rect 15304 7188 15332 7228
rect 15838 7216 15844 7268
rect 15896 7256 15902 7268
rect 16025 7259 16083 7265
rect 16025 7256 16037 7259
rect 15896 7228 16037 7256
rect 15896 7216 15902 7228
rect 16025 7225 16037 7228
rect 16071 7225 16083 7259
rect 16025 7219 16083 7225
rect 16117 7259 16175 7265
rect 16117 7225 16129 7259
rect 16163 7256 16175 7259
rect 16574 7256 16580 7268
rect 16163 7228 16580 7256
rect 16163 7225 16175 7228
rect 16117 7219 16175 7225
rect 14884 7160 15332 7188
rect 15381 7191 15439 7197
rect 14884 7148 14890 7160
rect 15381 7157 15393 7191
rect 15427 7188 15439 7191
rect 16132 7188 16160 7219
rect 16574 7216 16580 7228
rect 16632 7256 16638 7268
rect 18046 7256 18052 7268
rect 16632 7228 16988 7256
rect 18007 7228 18052 7256
rect 16632 7216 16638 7228
rect 16960 7200 16988 7228
rect 18046 7216 18052 7228
rect 18104 7216 18110 7268
rect 15427 7160 16160 7188
rect 15427 7157 15439 7160
rect 15381 7151 15439 7157
rect 16390 7148 16396 7200
rect 16448 7188 16454 7200
rect 16485 7191 16543 7197
rect 16485 7188 16497 7191
rect 16448 7160 16497 7188
rect 16448 7148 16454 7160
rect 16485 7157 16497 7160
rect 16531 7188 16543 7191
rect 16758 7188 16764 7200
rect 16531 7160 16764 7188
rect 16531 7157 16543 7160
rect 16485 7151 16543 7157
rect 16758 7148 16764 7160
rect 16816 7148 16822 7200
rect 16942 7188 16948 7200
rect 16903 7160 16948 7188
rect 16942 7148 16948 7160
rect 17000 7148 17006 7200
rect 17218 7188 17224 7200
rect 17179 7160 17224 7188
rect 17218 7148 17224 7160
rect 17276 7148 17282 7200
rect 18506 7188 18512 7200
rect 18467 7160 18512 7188
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2314 6984 2320 6996
rect 2275 6956 2320 6984
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 2961 6987 3019 6993
rect 2961 6984 2973 6987
rect 2924 6956 2973 6984
rect 2924 6944 2930 6956
rect 2961 6953 2973 6956
rect 3007 6953 3019 6987
rect 2961 6947 3019 6953
rect 3602 6944 3608 6996
rect 3660 6944 3666 6996
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 6086 6984 6092 6996
rect 4028 6956 4364 6984
rect 6047 6956 6092 6984
rect 4028 6944 4034 6956
rect 3234 6876 3240 6928
rect 3292 6916 3298 6928
rect 3620 6916 3648 6944
rect 4336 6925 4364 6956
rect 6086 6944 6092 6956
rect 6144 6944 6150 6996
rect 7374 6984 7380 6996
rect 7335 6956 7380 6984
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 7929 6987 7987 6993
rect 7929 6953 7941 6987
rect 7975 6984 7987 6987
rect 8202 6984 8208 6996
rect 7975 6956 8208 6984
rect 7975 6953 7987 6956
rect 7929 6947 7987 6953
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 9217 6987 9275 6993
rect 9217 6953 9229 6987
rect 9263 6984 9275 6987
rect 9490 6984 9496 6996
rect 9263 6956 9496 6984
rect 9263 6953 9275 6956
rect 9217 6947 9275 6953
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 9766 6944 9772 6996
rect 9824 6984 9830 6996
rect 10413 6987 10471 6993
rect 10413 6984 10425 6987
rect 9824 6956 10425 6984
rect 9824 6944 9830 6956
rect 10413 6953 10425 6956
rect 10459 6953 10471 6987
rect 14642 6984 14648 6996
rect 14603 6956 14648 6984
rect 10413 6947 10471 6953
rect 14642 6944 14648 6956
rect 14700 6944 14706 6996
rect 16942 6944 16948 6996
rect 17000 6984 17006 6996
rect 17773 6987 17831 6993
rect 17773 6984 17785 6987
rect 17000 6956 17785 6984
rect 17000 6944 17006 6956
rect 17773 6953 17785 6956
rect 17819 6953 17831 6987
rect 17773 6947 17831 6953
rect 3292 6888 3648 6916
rect 4321 6919 4379 6925
rect 3292 6876 3298 6888
rect 4321 6885 4333 6919
rect 4367 6885 4379 6919
rect 7193 6919 7251 6925
rect 7193 6916 7205 6919
rect 4321 6879 4379 6885
rect 6196 6888 7205 6916
rect 3050 6808 3056 6860
rect 3108 6848 3114 6860
rect 3513 6851 3571 6857
rect 3513 6848 3525 6851
rect 3108 6820 3525 6848
rect 3108 6808 3114 6820
rect 3513 6817 3525 6820
rect 3559 6848 3571 6851
rect 3602 6848 3608 6860
rect 3559 6820 3608 6848
rect 3559 6817 3571 6820
rect 3513 6811 3571 6817
rect 3602 6808 3608 6820
rect 3660 6808 3666 6860
rect 6196 6848 6224 6888
rect 7193 6885 7205 6888
rect 7239 6916 7251 6919
rect 8846 6916 8852 6928
rect 7239 6888 8852 6916
rect 7239 6885 7251 6888
rect 7193 6879 7251 6885
rect 8846 6876 8852 6888
rect 8904 6876 8910 6928
rect 11609 6919 11667 6925
rect 11609 6885 11621 6919
rect 11655 6885 11667 6919
rect 11609 6879 11667 6885
rect 3988 6820 6224 6848
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6780 1455 6783
rect 2222 6780 2228 6792
rect 1443 6752 2228 6780
rect 1443 6749 1455 6752
rect 1397 6743 1455 6749
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 2961 6783 3019 6789
rect 2961 6749 2973 6783
rect 3007 6780 3019 6783
rect 3142 6780 3148 6792
rect 3007 6752 3148 6780
rect 3007 6749 3019 6752
rect 2961 6743 3019 6749
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 3988 6780 4016 6820
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 7469 6851 7527 6857
rect 7469 6848 7481 6851
rect 6880 6820 7481 6848
rect 6880 6808 6886 6820
rect 7469 6817 7481 6820
rect 7515 6817 7527 6851
rect 7469 6811 7527 6817
rect 8389 6851 8447 6857
rect 8389 6817 8401 6851
rect 8435 6848 8447 6851
rect 9030 6848 9036 6860
rect 8435 6820 9036 6848
rect 8435 6817 8447 6820
rect 8389 6811 8447 6817
rect 9030 6808 9036 6820
rect 9088 6808 9094 6860
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6817 9735 6851
rect 10962 6848 10968 6860
rect 10923 6820 10968 6848
rect 9677 6811 9735 6817
rect 3528 6752 4016 6780
rect 4065 6783 4123 6789
rect 2501 6715 2559 6721
rect 2501 6681 2513 6715
rect 2547 6712 2559 6715
rect 3528 6712 3556 6752
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 8294 6780 8300 6792
rect 8255 6752 8300 6780
rect 4065 6743 4123 6749
rect 2547 6684 3556 6712
rect 2547 6681 2559 6684
rect 2501 6675 2559 6681
rect 3602 6672 3608 6724
rect 3660 6712 3666 6724
rect 4080 6712 4108 6743
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 6365 6715 6423 6721
rect 6365 6712 6377 6715
rect 3660 6684 4108 6712
rect 5000 6684 6377 6712
rect 3660 6672 3666 6684
rect 1949 6647 2007 6653
rect 1949 6613 1961 6647
rect 1995 6644 2007 6647
rect 2038 6644 2044 6656
rect 1995 6616 2044 6644
rect 1995 6613 2007 6616
rect 1949 6607 2007 6613
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 3881 6647 3939 6653
rect 3881 6613 3893 6647
rect 3927 6644 3939 6647
rect 3970 6644 3976 6656
rect 3927 6616 3976 6644
rect 3927 6613 3939 6616
rect 3881 6607 3939 6613
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 5000 6644 5028 6684
rect 6365 6681 6377 6684
rect 6411 6681 6423 6715
rect 6365 6675 6423 6681
rect 9490 6672 9496 6724
rect 9548 6712 9554 6724
rect 9692 6712 9720 6811
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11422 6848 11428 6860
rect 11383 6820 11428 6848
rect 11422 6808 11428 6820
rect 11480 6808 11486 6860
rect 11624 6848 11652 6879
rect 13630 6876 13636 6928
rect 13688 6916 13694 6928
rect 13688 6888 13768 6916
rect 13688 6876 13694 6888
rect 11974 6848 11980 6860
rect 11624 6820 11980 6848
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12342 6848 12348 6860
rect 12207 6820 12348 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 12710 6808 12716 6860
rect 12768 6848 12774 6860
rect 12877 6851 12935 6857
rect 12877 6848 12889 6851
rect 12768 6820 12889 6848
rect 12768 6808 12774 6820
rect 12877 6817 12889 6820
rect 12923 6817 12935 6851
rect 13740 6848 13768 6888
rect 14182 6876 14188 6928
rect 14240 6916 14246 6928
rect 14240 6888 15332 6916
rect 14240 6876 14246 6888
rect 15304 6857 15332 6888
rect 14921 6851 14979 6857
rect 14921 6848 14933 6851
rect 13740 6820 14933 6848
rect 12877 6811 12935 6817
rect 14921 6817 14933 6820
rect 14967 6817 14979 6851
rect 14921 6811 14979 6817
rect 15289 6851 15347 6857
rect 15289 6817 15301 6851
rect 15335 6848 15347 6851
rect 15378 6848 15384 6860
rect 15335 6820 15384 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 15933 6851 15991 6857
rect 15933 6817 15945 6851
rect 15979 6848 15991 6851
rect 16482 6848 16488 6860
rect 15979 6820 16488 6848
rect 15979 6817 15991 6820
rect 15933 6811 15991 6817
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 16666 6857 16672 6860
rect 16660 6848 16672 6857
rect 16627 6820 16672 6848
rect 16660 6811 16672 6820
rect 16666 6808 16672 6811
rect 16724 6808 16730 6860
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6780 10011 6783
rect 11054 6780 11060 6792
rect 9999 6752 11060 6780
rect 9999 6749 10011 6752
rect 9953 6743 10011 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11701 6783 11759 6789
rect 11701 6749 11713 6783
rect 11747 6780 11759 6783
rect 11882 6780 11888 6792
rect 11747 6752 11888 6780
rect 11747 6749 11759 6752
rect 11701 6743 11759 6749
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 12621 6783 12679 6789
rect 12621 6780 12633 6783
rect 12452 6752 12633 6780
rect 11149 6715 11207 6721
rect 11149 6712 11161 6715
rect 9548 6684 11161 6712
rect 9548 6672 9554 6684
rect 11149 6681 11161 6684
rect 11195 6681 11207 6715
rect 11149 6675 11207 6681
rect 12452 6656 12480 6752
rect 12621 6749 12633 6752
rect 12667 6749 12679 6783
rect 12621 6743 12679 6749
rect 13998 6740 14004 6792
rect 14056 6780 14062 6792
rect 14366 6780 14372 6792
rect 14056 6752 14372 6780
rect 14056 6740 14062 6752
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 16390 6780 16396 6792
rect 16351 6752 16396 6780
rect 16390 6740 16396 6752
rect 16448 6740 16454 6792
rect 18874 6780 18880 6792
rect 18835 6752 18880 6780
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 5442 6644 5448 6656
rect 4120 6616 5028 6644
rect 5403 6616 5448 6644
rect 4120 6604 4126 6616
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 6914 6644 6920 6656
rect 6875 6616 6920 6644
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 8386 6604 8392 6656
rect 8444 6644 8450 6656
rect 8573 6647 8631 6653
rect 8573 6644 8585 6647
rect 8444 6616 8585 6644
rect 8444 6604 8450 6616
rect 8573 6613 8585 6616
rect 8619 6613 8631 6647
rect 12434 6644 12440 6656
rect 12395 6616 12440 6644
rect 8573 6607 8631 6613
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 13998 6644 14004 6656
rect 13959 6616 14004 6644
rect 13998 6604 14004 6616
rect 14056 6604 14062 6656
rect 15470 6644 15476 6656
rect 15431 6616 15476 6644
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 16301 6647 16359 6653
rect 16301 6613 16313 6647
rect 16347 6644 16359 6647
rect 16390 6644 16396 6656
rect 16347 6616 16396 6644
rect 16347 6613 16359 6616
rect 16301 6607 16359 6613
rect 16390 6604 16396 6616
rect 16448 6644 16454 6656
rect 16666 6644 16672 6656
rect 16448 6616 16672 6644
rect 16448 6604 16454 6616
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 18322 6644 18328 6656
rect 18283 6616 18328 6644
rect 18322 6604 18328 6616
rect 18380 6604 18386 6656
rect 18690 6644 18696 6656
rect 18651 6616 18696 6644
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 19334 6644 19340 6656
rect 19295 6616 19340 6644
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 3694 6400 3700 6452
rect 3752 6440 3758 6452
rect 4246 6440 4252 6452
rect 3752 6412 4252 6440
rect 3752 6400 3758 6412
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 4617 6443 4675 6449
rect 4617 6409 4629 6443
rect 4663 6440 4675 6443
rect 4890 6440 4896 6452
rect 4663 6412 4896 6440
rect 4663 6409 4675 6412
rect 4617 6403 4675 6409
rect 2590 6372 2596 6384
rect 1412 6344 2596 6372
rect 1412 6245 1440 6344
rect 2590 6332 2596 6344
rect 2648 6332 2654 6384
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 4632 6372 4660 6403
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 5166 6440 5172 6452
rect 5127 6412 5172 6440
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 8297 6443 8355 6449
rect 8297 6409 8309 6443
rect 8343 6440 8355 6443
rect 8570 6440 8576 6452
rect 8343 6412 8576 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 3660 6344 4660 6372
rect 6917 6375 6975 6381
rect 3660 6332 3666 6344
rect 6917 6341 6929 6375
rect 6963 6372 6975 6375
rect 8018 6372 8024 6384
rect 6963 6344 8024 6372
rect 6963 6341 6975 6344
rect 6917 6335 6975 6341
rect 8018 6332 8024 6344
rect 8076 6332 8082 6384
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6205 1455 6239
rect 1397 6199 1455 6205
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 2547 6208 2605 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 2593 6205 2605 6208
rect 2639 6236 2651 6239
rect 3620 6236 3648 6332
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 5721 6307 5779 6313
rect 5721 6304 5733 6307
rect 5592 6276 5733 6304
rect 5592 6264 5598 6276
rect 5721 6273 5733 6276
rect 5767 6273 5779 6307
rect 5721 6267 5779 6273
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 6687 6276 7481 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 7469 6273 7481 6276
rect 7515 6304 7527 6307
rect 8202 6304 8208 6316
rect 7515 6276 8208 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 8404 6313 8432 6412
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 9732 6412 10517 6440
rect 9732 6400 9738 6412
rect 10505 6409 10517 6412
rect 10551 6440 10563 6443
rect 11422 6440 11428 6452
rect 10551 6412 11428 6440
rect 10551 6409 10563 6412
rect 10505 6403 10563 6409
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 13817 6443 13875 6449
rect 13817 6440 13829 6443
rect 12768 6412 13829 6440
rect 12768 6400 12774 6412
rect 13817 6409 13829 6412
rect 13863 6440 13875 6443
rect 14369 6443 14427 6449
rect 14369 6440 14381 6443
rect 13863 6412 14381 6440
rect 13863 6409 13875 6412
rect 13817 6403 13875 6409
rect 14369 6409 14381 6412
rect 14415 6409 14427 6443
rect 15378 6440 15384 6452
rect 15339 6412 15384 6440
rect 14369 6403 14427 6409
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 15746 6440 15752 6452
rect 15707 6412 15752 6440
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 15933 6443 15991 6449
rect 15933 6409 15945 6443
rect 15979 6440 15991 6443
rect 16114 6440 16120 6452
rect 15979 6412 16120 6440
rect 15979 6409 15991 6412
rect 15933 6403 15991 6409
rect 16114 6400 16120 6412
rect 16172 6400 16178 6452
rect 16758 6400 16764 6452
rect 16816 6440 16822 6452
rect 16853 6443 16911 6449
rect 16853 6440 16865 6443
rect 16816 6412 16865 6440
rect 16816 6400 16822 6412
rect 16853 6409 16865 6412
rect 16899 6440 16911 6443
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 16899 6412 17785 6440
rect 16899 6409 16911 6412
rect 16853 6403 16911 6409
rect 17773 6409 17785 6412
rect 17819 6409 17831 6443
rect 17773 6403 17831 6409
rect 10965 6375 11023 6381
rect 10965 6341 10977 6375
rect 11011 6372 11023 6375
rect 11974 6372 11980 6384
rect 11011 6344 11980 6372
rect 11011 6341 11023 6344
rect 10965 6335 11023 6341
rect 11974 6332 11980 6344
rect 12032 6332 12038 6384
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 11238 6304 11244 6316
rect 11199 6276 11244 6304
rect 8389 6267 8447 6273
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 16393 6307 16451 6313
rect 16393 6273 16405 6307
rect 16439 6304 16451 6307
rect 16482 6304 16488 6316
rect 16439 6276 16488 6304
rect 16439 6273 16451 6276
rect 16393 6267 16451 6273
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 17788 6304 17816 6403
rect 18046 6304 18052 6316
rect 17788 6276 18052 6304
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 2639 6208 3648 6236
rect 2639 6205 2651 6208
rect 2593 6199 2651 6205
rect 4890 6196 4896 6248
rect 4948 6236 4954 6248
rect 7742 6236 7748 6248
rect 4948 6208 7748 6236
rect 4948 6196 4954 6208
rect 7742 6196 7748 6208
rect 7800 6196 7806 6248
rect 10962 6196 10968 6248
rect 11020 6236 11026 6248
rect 11057 6239 11115 6245
rect 11057 6236 11069 6239
rect 11020 6208 11069 6236
rect 11020 6196 11026 6208
rect 11057 6205 11069 6208
rect 11103 6205 11115 6239
rect 12434 6236 12440 6248
rect 11057 6199 11115 6205
rect 12176 6208 12440 6236
rect 2133 6171 2191 6177
rect 2133 6137 2145 6171
rect 2179 6168 2191 6171
rect 2860 6171 2918 6177
rect 2860 6168 2872 6171
rect 2179 6140 2872 6168
rect 2179 6137 2191 6140
rect 2133 6131 2191 6137
rect 2860 6137 2872 6140
rect 2906 6168 2918 6171
rect 3602 6168 3608 6180
rect 2906 6140 3608 6168
rect 2906 6137 2918 6140
rect 2860 6131 2918 6137
rect 3602 6128 3608 6140
rect 3660 6128 3666 6180
rect 5074 6128 5080 6180
rect 5132 6168 5138 6180
rect 5445 6171 5503 6177
rect 5445 6168 5457 6171
rect 5132 6140 5457 6168
rect 5132 6128 5138 6140
rect 5445 6137 5457 6140
rect 5491 6137 5503 6171
rect 5445 6131 5503 6137
rect 6273 6171 6331 6177
rect 6273 6137 6285 6171
rect 6319 6168 6331 6171
rect 6822 6168 6828 6180
rect 6319 6140 6828 6168
rect 6319 6137 6331 6140
rect 6273 6131 6331 6137
rect 6822 6128 6828 6140
rect 6880 6128 6886 6180
rect 7190 6168 7196 6180
rect 7151 6140 7196 6168
rect 7190 6128 7196 6140
rect 7248 6128 7254 6180
rect 7374 6168 7380 6180
rect 7335 6140 7380 6168
rect 7374 6128 7380 6140
rect 7432 6128 7438 6180
rect 8634 6171 8692 6177
rect 8634 6168 8646 6171
rect 7852 6140 8646 6168
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 3970 6100 3976 6112
rect 3931 6072 3976 6100
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 4985 6103 5043 6109
rect 4985 6069 4997 6103
rect 5031 6100 5043 6103
rect 5629 6103 5687 6109
rect 5629 6100 5641 6103
rect 5031 6072 5641 6100
rect 5031 6069 5043 6072
rect 4985 6063 5043 6069
rect 5629 6069 5641 6072
rect 5675 6100 5687 6103
rect 6454 6100 6460 6112
rect 5675 6072 6460 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 6454 6060 6460 6072
rect 6512 6100 6518 6112
rect 6638 6100 6644 6112
rect 6512 6072 6644 6100
rect 6512 6060 6518 6072
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 7852 6109 7880 6140
rect 8634 6137 8646 6140
rect 8680 6137 8692 6171
rect 8634 6131 8692 6137
rect 10870 6128 10876 6180
rect 10928 6168 10934 6180
rect 12176 6177 12204 6208
rect 12434 6196 12440 6208
rect 12492 6196 12498 6248
rect 12161 6171 12219 6177
rect 12161 6168 12173 6171
rect 10928 6140 12173 6168
rect 10928 6128 10934 6140
rect 12161 6137 12173 6140
rect 12207 6137 12219 6171
rect 12161 6131 12219 6137
rect 12342 6128 12348 6180
rect 12400 6168 12406 6180
rect 12682 6171 12740 6177
rect 12682 6168 12694 6171
rect 12400 6140 12694 6168
rect 12400 6128 12406 6140
rect 12682 6137 12694 6140
rect 12728 6137 12740 6171
rect 12682 6131 12740 6137
rect 15013 6171 15071 6177
rect 15013 6137 15025 6171
rect 15059 6168 15071 6171
rect 16482 6168 16488 6180
rect 15059 6140 16488 6168
rect 15059 6137 15071 6140
rect 15013 6131 15071 6137
rect 16482 6128 16488 6140
rect 16540 6128 16546 6180
rect 18294 6171 18352 6177
rect 18294 6168 18306 6171
rect 17420 6140 18306 6168
rect 17420 6112 17448 6140
rect 18294 6137 18306 6140
rect 18340 6168 18352 6171
rect 18966 6168 18972 6180
rect 18340 6140 18972 6168
rect 18340 6137 18352 6140
rect 18294 6131 18352 6137
rect 18966 6128 18972 6140
rect 19024 6128 19030 6180
rect 7837 6103 7895 6109
rect 7837 6100 7849 6103
rect 7340 6072 7849 6100
rect 7340 6060 7346 6072
rect 7837 6069 7849 6072
rect 7883 6069 7895 6103
rect 7837 6063 7895 6069
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 9769 6103 9827 6109
rect 9769 6100 9781 6103
rect 9732 6072 9781 6100
rect 9732 6060 9738 6072
rect 9769 6069 9781 6072
rect 9815 6069 9827 6103
rect 11882 6100 11888 6112
rect 11843 6072 11888 6100
rect 9769 6063 9827 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 15746 6060 15752 6112
rect 15804 6100 15810 6112
rect 16393 6103 16451 6109
rect 16393 6100 16405 6103
rect 15804 6072 16405 6100
rect 15804 6060 15810 6072
rect 16393 6069 16405 6072
rect 16439 6069 16451 6103
rect 17402 6100 17408 6112
rect 17363 6072 17408 6100
rect 16393 6063 16451 6069
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 19426 6100 19432 6112
rect 19387 6072 19432 6100
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 3510 5896 3516 5908
rect 3471 5868 3516 5896
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3660 5868 3893 5896
rect 3660 5856 3666 5868
rect 3881 5865 3893 5868
rect 3927 5896 3939 5899
rect 5074 5896 5080 5908
rect 3927 5868 4752 5896
rect 5035 5868 5080 5896
rect 3927 5865 3939 5868
rect 3881 5859 3939 5865
rect 4724 5840 4752 5868
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 5534 5896 5540 5908
rect 5495 5868 5540 5896
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 7282 5896 7288 5908
rect 7243 5868 7288 5896
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 9490 5896 9496 5908
rect 9451 5868 9496 5896
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 12710 5856 12716 5908
rect 12768 5896 12774 5908
rect 13265 5899 13323 5905
rect 13265 5896 13277 5899
rect 12768 5868 13277 5896
rect 12768 5856 12774 5868
rect 13265 5865 13277 5868
rect 13311 5896 13323 5899
rect 15749 5899 15807 5905
rect 13311 5868 14136 5896
rect 13311 5865 13323 5868
rect 13265 5859 13323 5865
rect 2961 5831 3019 5837
rect 2961 5797 2973 5831
rect 3007 5828 3019 5831
rect 4062 5828 4068 5840
rect 3007 5800 4068 5828
rect 3007 5797 3019 5800
rect 2961 5791 3019 5797
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 4614 5828 4620 5840
rect 4575 5800 4620 5828
rect 4614 5788 4620 5800
rect 4672 5788 4678 5840
rect 4706 5788 4712 5840
rect 4764 5828 4770 5840
rect 5552 5828 5580 5856
rect 11232 5831 11290 5837
rect 4764 5800 5580 5828
rect 8404 5800 9996 5828
rect 4764 5788 4770 5800
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 2774 5760 2780 5772
rect 1912 5732 2780 5760
rect 1912 5720 1918 5732
rect 2774 5720 2780 5732
rect 2832 5760 2838 5772
rect 3053 5763 3111 5769
rect 3053 5760 3065 5763
rect 2832 5732 3065 5760
rect 2832 5720 2838 5732
rect 3053 5729 3065 5732
rect 3099 5760 3111 5763
rect 3970 5760 3976 5772
rect 3099 5732 3976 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 4430 5760 4436 5772
rect 4391 5732 4436 5760
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 5442 5760 5448 5772
rect 4540 5732 5448 5760
rect 2958 5692 2964 5704
rect 2919 5664 2964 5692
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 4246 5652 4252 5704
rect 4304 5692 4310 5704
rect 4540 5692 4568 5732
rect 5442 5720 5448 5732
rect 5500 5760 5506 5772
rect 6178 5769 6184 5772
rect 6172 5760 6184 5769
rect 5500 5732 6184 5760
rect 5500 5720 5506 5732
rect 6172 5723 6184 5732
rect 6178 5720 6184 5723
rect 6236 5720 6242 5772
rect 8404 5769 8432 5800
rect 9968 5772 9996 5800
rect 11232 5797 11244 5831
rect 11278 5828 11290 5831
rect 11422 5828 11428 5840
rect 11278 5800 11428 5828
rect 11278 5797 11290 5800
rect 11232 5791 11290 5797
rect 11422 5788 11428 5800
rect 11480 5788 11486 5840
rect 13998 5828 14004 5840
rect 13959 5800 14004 5828
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 14108 5837 14136 5868
rect 15749 5865 15761 5899
rect 15795 5896 15807 5899
rect 18966 5896 18972 5908
rect 15795 5868 16528 5896
rect 18927 5868 18972 5896
rect 15795 5865 15807 5868
rect 15749 5859 15807 5865
rect 16500 5840 16528 5868
rect 18966 5856 18972 5868
rect 19024 5856 19030 5908
rect 19518 5856 19524 5908
rect 19576 5896 19582 5908
rect 19613 5899 19671 5905
rect 19613 5896 19625 5899
rect 19576 5868 19625 5896
rect 19576 5856 19582 5868
rect 19613 5865 19625 5868
rect 19659 5865 19671 5899
rect 19613 5859 19671 5865
rect 14093 5831 14151 5837
rect 14093 5797 14105 5831
rect 14139 5797 14151 5831
rect 14093 5791 14151 5797
rect 15930 5788 15936 5840
rect 15988 5828 15994 5840
rect 16209 5831 16267 5837
rect 16209 5828 16221 5831
rect 15988 5800 16221 5828
rect 15988 5788 15994 5800
rect 16209 5797 16221 5800
rect 16255 5797 16267 5831
rect 16390 5828 16396 5840
rect 16351 5800 16396 5828
rect 16209 5791 16267 5797
rect 16390 5788 16396 5800
rect 16448 5788 16454 5840
rect 16482 5788 16488 5840
rect 16540 5828 16546 5840
rect 16540 5800 16585 5828
rect 16540 5788 16546 5800
rect 8389 5763 8447 5769
rect 8389 5729 8401 5763
rect 8435 5729 8447 5763
rect 9674 5760 9680 5772
rect 9635 5732 9680 5760
rect 8389 5723 8447 5729
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 9950 5760 9956 5772
rect 9911 5732 9956 5760
rect 9950 5720 9956 5732
rect 10008 5720 10014 5772
rect 10870 5720 10876 5772
rect 10928 5760 10934 5772
rect 10965 5763 11023 5769
rect 10965 5760 10977 5763
rect 10928 5732 10977 5760
rect 10928 5720 10934 5732
rect 10965 5729 10977 5732
rect 11011 5729 11023 5763
rect 10965 5723 11023 5729
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 14829 5763 14887 5769
rect 14829 5760 14841 5763
rect 13872 5732 14841 5760
rect 13872 5720 13878 5732
rect 14829 5729 14841 5732
rect 14875 5729 14887 5763
rect 14829 5723 14887 5729
rect 15654 5720 15660 5772
rect 15712 5760 15718 5772
rect 16408 5760 16436 5788
rect 17862 5769 17868 5772
rect 15712 5732 16436 5760
rect 17129 5763 17187 5769
rect 15712 5720 15718 5732
rect 17129 5729 17141 5763
rect 17175 5760 17187 5763
rect 17497 5763 17555 5769
rect 17497 5760 17509 5763
rect 17175 5732 17509 5760
rect 17175 5729 17187 5732
rect 17129 5723 17187 5729
rect 17497 5729 17509 5732
rect 17543 5760 17555 5763
rect 17856 5760 17868 5769
rect 17543 5732 17868 5760
rect 17543 5729 17555 5732
rect 17497 5723 17555 5729
rect 17856 5723 17868 5732
rect 17862 5720 17868 5723
rect 17920 5720 17926 5772
rect 4304 5664 4568 5692
rect 5905 5695 5963 5701
rect 4304 5652 4310 5664
rect 5905 5661 5917 5695
rect 5951 5661 5963 5695
rect 13906 5692 13912 5704
rect 13867 5664 13912 5692
rect 5905 5655 5963 5661
rect 2317 5627 2375 5633
rect 2317 5593 2329 5627
rect 2363 5624 2375 5627
rect 3050 5624 3056 5636
rect 2363 5596 3056 5624
rect 2363 5593 2375 5596
rect 2317 5587 2375 5593
rect 3050 5584 3056 5596
rect 3108 5584 3114 5636
rect 4154 5624 4160 5636
rect 4115 5596 4160 5624
rect 4154 5584 4160 5596
rect 4212 5584 4218 5636
rect 1946 5556 1952 5568
rect 1907 5528 1952 5556
rect 1946 5516 1952 5528
rect 2004 5516 2010 5568
rect 2501 5559 2559 5565
rect 2501 5525 2513 5559
rect 2547 5556 2559 5559
rect 2682 5556 2688 5568
rect 2547 5528 2688 5556
rect 2547 5525 2559 5528
rect 2501 5519 2559 5525
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 5534 5516 5540 5568
rect 5592 5556 5598 5568
rect 5920 5556 5948 5655
rect 13906 5652 13912 5664
rect 13964 5652 13970 5704
rect 17586 5692 17592 5704
rect 17547 5664 17592 5692
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 20346 5692 20352 5704
rect 20307 5664 20352 5692
rect 20346 5652 20352 5664
rect 20404 5652 20410 5704
rect 7834 5624 7840 5636
rect 7795 5596 7840 5624
rect 7834 5584 7840 5596
rect 7892 5584 7898 5636
rect 11974 5584 11980 5636
rect 12032 5624 12038 5636
rect 13541 5627 13599 5633
rect 13541 5624 13553 5627
rect 12032 5596 13553 5624
rect 12032 5584 12038 5596
rect 13541 5593 13553 5596
rect 13587 5593 13599 5627
rect 13541 5587 13599 5593
rect 14274 5584 14280 5636
rect 14332 5624 14338 5636
rect 15746 5624 15752 5636
rect 14332 5596 15752 5624
rect 14332 5584 14338 5596
rect 15746 5584 15752 5596
rect 15804 5584 15810 5636
rect 15838 5584 15844 5636
rect 15896 5624 15902 5636
rect 15933 5627 15991 5633
rect 15933 5624 15945 5627
rect 15896 5596 15945 5624
rect 15896 5584 15902 5596
rect 15933 5593 15945 5596
rect 15979 5593 15991 5627
rect 15933 5587 15991 5593
rect 6086 5556 6092 5568
rect 5592 5528 6092 5556
rect 5592 5516 5598 5528
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 8294 5556 8300 5568
rect 8255 5528 8300 5556
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8570 5556 8576 5568
rect 8531 5528 8576 5556
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 9030 5556 9036 5568
rect 8991 5528 9036 5556
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 9766 5516 9772 5568
rect 9824 5556 9830 5568
rect 10413 5559 10471 5565
rect 10413 5556 10425 5559
rect 9824 5528 10425 5556
rect 9824 5516 9830 5528
rect 10413 5525 10425 5528
rect 10459 5525 10471 5559
rect 10870 5556 10876 5568
rect 10831 5528 10876 5556
rect 10413 5519 10471 5525
rect 10870 5516 10876 5528
rect 10928 5516 10934 5568
rect 12342 5556 12348 5568
rect 12303 5528 12348 5556
rect 12342 5516 12348 5528
rect 12400 5556 12406 5568
rect 12897 5559 12955 5565
rect 12897 5556 12909 5559
rect 12400 5528 12909 5556
rect 12400 5516 12406 5528
rect 12897 5525 12909 5528
rect 12943 5525 12955 5559
rect 12897 5519 12955 5525
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 14461 5559 14519 5565
rect 14461 5556 14473 5559
rect 13872 5528 14473 5556
rect 13872 5516 13878 5528
rect 14461 5525 14473 5528
rect 14507 5525 14519 5559
rect 20070 5556 20076 5568
rect 20031 5528 20076 5556
rect 14461 5519 14519 5525
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1854 5352 1860 5364
rect 1815 5324 1860 5352
rect 1854 5312 1860 5324
rect 1912 5312 1918 5364
rect 4062 5352 4068 5364
rect 4023 5324 4068 5352
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4522 5312 4528 5364
rect 4580 5352 4586 5364
rect 5721 5355 5779 5361
rect 5721 5352 5733 5355
rect 4580 5324 5733 5352
rect 4580 5312 4586 5324
rect 5721 5321 5733 5324
rect 5767 5321 5779 5355
rect 7006 5352 7012 5364
rect 6967 5324 7012 5352
rect 5721 5315 5779 5321
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7282 5312 7288 5364
rect 7340 5352 7346 5364
rect 7929 5355 7987 5361
rect 7929 5352 7941 5355
rect 7340 5324 7941 5352
rect 7340 5312 7346 5324
rect 2501 5287 2559 5293
rect 2501 5253 2513 5287
rect 2547 5284 2559 5287
rect 2590 5284 2596 5296
rect 2547 5256 2596 5284
rect 2547 5253 2559 5256
rect 2501 5247 2559 5253
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 3513 5287 3571 5293
rect 3513 5253 3525 5287
rect 3559 5284 3571 5287
rect 4614 5284 4620 5296
rect 3559 5256 4620 5284
rect 3559 5253 3571 5256
rect 3513 5247 3571 5253
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 5074 5244 5080 5296
rect 5132 5284 5138 5296
rect 6549 5287 6607 5293
rect 6549 5284 6561 5287
rect 5132 5256 6561 5284
rect 5132 5244 5138 5256
rect 6549 5253 6561 5256
rect 6595 5253 6607 5287
rect 6549 5247 6607 5253
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 2869 5219 2927 5225
rect 2869 5216 2881 5219
rect 2832 5188 2881 5216
rect 2832 5176 2838 5188
rect 2869 5185 2881 5188
rect 2915 5185 2927 5219
rect 2869 5179 2927 5185
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5216 3111 5219
rect 4062 5216 4068 5228
rect 3099 5188 4068 5216
rect 3099 5185 3111 5188
rect 3053 5179 3111 5185
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5148 2375 5151
rect 3068 5148 3096 5179
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5216 4583 5219
rect 5442 5216 5448 5228
rect 4571 5188 5448 5216
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 2363 5120 3096 5148
rect 2363 5117 2375 5120
rect 2317 5111 2375 5117
rect 3602 5108 3608 5160
rect 3660 5148 3666 5160
rect 4540 5148 4568 5179
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 6564 5216 6592 5247
rect 7576 5225 7604 5324
rect 7929 5321 7941 5324
rect 7975 5321 7987 5355
rect 8478 5352 8484 5364
rect 8439 5324 8484 5352
rect 7929 5315 7987 5321
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 9916 5324 10057 5352
rect 9916 5312 9922 5324
rect 10045 5321 10057 5324
rect 10091 5321 10103 5355
rect 10962 5352 10968 5364
rect 10923 5324 10968 5352
rect 10045 5315 10103 5321
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 12989 5355 13047 5361
rect 12989 5352 13001 5355
rect 12492 5324 13001 5352
rect 12492 5312 12498 5324
rect 12989 5321 13001 5324
rect 13035 5321 13047 5355
rect 12989 5315 13047 5321
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 6564 5188 7389 5216
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5185 7619 5219
rect 8496 5216 8524 5312
rect 8665 5219 8723 5225
rect 8665 5216 8677 5219
rect 8496 5188 8677 5216
rect 7561 5179 7619 5185
rect 8665 5185 8677 5188
rect 8711 5185 8723 5219
rect 13004 5216 13032 5315
rect 14458 5312 14464 5364
rect 14516 5352 14522 5364
rect 15378 5352 15384 5364
rect 14516 5324 15384 5352
rect 14516 5312 14522 5324
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 15930 5352 15936 5364
rect 15891 5324 15936 5352
rect 15930 5312 15936 5324
rect 15988 5312 15994 5364
rect 16301 5355 16359 5361
rect 16301 5321 16313 5355
rect 16347 5352 16359 5355
rect 16390 5352 16396 5364
rect 16347 5324 16396 5352
rect 16347 5321 16359 5324
rect 16301 5315 16359 5321
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 18874 5312 18880 5364
rect 18932 5352 18938 5364
rect 19061 5355 19119 5361
rect 19061 5352 19073 5355
rect 18932 5324 19073 5352
rect 18932 5312 18938 5324
rect 19061 5321 19073 5324
rect 19107 5321 19119 5355
rect 19426 5352 19432 5364
rect 19387 5324 19432 5352
rect 19061 5315 19119 5321
rect 19426 5312 19432 5324
rect 19484 5352 19490 5364
rect 19978 5352 19984 5364
rect 19484 5324 19984 5352
rect 19484 5312 19490 5324
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 20990 5352 20996 5364
rect 20951 5324 20996 5352
rect 20990 5312 20996 5324
rect 21048 5312 21054 5364
rect 16482 5284 16488 5296
rect 16443 5256 16488 5284
rect 16482 5244 16488 5256
rect 16540 5244 16546 5296
rect 18141 5287 18199 5293
rect 18141 5253 18153 5287
rect 18187 5253 18199 5287
rect 18141 5247 18199 5253
rect 13354 5216 13360 5228
rect 13004 5188 13360 5216
rect 8665 5179 8723 5185
rect 13354 5176 13360 5188
rect 13412 5216 13418 5228
rect 13541 5219 13599 5225
rect 13541 5216 13553 5219
rect 13412 5188 13553 5216
rect 13412 5176 13418 5188
rect 13541 5185 13553 5188
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5216 17003 5219
rect 17218 5216 17224 5228
rect 16991 5188 17224 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 17218 5176 17224 5188
rect 17276 5216 17282 5228
rect 18156 5216 18184 5247
rect 17276 5188 18184 5216
rect 18601 5219 18659 5225
rect 17276 5176 17282 5188
rect 18601 5185 18613 5219
rect 18647 5216 18659 5219
rect 18892 5216 18920 5312
rect 19518 5244 19524 5296
rect 19576 5284 19582 5296
rect 19705 5287 19763 5293
rect 19705 5284 19717 5287
rect 19576 5256 19717 5284
rect 19576 5244 19582 5256
rect 19705 5253 19717 5256
rect 19751 5253 19763 5287
rect 19705 5247 19763 5253
rect 18647 5188 18920 5216
rect 18647 5185 18659 5188
rect 18601 5179 18659 5185
rect 20070 5176 20076 5228
rect 20128 5216 20134 5228
rect 20257 5219 20315 5225
rect 20257 5216 20269 5219
rect 20128 5188 20269 5216
rect 20128 5176 20134 5188
rect 20257 5185 20269 5188
rect 20303 5185 20315 5219
rect 20257 5179 20315 5185
rect 3660 5120 4568 5148
rect 4617 5151 4675 5157
rect 3660 5108 3666 5120
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 4706 5148 4712 5160
rect 4663 5120 4712 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5148 5595 5151
rect 6086 5148 6092 5160
rect 5583 5120 6092 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 6086 5108 6092 5120
rect 6144 5108 6150 5160
rect 6273 5151 6331 5157
rect 6273 5117 6285 5151
rect 6319 5148 6331 5151
rect 11146 5148 11152 5160
rect 6319 5120 7512 5148
rect 11107 5120 11152 5148
rect 6319 5117 6331 5120
rect 6273 5111 6331 5117
rect 3326 5080 3332 5092
rect 3239 5052 3332 5080
rect 3326 5040 3332 5052
rect 3384 5080 3390 5092
rect 3786 5080 3792 5092
rect 3384 5052 3792 5080
rect 3384 5040 3390 5052
rect 3786 5040 3792 5052
rect 3844 5040 3850 5092
rect 4154 5040 4160 5092
rect 4212 5080 4218 5092
rect 4525 5083 4583 5089
rect 4525 5080 4537 5083
rect 4212 5052 4537 5080
rect 4212 5040 4218 5052
rect 4525 5049 4537 5052
rect 4571 5080 4583 5083
rect 4985 5083 5043 5089
rect 4985 5080 4997 5083
rect 4571 5052 4997 5080
rect 4571 5049 4583 5052
rect 4525 5043 4583 5049
rect 4985 5049 4997 5052
rect 5031 5080 5043 5083
rect 6730 5080 6736 5092
rect 5031 5052 6736 5080
rect 5031 5049 5043 5052
rect 4985 5043 5043 5049
rect 6730 5040 6736 5052
rect 6788 5040 6794 5092
rect 7484 5089 7512 5120
rect 11146 5108 11152 5120
rect 11204 5148 11210 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11204 5120 12081 5148
rect 11204 5108 11210 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 13808 5151 13866 5157
rect 12492 5120 12537 5148
rect 12492 5108 12498 5120
rect 13808 5117 13820 5151
rect 13854 5148 13866 5151
rect 14090 5148 14096 5160
rect 13854 5120 14096 5148
rect 13854 5117 13866 5120
rect 13808 5111 13866 5117
rect 14090 5108 14096 5120
rect 14148 5108 14154 5160
rect 15565 5151 15623 5157
rect 15565 5117 15577 5151
rect 15611 5148 15623 5151
rect 17037 5151 17095 5157
rect 17037 5148 17049 5151
rect 15611 5120 17049 5148
rect 15611 5117 15623 5120
rect 15565 5111 15623 5117
rect 17037 5117 17049 5120
rect 17083 5148 17095 5151
rect 17402 5148 17408 5160
rect 17083 5120 17408 5148
rect 17083 5117 17095 5120
rect 17037 5111 17095 5117
rect 17402 5108 17408 5120
rect 17460 5108 17466 5160
rect 17954 5108 17960 5160
rect 18012 5148 18018 5160
rect 18506 5148 18512 5160
rect 18012 5120 18512 5148
rect 18012 5108 18018 5120
rect 18506 5108 18512 5120
rect 18564 5148 18570 5160
rect 18693 5151 18751 5157
rect 18693 5148 18705 5151
rect 18564 5120 18705 5148
rect 18564 5108 18570 5120
rect 18693 5117 18705 5120
rect 18739 5148 18751 5151
rect 20088 5148 20116 5176
rect 20714 5148 20720 5160
rect 18739 5120 20116 5148
rect 20675 5120 20720 5148
rect 18739 5117 18751 5120
rect 18693 5111 18751 5117
rect 20714 5108 20720 5120
rect 20772 5108 20778 5160
rect 7469 5083 7527 5089
rect 7469 5049 7481 5083
rect 7515 5080 7527 5083
rect 7650 5080 7656 5092
rect 7515 5052 7656 5080
rect 7515 5049 7527 5052
rect 7469 5043 7527 5049
rect 7650 5040 7656 5052
rect 7708 5040 7714 5092
rect 8754 5040 8760 5092
rect 8812 5080 8818 5092
rect 8910 5083 8968 5089
rect 8910 5080 8922 5083
rect 8812 5052 8922 5080
rect 8812 5040 8818 5052
rect 8910 5049 8922 5052
rect 8956 5080 8968 5083
rect 9582 5080 9588 5092
rect 8956 5052 9588 5080
rect 8956 5049 8968 5052
rect 8910 5043 8968 5049
rect 9582 5040 9588 5052
rect 9640 5040 9646 5092
rect 12710 5040 12716 5092
rect 12768 5080 12774 5092
rect 13357 5083 13415 5089
rect 13357 5080 13369 5083
rect 12768 5052 13369 5080
rect 12768 5040 12774 5052
rect 13357 5049 13369 5052
rect 13403 5049 13415 5083
rect 13357 5043 13415 5049
rect 2961 5015 3019 5021
rect 2961 4981 2973 5015
rect 3007 5012 3019 5015
rect 3344 5012 3372 5040
rect 3007 4984 3372 5012
rect 3881 5015 3939 5021
rect 3007 4981 3019 4984
rect 2961 4975 3019 4981
rect 3881 4981 3893 5015
rect 3927 5012 3939 5015
rect 4430 5012 4436 5024
rect 3927 4984 4436 5012
rect 3927 4981 3939 4984
rect 3881 4975 3939 4981
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 5442 5012 5448 5024
rect 5403 4984 5448 5012
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 6086 4972 6092 5024
rect 6144 5012 6150 5024
rect 8662 5012 8668 5024
rect 6144 4984 8668 5012
rect 6144 4972 6150 4984
rect 8662 4972 8668 4984
rect 8720 5012 8726 5024
rect 9122 5012 9128 5024
rect 8720 4984 9128 5012
rect 8720 4972 8726 4984
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 10686 5012 10692 5024
rect 10647 4984 10692 5012
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 11330 5012 11336 5024
rect 11291 4984 11336 5012
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 11422 4972 11428 5024
rect 11480 5012 11486 5024
rect 11698 5012 11704 5024
rect 11480 4984 11704 5012
rect 11480 4972 11486 4984
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 12618 5012 12624 5024
rect 12579 4984 12624 5012
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 13372 5012 13400 5043
rect 14274 5040 14280 5092
rect 14332 5080 14338 5092
rect 17773 5083 17831 5089
rect 17773 5080 17785 5083
rect 14332 5052 17785 5080
rect 14332 5040 14338 5052
rect 17773 5049 17785 5052
rect 17819 5080 17831 5083
rect 18598 5080 18604 5092
rect 17819 5052 18604 5080
rect 17819 5049 17831 5052
rect 17773 5043 17831 5049
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 19610 5040 19616 5092
rect 19668 5040 19674 5092
rect 19978 5080 19984 5092
rect 19939 5052 19984 5080
rect 19978 5040 19984 5052
rect 20036 5040 20042 5092
rect 13906 5012 13912 5024
rect 13372 4984 13912 5012
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 14826 4972 14832 5024
rect 14884 5012 14890 5024
rect 14921 5015 14979 5021
rect 14921 5012 14933 5015
rect 14884 4984 14933 5012
rect 14884 4972 14890 4984
rect 14921 4981 14933 4984
rect 14967 4981 14979 5015
rect 16942 5012 16948 5024
rect 16903 4984 16948 5012
rect 14921 4975 14979 4981
rect 16942 4972 16948 4984
rect 17000 4972 17006 5024
rect 17218 4972 17224 5024
rect 17276 5012 17282 5024
rect 17405 5015 17463 5021
rect 17405 5012 17417 5015
rect 17276 4984 17417 5012
rect 17276 4972 17282 4984
rect 17405 4981 17417 4984
rect 17451 5012 17463 5015
rect 17586 5012 17592 5024
rect 17451 4984 17592 5012
rect 17451 4981 17463 4984
rect 17405 4975 17463 4981
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 19628 5012 19656 5040
rect 20165 5015 20223 5021
rect 20165 5012 20177 5015
rect 19628 4984 20177 5012
rect 20165 4981 20177 4984
rect 20211 5012 20223 5015
rect 20438 5012 20444 5024
rect 20211 4984 20444 5012
rect 20211 4981 20223 4984
rect 20165 4975 20223 4981
rect 20438 4972 20444 4984
rect 20496 4972 20502 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 4614 4808 4620 4820
rect 4575 4780 4620 4808
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 5905 4811 5963 4817
rect 5905 4808 5917 4811
rect 5592 4780 5917 4808
rect 5592 4768 5598 4780
rect 5905 4777 5917 4780
rect 5951 4777 5963 4811
rect 5905 4771 5963 4777
rect 2958 4740 2964 4752
rect 2919 4712 2964 4740
rect 2958 4700 2964 4712
rect 3016 4700 3022 4752
rect 3881 4743 3939 4749
rect 3881 4709 3893 4743
rect 3927 4740 3939 4743
rect 4706 4740 4712 4752
rect 3927 4712 4712 4740
rect 3927 4709 3939 4712
rect 3881 4703 3939 4709
rect 3896 4616 3924 4703
rect 4706 4700 4712 4712
rect 4764 4700 4770 4752
rect 4062 4632 4068 4684
rect 4120 4672 4126 4684
rect 4433 4675 4491 4681
rect 4433 4672 4445 4675
rect 4120 4644 4445 4672
rect 4120 4632 4126 4644
rect 4433 4641 4445 4644
rect 4479 4641 4491 4675
rect 5920 4672 5948 4771
rect 6178 4768 6184 4820
rect 6236 4808 6242 4820
rect 6273 4811 6331 4817
rect 6273 4808 6285 4811
rect 6236 4780 6285 4808
rect 6236 4768 6242 4780
rect 6273 4777 6285 4780
rect 6319 4777 6331 4811
rect 8754 4808 8760 4820
rect 8715 4780 8760 4808
rect 6273 4771 6331 4777
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 10134 4768 10140 4820
rect 10192 4808 10198 4820
rect 10229 4811 10287 4817
rect 10229 4808 10241 4811
rect 10192 4780 10241 4808
rect 10192 4768 10198 4780
rect 10229 4777 10241 4780
rect 10275 4777 10287 4811
rect 10229 4771 10287 4777
rect 12069 4811 12127 4817
rect 12069 4777 12081 4811
rect 12115 4808 12127 4811
rect 12158 4808 12164 4820
rect 12115 4780 12164 4808
rect 12115 4777 12127 4780
rect 12069 4771 12127 4777
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 14090 4808 14096 4820
rect 14051 4780 14096 4808
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 15562 4768 15568 4820
rect 15620 4808 15626 4820
rect 16117 4811 16175 4817
rect 16117 4808 16129 4811
rect 15620 4780 16129 4808
rect 15620 4768 15626 4780
rect 16117 4777 16129 4780
rect 16163 4777 16175 4811
rect 16117 4771 16175 4777
rect 16942 4768 16948 4820
rect 17000 4808 17006 4820
rect 19061 4811 19119 4817
rect 19061 4808 19073 4811
rect 17000 4780 19073 4808
rect 17000 4768 17006 4780
rect 19061 4777 19073 4780
rect 19107 4808 19119 4811
rect 19518 4808 19524 4820
rect 19107 4780 19524 4808
rect 19107 4777 19119 4780
rect 19061 4771 19119 4777
rect 19518 4768 19524 4780
rect 19576 4768 19582 4820
rect 6822 4749 6828 4752
rect 6816 4740 6828 4749
rect 6783 4712 6828 4740
rect 6816 4703 6828 4712
rect 6822 4700 6828 4703
rect 6880 4700 6886 4752
rect 12989 4743 13047 4749
rect 12989 4709 13001 4743
rect 13035 4740 13047 4743
rect 13538 4740 13544 4752
rect 13035 4712 13544 4740
rect 13035 4709 13047 4712
rect 12989 4703 13047 4709
rect 13538 4700 13544 4712
rect 13596 4740 13602 4752
rect 13725 4743 13783 4749
rect 13725 4740 13737 4743
rect 13596 4712 13737 4740
rect 13596 4700 13602 4712
rect 13725 4709 13737 4712
rect 13771 4709 13783 4743
rect 13725 4703 13783 4709
rect 6546 4672 6552 4684
rect 5920 4644 6552 4672
rect 4433 4635 4491 4641
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 9950 4632 9956 4684
rect 10008 4672 10014 4684
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 10008 4644 10057 4672
rect 10008 4632 10014 4644
rect 10045 4641 10057 4644
rect 10091 4641 10103 4675
rect 10045 4635 10103 4641
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 12161 4675 12219 4681
rect 12161 4672 12173 4675
rect 11471 4644 12173 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 12161 4641 12173 4644
rect 12207 4672 12219 4675
rect 12342 4672 12348 4684
rect 12207 4644 12348 4672
rect 12207 4641 12219 4644
rect 12161 4635 12219 4641
rect 12342 4632 12348 4644
rect 12400 4632 12406 4684
rect 13262 4632 13268 4684
rect 13320 4672 13326 4684
rect 13449 4675 13507 4681
rect 13449 4672 13461 4675
rect 13320 4644 13461 4672
rect 13320 4632 13326 4644
rect 13449 4641 13461 4644
rect 13495 4641 13507 4675
rect 13449 4635 13507 4641
rect 15105 4675 15163 4681
rect 15105 4641 15117 4675
rect 15151 4672 15163 4675
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 15151 4644 16221 4672
rect 15151 4641 15163 4644
rect 15105 4635 15163 4641
rect 16209 4641 16221 4644
rect 16255 4672 16267 4675
rect 16577 4675 16635 4681
rect 16577 4672 16589 4675
rect 16255 4644 16589 4672
rect 16255 4641 16267 4644
rect 16209 4635 16267 4641
rect 16577 4641 16589 4644
rect 16623 4672 16635 4675
rect 16666 4672 16672 4684
rect 16623 4644 16672 4672
rect 16623 4641 16635 4644
rect 16577 4635 16635 4641
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 17218 4632 17224 4684
rect 17276 4632 17282 4684
rect 17402 4681 17408 4684
rect 17396 4672 17408 4681
rect 17363 4644 17408 4672
rect 17396 4635 17408 4644
rect 17402 4632 17408 4635
rect 17460 4632 17466 4684
rect 19610 4672 19616 4684
rect 19571 4644 19616 4672
rect 19610 4632 19616 4644
rect 19668 4632 19674 4684
rect 20898 4672 20904 4684
rect 20859 4644 20904 4672
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 2225 4607 2283 4613
rect 2225 4604 2237 4607
rect 1443 4576 2237 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 2225 4573 2237 4576
rect 2271 4604 2283 4607
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2271 4576 2881 4604
rect 2271 4573 2283 4576
rect 2225 4567 2283 4573
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4573 3111 4607
rect 3053 4567 3111 4573
rect 2498 4536 2504 4548
rect 2459 4508 2504 4536
rect 2498 4496 2504 4508
rect 2556 4496 2562 4548
rect 1762 4428 1768 4480
rect 1820 4468 1826 4480
rect 1857 4471 1915 4477
rect 1857 4468 1869 4471
rect 1820 4440 1869 4468
rect 1820 4428 1826 4440
rect 1857 4437 1869 4440
rect 1903 4468 1915 4471
rect 2866 4468 2872 4480
rect 1903 4440 2872 4468
rect 1903 4437 1915 4440
rect 1857 4431 1915 4437
rect 2866 4428 2872 4440
rect 2924 4468 2930 4480
rect 3068 4468 3096 4567
rect 3878 4564 3884 4616
rect 3936 4564 3942 4616
rect 9858 4564 9864 4616
rect 9916 4604 9922 4616
rect 10321 4607 10379 4613
rect 10321 4604 10333 4607
rect 9916 4576 10333 4604
rect 9916 4564 9922 4576
rect 10321 4573 10333 4576
rect 10367 4573 10379 4607
rect 12066 4604 12072 4616
rect 12027 4576 12072 4604
rect 10321 4567 10379 4573
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 12529 4607 12587 4613
rect 12529 4604 12541 4607
rect 12360 4576 12541 4604
rect 12360 4548 12388 4576
rect 12529 4573 12541 4576
rect 12575 4573 12587 4607
rect 12529 4567 12587 4573
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4573 16175 4607
rect 16117 4567 16175 4573
rect 17129 4607 17187 4613
rect 17129 4573 17141 4607
rect 17175 4604 17187 4607
rect 17236 4604 17264 4632
rect 17175 4576 17264 4604
rect 20257 4607 20315 4613
rect 17175 4573 17187 4576
rect 17129 4567 17187 4573
rect 20257 4573 20269 4607
rect 20303 4604 20315 4607
rect 20530 4604 20536 4616
rect 20303 4576 20536 4604
rect 20303 4573 20315 4576
rect 20257 4567 20315 4573
rect 4157 4539 4215 4545
rect 4157 4505 4169 4539
rect 4203 4536 4215 4539
rect 4798 4536 4804 4548
rect 4203 4508 4804 4536
rect 4203 4505 4215 4508
rect 4157 4499 4215 4505
rect 4798 4496 4804 4508
rect 4856 4496 4862 4548
rect 9766 4536 9772 4548
rect 9727 4508 9772 4536
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 12342 4496 12348 4548
rect 12400 4496 12406 4548
rect 13998 4536 14004 4548
rect 12452 4508 14004 4536
rect 3510 4468 3516 4480
rect 2924 4440 3516 4468
rect 2924 4428 2930 4440
rect 3510 4428 3516 4440
rect 3568 4428 3574 4480
rect 4338 4428 4344 4480
rect 4396 4468 4402 4480
rect 5077 4471 5135 4477
rect 5077 4468 5089 4471
rect 4396 4440 5089 4468
rect 4396 4428 4402 4440
rect 5077 4437 5089 4440
rect 5123 4468 5135 4471
rect 5445 4471 5503 4477
rect 5445 4468 5457 4471
rect 5123 4440 5457 4468
rect 5123 4437 5135 4440
rect 5077 4431 5135 4437
rect 5445 4437 5457 4440
rect 5491 4437 5503 4471
rect 5445 4431 5503 4437
rect 6730 4428 6736 4480
rect 6788 4468 6794 4480
rect 7929 4471 7987 4477
rect 7929 4468 7941 4471
rect 6788 4440 7941 4468
rect 6788 4428 6794 4440
rect 7929 4437 7941 4440
rect 7975 4437 7987 4471
rect 7929 4431 7987 4437
rect 8938 4428 8944 4480
rect 8996 4468 9002 4480
rect 9125 4471 9183 4477
rect 9125 4468 9137 4471
rect 8996 4440 9137 4468
rect 8996 4428 9002 4440
rect 9125 4437 9137 4440
rect 9171 4468 9183 4471
rect 9401 4471 9459 4477
rect 9401 4468 9413 4471
rect 9171 4440 9413 4468
rect 9171 4437 9183 4440
rect 9125 4431 9183 4437
rect 9401 4437 9413 4440
rect 9447 4437 9459 4471
rect 9401 4431 9459 4437
rect 10781 4471 10839 4477
rect 10781 4437 10793 4471
rect 10827 4468 10839 4471
rect 10962 4468 10968 4480
rect 10827 4440 10968 4468
rect 10827 4437 10839 4440
rect 10781 4431 10839 4437
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 11609 4471 11667 4477
rect 11609 4437 11621 4471
rect 11655 4468 11667 4471
rect 12452 4468 12480 4508
rect 13998 4496 14004 4508
rect 14056 4536 14062 4548
rect 14461 4539 14519 4545
rect 14461 4536 14473 4539
rect 14056 4508 14473 4536
rect 14056 4496 14062 4508
rect 14461 4505 14473 4508
rect 14507 4505 14519 4539
rect 16132 4536 16160 4567
rect 16206 4536 16212 4548
rect 16132 4508 16212 4536
rect 14461 4499 14519 4505
rect 16206 4496 16212 4508
rect 16264 4496 16270 4548
rect 16574 4496 16580 4548
rect 16632 4536 16638 4548
rect 17144 4536 17172 4567
rect 20530 4564 20536 4576
rect 20588 4564 20594 4616
rect 18506 4536 18512 4548
rect 16632 4508 17172 4536
rect 18467 4508 18512 4536
rect 16632 4496 16638 4508
rect 18506 4496 18512 4508
rect 18564 4496 18570 4548
rect 19797 4539 19855 4545
rect 19797 4505 19809 4539
rect 19843 4536 19855 4539
rect 20714 4536 20720 4548
rect 19843 4508 20720 4536
rect 19843 4505 19855 4508
rect 19797 4499 19855 4505
rect 20714 4496 20720 4508
rect 20772 4496 20778 4548
rect 11655 4440 12480 4468
rect 13173 4471 13231 4477
rect 11655 4437 11667 4440
rect 11609 4431 11667 4437
rect 13173 4437 13185 4471
rect 13219 4468 13231 4471
rect 13722 4468 13728 4480
rect 13219 4440 13728 4468
rect 13219 4437 13231 4440
rect 13173 4431 13231 4437
rect 13722 4428 13728 4440
rect 13780 4428 13786 4480
rect 15654 4468 15660 4480
rect 15615 4440 15660 4468
rect 15654 4428 15660 4440
rect 15712 4428 15718 4480
rect 16850 4428 16856 4480
rect 16908 4468 16914 4480
rect 16945 4471 17003 4477
rect 16945 4468 16957 4471
rect 16908 4440 16957 4468
rect 16908 4428 16914 4440
rect 16945 4437 16957 4440
rect 16991 4437 17003 4471
rect 19426 4468 19432 4480
rect 19387 4440 19432 4468
rect 16945 4431 17003 4437
rect 19426 4428 19432 4440
rect 19484 4428 19490 4480
rect 19886 4428 19892 4480
rect 19944 4468 19950 4480
rect 20533 4471 20591 4477
rect 20533 4468 20545 4471
rect 19944 4440 20545 4468
rect 19944 4428 19950 4440
rect 20533 4437 20545 4440
rect 20579 4437 20591 4471
rect 21082 4468 21088 4480
rect 21043 4440 21088 4468
rect 20533 4431 20591 4437
rect 21082 4428 21088 4440
rect 21140 4428 21146 4480
rect 21450 4468 21456 4480
rect 21411 4440 21456 4468
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 2958 4224 2964 4276
rect 3016 4264 3022 4276
rect 3145 4267 3203 4273
rect 3145 4264 3157 4267
rect 3016 4236 3157 4264
rect 3016 4224 3022 4236
rect 3145 4233 3157 4236
rect 3191 4264 3203 4267
rect 4614 4264 4620 4276
rect 3191 4236 4620 4264
rect 3191 4233 3203 4236
rect 3145 4227 3203 4233
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 6273 4267 6331 4273
rect 6273 4233 6285 4267
rect 6319 4264 6331 4267
rect 6822 4264 6828 4276
rect 6319 4236 6828 4264
rect 6319 4233 6331 4236
rect 6273 4227 6331 4233
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 10134 4264 10140 4276
rect 10095 4236 10140 4264
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 11701 4267 11759 4273
rect 11701 4233 11713 4267
rect 11747 4264 11759 4267
rect 12066 4264 12072 4276
rect 11747 4236 12072 4264
rect 11747 4233 11759 4236
rect 11701 4227 11759 4233
rect 12066 4224 12072 4236
rect 12124 4224 12130 4276
rect 13265 4267 13323 4273
rect 13265 4233 13277 4267
rect 13311 4264 13323 4267
rect 13630 4264 13636 4276
rect 13311 4236 13636 4264
rect 13311 4233 13323 4236
rect 13265 4227 13323 4233
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 14458 4264 14464 4276
rect 13832 4236 14464 4264
rect 6546 4196 6552 4208
rect 6507 4168 6552 4196
rect 6546 4156 6552 4168
rect 6604 4196 6610 4208
rect 7282 4196 7288 4208
rect 6604 4168 7288 4196
rect 6604 4156 6610 4168
rect 7282 4156 7288 4168
rect 7340 4196 7346 4208
rect 7929 4199 7987 4205
rect 7929 4196 7941 4199
rect 7340 4168 7941 4196
rect 7340 4156 7346 4168
rect 7929 4165 7941 4168
rect 7975 4196 7987 4199
rect 10686 4196 10692 4208
rect 7975 4168 8156 4196
rect 10647 4168 10692 4196
rect 7975 4165 7987 4168
rect 7929 4159 7987 4165
rect 2130 4088 2136 4140
rect 2188 4088 2194 4140
rect 2222 4088 2228 4140
rect 2280 4128 2286 4140
rect 3513 4131 3571 4137
rect 3513 4128 3525 4131
rect 2280 4100 3525 4128
rect 2280 4088 2286 4100
rect 3513 4097 3525 4100
rect 3559 4128 3571 4131
rect 4062 4128 4068 4140
rect 3559 4100 4068 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5718 4128 5724 4140
rect 5123 4100 5724 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 7374 4128 7380 4140
rect 5859 4100 7380 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 7374 4088 7380 4100
rect 7432 4128 7438 4140
rect 8128 4137 8156 4168
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 11974 4156 11980 4208
rect 12032 4196 12038 4208
rect 13832 4196 13860 4236
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 15562 4224 15568 4276
rect 15620 4264 15626 4276
rect 15749 4267 15807 4273
rect 15749 4264 15761 4267
rect 15620 4236 15761 4264
rect 15620 4224 15626 4236
rect 15749 4233 15761 4236
rect 15795 4233 15807 4267
rect 15749 4227 15807 4233
rect 16574 4224 16580 4276
rect 16632 4264 16638 4276
rect 17313 4267 17371 4273
rect 17313 4264 17325 4267
rect 16632 4236 17325 4264
rect 16632 4224 16638 4236
rect 17313 4233 17325 4236
rect 17359 4233 17371 4267
rect 17313 4227 17371 4233
rect 19518 4224 19524 4276
rect 19576 4264 19582 4276
rect 20254 4264 20260 4276
rect 19576 4236 20260 4264
rect 19576 4224 19582 4236
rect 20254 4224 20260 4236
rect 20312 4224 20318 4276
rect 20898 4224 20904 4276
rect 20956 4264 20962 4276
rect 21085 4267 21143 4273
rect 21085 4264 21097 4267
rect 20956 4236 21097 4264
rect 20956 4224 20962 4236
rect 21085 4233 21097 4236
rect 21131 4233 21143 4267
rect 21085 4227 21143 4233
rect 12032 4168 13860 4196
rect 12032 4156 12038 4168
rect 15654 4156 15660 4208
rect 15712 4196 15718 4208
rect 19610 4196 19616 4208
rect 15712 4168 16528 4196
rect 19571 4168 19616 4196
rect 15712 4156 15718 4168
rect 7561 4131 7619 4137
rect 7561 4128 7573 4131
rect 7432 4100 7573 4128
rect 7432 4088 7438 4100
rect 7561 4097 7573 4100
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 12069 4131 12127 4137
rect 12069 4097 12081 4131
rect 12115 4128 12127 4131
rect 12158 4128 12164 4140
rect 12115 4100 12164 4128
rect 12115 4097 12127 4100
rect 12069 4091 12127 4097
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 13354 4088 13360 4140
rect 13412 4128 13418 4140
rect 13633 4131 13691 4137
rect 13633 4128 13645 4131
rect 13412 4100 13645 4128
rect 13412 4088 13418 4100
rect 13633 4097 13645 4100
rect 13679 4128 13691 4131
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13679 4100 13829 4128
rect 13679 4097 13691 4100
rect 13633 4091 13691 4097
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 16500 4128 16528 4168
rect 19610 4156 19616 4168
rect 19668 4156 19674 4208
rect 16761 4131 16819 4137
rect 16761 4128 16773 4131
rect 16500 4100 16773 4128
rect 13817 4091 13875 4097
rect 16761 4097 16773 4100
rect 16807 4128 16819 4131
rect 18785 4131 18843 4137
rect 18785 4128 18797 4131
rect 16807 4100 18797 4128
rect 16807 4097 16819 4100
rect 16761 4091 16819 4097
rect 18785 4097 18797 4100
rect 18831 4097 18843 4131
rect 18785 4091 18843 4097
rect 2148 4060 2176 4088
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 2148 4032 2421 4060
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 2866 4060 2872 4072
rect 2731 4032 2872 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 3970 4060 3976 4072
rect 3931 4032 3976 4060
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 5243 4063 5301 4069
rect 5243 4029 5255 4063
rect 5289 4060 5301 4063
rect 6454 4060 6460 4072
rect 5289 4032 6460 4060
rect 5289 4029 5301 4032
rect 5243 4023 5301 4029
rect 6454 4020 6460 4032
rect 6512 4020 6518 4072
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 2115 3995 2173 4001
rect 2115 3961 2127 3995
rect 2161 3992 2173 3995
rect 2222 3992 2228 4004
rect 2161 3964 2228 3992
rect 2161 3961 2173 3964
rect 2115 3955 2173 3961
rect 2222 3952 2228 3964
rect 2280 3952 2286 4004
rect 2774 3952 2780 4004
rect 2832 3992 2838 4004
rect 4249 3995 4307 4001
rect 4249 3992 4261 3995
rect 2832 3964 4261 3992
rect 2832 3952 2838 3964
rect 4249 3961 4261 3964
rect 4295 3992 4307 3995
rect 4338 3992 4344 4004
rect 4295 3964 4344 3992
rect 4295 3961 4307 3964
rect 4249 3955 4307 3961
rect 4338 3952 4344 3964
rect 4396 3952 4402 4004
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 6270 3992 6276 4004
rect 5592 3964 6276 3992
rect 5592 3952 5598 3964
rect 6270 3952 6276 3964
rect 6328 3992 6334 4004
rect 6840 3992 6868 4023
rect 9858 4020 9864 4072
rect 9916 4060 9922 4072
rect 11241 4063 11299 4069
rect 11241 4060 11253 4063
rect 9916 4032 11253 4060
rect 9916 4020 9922 4032
rect 11241 4029 11253 4032
rect 11287 4029 11299 4063
rect 11241 4023 11299 4029
rect 11882 4020 11888 4072
rect 11940 4060 11946 4072
rect 12342 4060 12348 4072
rect 11940 4032 12348 4060
rect 11940 4020 11946 4032
rect 12342 4020 12348 4032
rect 12400 4060 12406 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12400 4032 12449 4060
rect 12400 4020 12406 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 16375 4063 16433 4069
rect 16375 4029 16387 4063
rect 16421 4060 16433 4063
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 16421 4032 18061 4060
rect 16421 4029 16433 4032
rect 16375 4023 16433 4029
rect 18049 4029 18061 4032
rect 18095 4060 18107 4063
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 18095 4032 19165 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 20162 4060 20168 4072
rect 20123 4032 20168 4060
rect 19153 4023 19211 4029
rect 20162 4020 20168 4032
rect 20220 4060 20226 4072
rect 20717 4063 20775 4069
rect 20717 4060 20729 4063
rect 20220 4032 20729 4060
rect 20220 4020 20226 4032
rect 20717 4029 20729 4032
rect 20763 4029 20775 4063
rect 21266 4060 21272 4072
rect 21227 4032 21272 4060
rect 20717 4023 20775 4029
rect 21266 4020 21272 4032
rect 21324 4060 21330 4072
rect 21821 4063 21879 4069
rect 21821 4060 21833 4063
rect 21324 4032 21833 4060
rect 21324 4020 21330 4032
rect 21821 4029 21833 4032
rect 21867 4029 21879 4063
rect 21821 4023 21879 4029
rect 7098 3992 7104 4004
rect 6328 3964 6868 3992
rect 7059 3964 7104 3992
rect 6328 3952 6334 3964
rect 7098 3952 7104 3964
rect 7156 3952 7162 4004
rect 8380 3995 8438 4001
rect 8380 3961 8392 3995
rect 8426 3992 8438 3995
rect 8938 3992 8944 4004
rect 8426 3964 8944 3992
rect 8426 3961 8438 3964
rect 8380 3955 8438 3961
rect 8938 3952 8944 3964
rect 8996 3952 9002 4004
rect 10965 3995 11023 4001
rect 10965 3961 10977 3995
rect 11011 3961 11023 3995
rect 12250 3992 12256 4004
rect 10965 3955 11023 3961
rect 11348 3964 12256 3992
rect 1949 3927 2007 3933
rect 1949 3893 1961 3927
rect 1995 3924 2007 3927
rect 2590 3924 2596 3936
rect 1995 3896 2596 3924
rect 1995 3893 2007 3896
rect 1949 3887 2007 3893
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 3687 3927 3745 3933
rect 3687 3893 3699 3927
rect 3733 3924 3745 3927
rect 4062 3924 4068 3936
rect 3733 3896 4068 3924
rect 3733 3893 3745 3896
rect 3687 3887 3745 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4154 3884 4160 3936
rect 4212 3924 4218 3936
rect 4212 3896 4257 3924
rect 4212 3884 4218 3896
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 5721 3927 5779 3933
rect 5721 3924 5733 3927
rect 5684 3896 5733 3924
rect 5684 3884 5690 3896
rect 5721 3893 5733 3896
rect 5767 3893 5779 3927
rect 5721 3887 5779 3893
rect 8202 3884 8208 3936
rect 8260 3924 8266 3936
rect 9490 3924 9496 3936
rect 8260 3896 9496 3924
rect 8260 3884 8266 3896
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10413 3927 10471 3933
rect 10413 3924 10425 3927
rect 10192 3896 10425 3924
rect 10192 3884 10198 3896
rect 10413 3893 10425 3896
rect 10459 3924 10471 3927
rect 10980 3924 11008 3955
rect 10459 3896 11008 3924
rect 10459 3893 10471 3896
rect 10413 3887 10471 3893
rect 11054 3884 11060 3936
rect 11112 3924 11118 3936
rect 11149 3927 11207 3933
rect 11149 3924 11161 3927
rect 11112 3896 11161 3924
rect 11112 3884 11118 3896
rect 11149 3893 11161 3896
rect 11195 3924 11207 3927
rect 11348 3924 11376 3964
rect 12250 3952 12256 3964
rect 12308 3952 12314 4004
rect 12710 3992 12716 4004
rect 12671 3964 12716 3992
rect 12710 3952 12716 3964
rect 12768 3952 12774 4004
rect 13538 3952 13544 4004
rect 13596 3992 13602 4004
rect 14084 3995 14142 4001
rect 14084 3992 14096 3995
rect 13596 3964 14096 3992
rect 13596 3952 13602 3964
rect 14084 3961 14096 3964
rect 14130 3992 14142 3995
rect 14366 3992 14372 4004
rect 14130 3964 14372 3992
rect 14130 3961 14142 3964
rect 14084 3955 14142 3961
rect 14366 3952 14372 3964
rect 14424 3952 14430 4004
rect 16942 3992 16948 4004
rect 16903 3964 16948 3992
rect 16942 3952 16948 3964
rect 17000 3992 17006 4004
rect 17402 3992 17408 4004
rect 17000 3964 17408 3992
rect 17000 3952 17006 3964
rect 17402 3952 17408 3964
rect 17460 3992 17466 4004
rect 17681 3995 17739 4001
rect 17681 3992 17693 3995
rect 17460 3964 17693 3992
rect 17460 3952 17466 3964
rect 17681 3961 17693 3964
rect 17727 3961 17739 3995
rect 18322 3992 18328 4004
rect 18283 3964 18328 3992
rect 17681 3955 17739 3961
rect 18322 3952 18328 3964
rect 18380 3952 18386 4004
rect 19426 3952 19432 4004
rect 19484 3992 19490 4004
rect 19981 3995 20039 4001
rect 19981 3992 19993 3995
rect 19484 3964 19993 3992
rect 19484 3952 19490 3964
rect 19981 3961 19993 3964
rect 20027 3961 20039 3995
rect 19981 3955 20039 3961
rect 20070 3952 20076 4004
rect 20128 3992 20134 4004
rect 20128 3964 21496 3992
rect 20128 3952 20134 3964
rect 11195 3896 11376 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 13170 3884 13176 3936
rect 13228 3924 13234 3936
rect 13630 3924 13636 3936
rect 13228 3896 13636 3924
rect 13228 3884 13234 3896
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 14458 3884 14464 3936
rect 14516 3924 14522 3936
rect 15197 3927 15255 3933
rect 15197 3924 15209 3927
rect 14516 3896 15209 3924
rect 14516 3884 14522 3896
rect 15197 3893 15209 3896
rect 15243 3893 15255 3927
rect 16206 3924 16212 3936
rect 16167 3896 16212 3924
rect 15197 3887 15255 3893
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 16850 3924 16856 3936
rect 16811 3896 16856 3924
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 20346 3924 20352 3936
rect 20307 3896 20352 3924
rect 20346 3884 20352 3896
rect 20404 3884 20410 3936
rect 21468 3933 21496 3964
rect 21453 3927 21511 3933
rect 21453 3893 21465 3927
rect 21499 3893 21511 3927
rect 22370 3924 22376 3936
rect 22331 3896 22376 3924
rect 21453 3887 21511 3893
rect 22370 3884 22376 3896
rect 22428 3884 22434 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 2130 3720 2136 3732
rect 2091 3692 2136 3720
rect 2130 3680 2136 3692
rect 2188 3680 2194 3732
rect 2961 3723 3019 3729
rect 2961 3689 2973 3723
rect 3007 3720 3019 3723
rect 3234 3720 3240 3732
rect 3007 3692 3240 3720
rect 3007 3689 3019 3692
rect 2961 3683 3019 3689
rect 3234 3680 3240 3692
rect 3292 3680 3298 3732
rect 3878 3720 3884 3732
rect 3839 3692 3884 3720
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 5994 3720 6000 3732
rect 5592 3692 6000 3720
rect 5592 3680 5598 3692
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 6454 3720 6460 3732
rect 6415 3692 6460 3720
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 8478 3720 8484 3732
rect 6564 3692 8484 3720
rect 2590 3612 2596 3664
rect 2648 3652 2654 3664
rect 2777 3655 2835 3661
rect 2777 3652 2789 3655
rect 2648 3624 2789 3652
rect 2648 3612 2654 3624
rect 2777 3621 2789 3624
rect 2823 3652 2835 3655
rect 3602 3652 3608 3664
rect 2823 3624 3608 3652
rect 2823 3621 2835 3624
rect 2777 3615 2835 3621
rect 3602 3612 3608 3624
rect 3660 3612 3666 3664
rect 4062 3612 4068 3664
rect 4120 3652 4126 3664
rect 4433 3655 4491 3661
rect 4433 3652 4445 3655
rect 4120 3624 4445 3652
rect 4120 3612 4126 3624
rect 4433 3621 4445 3624
rect 4479 3621 4491 3655
rect 4614 3652 4620 3664
rect 4575 3624 4620 3652
rect 4433 3615 4491 3621
rect 4614 3612 4620 3624
rect 4672 3612 4678 3664
rect 6086 3612 6092 3664
rect 6144 3652 6150 3664
rect 6564 3661 6592 3692
rect 6273 3655 6331 3661
rect 6273 3652 6285 3655
rect 6144 3624 6285 3652
rect 6144 3612 6150 3624
rect 6273 3621 6285 3624
rect 6319 3621 6331 3655
rect 6273 3615 6331 3621
rect 6549 3655 6607 3661
rect 6549 3621 6561 3655
rect 6595 3621 6607 3655
rect 6549 3615 6607 3621
rect 7193 3655 7251 3661
rect 7193 3621 7205 3655
rect 7239 3652 7251 3655
rect 7282 3652 7288 3664
rect 7239 3624 7288 3652
rect 7239 3621 7251 3624
rect 7193 3615 7251 3621
rect 7282 3612 7288 3624
rect 7340 3612 7346 3664
rect 8128 3661 8156 3692
rect 8478 3680 8484 3692
rect 8536 3720 8542 3732
rect 8938 3720 8944 3732
rect 8536 3692 8944 3720
rect 8536 3680 8542 3692
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10229 3723 10287 3729
rect 10229 3720 10241 3723
rect 10008 3692 10241 3720
rect 10008 3680 10014 3692
rect 10229 3689 10241 3692
rect 10275 3720 10287 3723
rect 10778 3720 10784 3732
rect 10275 3692 10784 3720
rect 10275 3689 10287 3692
rect 10229 3683 10287 3689
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 12161 3723 12219 3729
rect 12161 3689 12173 3723
rect 12207 3720 12219 3723
rect 12618 3720 12624 3732
rect 12207 3692 12624 3720
rect 12207 3689 12219 3692
rect 12161 3683 12219 3689
rect 8021 3655 8079 3661
rect 8021 3621 8033 3655
rect 8067 3621 8079 3655
rect 8021 3615 8079 3621
rect 8113 3655 8171 3661
rect 8113 3621 8125 3655
rect 8159 3621 8171 3655
rect 8113 3615 8171 3621
rect 9493 3655 9551 3661
rect 9493 3621 9505 3655
rect 9539 3652 9551 3655
rect 9858 3652 9864 3664
rect 9539 3624 9864 3652
rect 9539 3621 9551 3624
rect 9493 3615 9551 3621
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 3053 3587 3111 3593
rect 3053 3553 3065 3587
rect 3099 3584 3111 3587
rect 3510 3584 3516 3596
rect 3099 3556 3516 3584
rect 3099 3553 3111 3556
rect 3053 3547 3111 3553
rect 3510 3544 3516 3556
rect 3568 3584 3574 3596
rect 3970 3584 3976 3596
rect 3568 3556 3976 3584
rect 3568 3544 3574 3556
rect 3970 3544 3976 3556
rect 4028 3584 4034 3596
rect 5629 3587 5687 3593
rect 5629 3584 5641 3587
rect 4028 3556 5641 3584
rect 4028 3544 4034 3556
rect 5629 3553 5641 3556
rect 5675 3584 5687 3587
rect 6730 3584 6736 3596
rect 5675 3556 6736 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 7834 3584 7840 3596
rect 7795 3556 7840 3584
rect 7834 3544 7840 3556
rect 7892 3544 7898 3596
rect 4706 3516 4712 3528
rect 4667 3488 4712 3516
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 7466 3516 7472 3528
rect 6604 3488 7472 3516
rect 6604 3476 6610 3488
rect 7466 3476 7472 3488
rect 7524 3516 7530 3528
rect 8036 3516 8064 3615
rect 9858 3612 9864 3624
rect 9916 3652 9922 3664
rect 10597 3655 10655 3661
rect 10597 3652 10609 3655
rect 9916 3624 10609 3652
rect 9916 3612 9922 3624
rect 10597 3621 10609 3624
rect 10643 3652 10655 3655
rect 12176 3652 12204 3683
rect 12618 3680 12624 3692
rect 12676 3720 12682 3732
rect 12713 3723 12771 3729
rect 12713 3720 12725 3723
rect 12676 3692 12725 3720
rect 12676 3680 12682 3692
rect 12713 3689 12725 3692
rect 12759 3689 12771 3723
rect 13814 3720 13820 3732
rect 13775 3692 13820 3720
rect 12713 3683 12771 3689
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 14826 3680 14832 3732
rect 14884 3720 14890 3732
rect 14921 3723 14979 3729
rect 14921 3720 14933 3723
rect 14884 3692 14933 3720
rect 14884 3680 14890 3692
rect 14921 3689 14933 3692
rect 14967 3689 14979 3723
rect 14921 3683 14979 3689
rect 16393 3723 16451 3729
rect 16393 3689 16405 3723
rect 16439 3720 16451 3723
rect 16942 3720 16948 3732
rect 16439 3692 16948 3720
rect 16439 3689 16451 3692
rect 16393 3683 16451 3689
rect 16942 3680 16948 3692
rect 17000 3720 17006 3732
rect 17957 3723 18015 3729
rect 17957 3720 17969 3723
rect 17000 3692 17969 3720
rect 17000 3680 17006 3692
rect 17957 3689 17969 3692
rect 18003 3689 18015 3723
rect 17957 3683 18015 3689
rect 21358 3680 21364 3732
rect 21416 3720 21422 3732
rect 21453 3723 21511 3729
rect 21453 3720 21465 3723
rect 21416 3692 21465 3720
rect 21416 3680 21422 3692
rect 21453 3689 21465 3692
rect 21499 3689 21511 3723
rect 21453 3683 21511 3689
rect 10643 3624 12204 3652
rect 13173 3655 13231 3661
rect 10643 3621 10655 3624
rect 10597 3615 10655 3621
rect 13173 3621 13185 3655
rect 13219 3652 13231 3655
rect 13262 3652 13268 3664
rect 13219 3624 13268 3652
rect 13219 3621 13231 3624
rect 13173 3615 13231 3621
rect 13262 3612 13268 3624
rect 13320 3612 13326 3664
rect 13633 3655 13691 3661
rect 13633 3621 13645 3655
rect 13679 3652 13691 3655
rect 13722 3652 13728 3664
rect 13679 3624 13728 3652
rect 13679 3621 13691 3624
rect 13633 3615 13691 3621
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 15565 3655 15623 3661
rect 15565 3621 15577 3655
rect 15611 3652 15623 3655
rect 16022 3652 16028 3664
rect 15611 3624 16028 3652
rect 15611 3621 15623 3624
rect 15565 3615 15623 3621
rect 16022 3612 16028 3624
rect 16080 3612 16086 3664
rect 16482 3652 16488 3664
rect 16224 3624 16488 3652
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 10781 3587 10839 3593
rect 10781 3553 10793 3587
rect 10827 3584 10839 3587
rect 10870 3584 10876 3596
rect 10827 3556 10876 3584
rect 10827 3553 10839 3556
rect 10781 3547 10839 3553
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 11054 3593 11060 3596
rect 11048 3584 11060 3593
rect 11015 3556 11060 3584
rect 11048 3547 11060 3556
rect 11054 3544 11060 3547
rect 11112 3544 11118 3596
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3584 15347 3587
rect 16224 3584 16252 3624
rect 16482 3612 16488 3624
rect 16540 3652 16546 3664
rect 18877 3655 18935 3661
rect 18877 3652 18889 3655
rect 16540 3624 18889 3652
rect 16540 3612 16546 3624
rect 18877 3621 18889 3624
rect 18923 3621 18935 3655
rect 18877 3615 18935 3621
rect 15335 3556 16252 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 16666 3544 16672 3596
rect 16724 3584 16730 3596
rect 16833 3587 16891 3593
rect 16833 3584 16845 3587
rect 16724 3556 16845 3584
rect 16724 3544 16730 3556
rect 16833 3553 16845 3556
rect 16879 3584 16891 3587
rect 18509 3587 18567 3593
rect 18509 3584 18521 3587
rect 16879 3556 18521 3584
rect 16879 3553 16891 3556
rect 16833 3547 16891 3553
rect 18509 3553 18521 3556
rect 18555 3584 18567 3587
rect 18690 3584 18696 3596
rect 18555 3556 18696 3584
rect 18555 3553 18567 3556
rect 18509 3547 18567 3553
rect 18690 3544 18696 3556
rect 18748 3544 18754 3596
rect 19058 3584 19064 3596
rect 19019 3556 19064 3584
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 20898 3584 20904 3596
rect 20859 3556 20904 3584
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 22002 3584 22008 3596
rect 21963 3556 22008 3584
rect 22002 3544 22008 3556
rect 22060 3544 22066 3596
rect 7524 3488 8064 3516
rect 13909 3519 13967 3525
rect 7524 3476 7530 3488
rect 13909 3485 13921 3519
rect 13955 3516 13967 3519
rect 14458 3516 14464 3528
rect 13955 3488 14464 3516
rect 13955 3485 13967 3488
rect 13909 3479 13967 3485
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 16574 3516 16580 3528
rect 16535 3488 16580 3516
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 19610 3516 19616 3528
rect 19571 3488 19616 3516
rect 19610 3476 19616 3488
rect 19668 3476 19674 3528
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 3878 3448 3884 3460
rect 3752 3420 3884 3448
rect 3752 3408 3758 3420
rect 3878 3408 3884 3420
rect 3936 3408 3942 3460
rect 4157 3451 4215 3457
rect 4157 3417 4169 3451
rect 4203 3448 4215 3451
rect 4246 3448 4252 3460
rect 4203 3420 4252 3448
rect 4203 3417 4215 3420
rect 4157 3411 4215 3417
rect 4246 3408 4252 3420
rect 4304 3408 4310 3460
rect 5261 3451 5319 3457
rect 5261 3417 5273 3451
rect 5307 3448 5319 3451
rect 5626 3448 5632 3460
rect 5307 3420 5632 3448
rect 5307 3417 5319 3420
rect 5261 3411 5319 3417
rect 5626 3408 5632 3420
rect 5684 3448 5690 3460
rect 6178 3448 6184 3460
rect 5684 3420 6184 3448
rect 5684 3408 5690 3420
rect 6178 3408 6184 3420
rect 6236 3408 6242 3460
rect 7374 3408 7380 3460
rect 7432 3448 7438 3460
rect 8294 3448 8300 3460
rect 7432 3420 8300 3448
rect 7432 3408 7438 3420
rect 8294 3408 8300 3420
rect 8352 3448 8358 3460
rect 8481 3451 8539 3457
rect 8481 3448 8493 3451
rect 8352 3420 8493 3448
rect 8352 3408 8358 3420
rect 8481 3417 8493 3420
rect 8527 3417 8539 3451
rect 13354 3448 13360 3460
rect 13315 3420 13360 3448
rect 8481 3411 8539 3417
rect 13354 3408 13360 3420
rect 13412 3408 13418 3460
rect 14366 3448 14372 3460
rect 14279 3420 14372 3448
rect 14366 3408 14372 3420
rect 14424 3448 14430 3460
rect 16482 3448 16488 3460
rect 14424 3420 16488 3448
rect 14424 3408 14430 3420
rect 16482 3408 16488 3420
rect 16540 3408 16546 3460
rect 21085 3451 21143 3457
rect 21085 3417 21097 3451
rect 21131 3448 21143 3451
rect 22738 3448 22744 3460
rect 21131 3420 22744 3448
rect 21131 3417 21143 3420
rect 21085 3411 21143 3417
rect 22738 3408 22744 3420
rect 22796 3408 22802 3460
rect 2498 3380 2504 3392
rect 2459 3352 2504 3380
rect 2498 3340 2504 3352
rect 2556 3340 2562 3392
rect 5997 3383 6055 3389
rect 5997 3349 6009 3383
rect 6043 3380 6055 3383
rect 6362 3380 6368 3392
rect 6043 3352 6368 3380
rect 6043 3349 6055 3352
rect 5997 3343 6055 3349
rect 6362 3340 6368 3352
rect 6420 3340 6426 3392
rect 7190 3340 7196 3392
rect 7248 3380 7254 3392
rect 7561 3383 7619 3389
rect 7561 3380 7573 3383
rect 7248 3352 7573 3380
rect 7248 3340 7254 3352
rect 7561 3349 7573 3352
rect 7607 3349 7619 3383
rect 7561 3343 7619 3349
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 9861 3383 9919 3389
rect 9861 3380 9873 3383
rect 9732 3352 9873 3380
rect 9732 3340 9738 3352
rect 9861 3349 9873 3352
rect 9907 3349 9919 3383
rect 19242 3380 19248 3392
rect 19203 3352 19248 3380
rect 9861 3343 9919 3349
rect 19242 3340 19248 3352
rect 19300 3340 19306 3392
rect 19978 3380 19984 3392
rect 19939 3352 19984 3380
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 20254 3340 20260 3392
rect 20312 3380 20318 3392
rect 20349 3383 20407 3389
rect 20349 3380 20361 3383
rect 20312 3352 20361 3380
rect 20312 3340 20318 3352
rect 20349 3349 20361 3352
rect 20395 3349 20407 3383
rect 21818 3380 21824 3392
rect 21779 3352 21824 3380
rect 20349 3343 20407 3349
rect 21818 3340 21824 3352
rect 21876 3340 21882 3392
rect 22186 3380 22192 3392
rect 22147 3352 22192 3380
rect 22186 3340 22192 3352
rect 22244 3340 22250 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1762 3176 1768 3188
rect 1723 3148 1768 3176
rect 1762 3136 1768 3148
rect 1820 3136 1826 3188
rect 2133 3179 2191 3185
rect 2133 3145 2145 3179
rect 2179 3176 2191 3179
rect 2590 3176 2596 3188
rect 2179 3148 2596 3176
rect 2179 3145 2191 3148
rect 2133 3139 2191 3145
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 3234 3176 3240 3188
rect 3195 3148 3240 3176
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 5997 3179 6055 3185
rect 5997 3145 6009 3179
rect 6043 3176 6055 3179
rect 6086 3176 6092 3188
rect 6043 3148 6092 3176
rect 6043 3145 6055 3148
rect 5997 3139 6055 3145
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 7282 3176 7288 3188
rect 7116 3148 7288 3176
rect 2314 3108 2320 3120
rect 2275 3080 2320 3108
rect 2314 3068 2320 3080
rect 2372 3068 2378 3120
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 7116 3049 7144 3148
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 8478 3176 8484 3188
rect 8439 3148 8484 3176
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 10870 3136 10876 3188
rect 10928 3176 10934 3188
rect 11517 3179 11575 3185
rect 11517 3176 11529 3179
rect 10928 3148 11529 3176
rect 10928 3136 10934 3148
rect 11517 3145 11529 3148
rect 11563 3176 11575 3179
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 11563 3148 12173 3176
rect 11563 3145 11575 3148
rect 11517 3139 11575 3145
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 14458 3176 14464 3188
rect 14419 3148 14464 3176
rect 12161 3139 12219 3145
rect 2869 3043 2927 3049
rect 2869 3040 2881 3043
rect 2832 3012 2881 3040
rect 2832 3000 2838 3012
rect 2869 3009 2881 3012
rect 2915 3009 2927 3043
rect 2869 3003 2927 3009
rect 7101 3043 7159 3049
rect 7101 3009 7113 3043
rect 7147 3009 7159 3043
rect 12176 3040 12204 3139
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 18141 3179 18199 3185
rect 18141 3176 18153 3179
rect 16908 3148 18153 3176
rect 16908 3136 16914 3148
rect 18141 3145 18153 3148
rect 18187 3145 18199 3179
rect 19058 3176 19064 3188
rect 19019 3148 19064 3176
rect 18141 3139 18199 3145
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 19429 3179 19487 3185
rect 19429 3176 19441 3179
rect 19392 3148 19441 3176
rect 19392 3136 19398 3148
rect 19429 3145 19441 3148
rect 19475 3145 19487 3179
rect 19429 3139 19487 3145
rect 17126 3068 17132 3120
rect 17184 3108 17190 3120
rect 17405 3111 17463 3117
rect 17405 3108 17417 3111
rect 17184 3080 17417 3108
rect 17184 3068 17190 3080
rect 17405 3077 17417 3080
rect 17451 3077 17463 3111
rect 17405 3071 17463 3077
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 12176 3012 12449 3040
rect 7101 3003 7159 3009
rect 12437 3009 12449 3012
rect 12483 3009 12495 3043
rect 12437 3003 12495 3009
rect 2222 2932 2228 2984
rect 2280 2972 2286 2984
rect 2590 2972 2596 2984
rect 2280 2944 2596 2972
rect 2280 2932 2286 2944
rect 2590 2932 2596 2944
rect 2648 2932 2654 2984
rect 3789 2975 3847 2981
rect 3789 2972 3801 2975
rect 3712 2944 3801 2972
rect 3712 2848 3740 2944
rect 3789 2941 3801 2944
rect 3835 2941 3847 2975
rect 6546 2972 6552 2984
rect 6507 2944 6552 2972
rect 3789 2935 3847 2941
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 7374 2981 7380 2984
rect 7368 2972 7380 2981
rect 7335 2944 7380 2972
rect 7368 2935 7380 2944
rect 7374 2932 7380 2935
rect 7432 2932 7438 2984
rect 7834 2932 7840 2984
rect 7892 2972 7898 2984
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 7892 2944 9045 2972
rect 7892 2932 7898 2944
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 9493 2975 9551 2981
rect 9493 2941 9505 2975
rect 9539 2972 9551 2975
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 9539 2944 9597 2972
rect 9539 2941 9551 2944
rect 9493 2935 9551 2941
rect 9585 2941 9597 2944
rect 9631 2972 9643 2975
rect 10870 2972 10876 2984
rect 9631 2944 10876 2972
rect 9631 2941 9643 2944
rect 9585 2935 9643 2941
rect 10870 2932 10876 2944
rect 10928 2932 10934 2984
rect 12452 2972 12480 3003
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 12452 2944 14749 2972
rect 14737 2941 14749 2944
rect 14783 2972 14795 2975
rect 14918 2972 14924 2984
rect 14783 2944 14924 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 14918 2932 14924 2944
rect 14976 2972 14982 2984
rect 16574 2972 16580 2984
rect 14976 2944 16580 2972
rect 14976 2932 14982 2944
rect 16574 2932 16580 2944
rect 16632 2972 16638 2984
rect 16853 2975 16911 2981
rect 16853 2972 16865 2975
rect 16632 2944 16865 2972
rect 16632 2932 16638 2944
rect 16853 2941 16865 2944
rect 16899 2941 16911 2975
rect 16853 2935 16911 2941
rect 3970 2864 3976 2916
rect 4028 2913 4034 2916
rect 4028 2907 4092 2913
rect 4028 2873 4046 2907
rect 4080 2873 4092 2907
rect 9830 2907 9888 2913
rect 9830 2904 9842 2907
rect 4028 2867 4092 2873
rect 9508 2876 9842 2904
rect 4028 2864 4034 2867
rect 9508 2848 9536 2876
rect 9830 2873 9842 2876
rect 9876 2873 9888 2907
rect 9830 2867 9888 2873
rect 9950 2864 9956 2916
rect 10008 2904 10014 2916
rect 12066 2904 12072 2916
rect 10008 2876 12072 2904
rect 10008 2864 10014 2876
rect 12066 2864 12072 2876
rect 12124 2864 12130 2916
rect 12618 2864 12624 2916
rect 12676 2913 12682 2916
rect 12676 2907 12740 2913
rect 12676 2873 12694 2907
rect 12728 2873 12740 2907
rect 12676 2867 12740 2873
rect 12676 2864 12682 2867
rect 14826 2864 14832 2916
rect 14884 2904 14890 2916
rect 15166 2907 15224 2913
rect 15166 2904 15178 2907
rect 14884 2876 15178 2904
rect 14884 2864 14890 2876
rect 15166 2873 15178 2876
rect 15212 2873 15224 2907
rect 17420 2904 17448 3071
rect 17865 3043 17923 3049
rect 17865 3009 17877 3043
rect 17911 3040 17923 3043
rect 18138 3040 18144 3052
rect 17911 3012 18144 3040
rect 17911 3009 17923 3012
rect 17865 3003 17923 3009
rect 18138 3000 18144 3012
rect 18196 3040 18202 3052
rect 18509 3043 18567 3049
rect 18509 3040 18521 3043
rect 18196 3012 18521 3040
rect 18196 3000 18202 3012
rect 18509 3009 18521 3012
rect 18555 3009 18567 3043
rect 18690 3040 18696 3052
rect 18651 3012 18696 3040
rect 18509 3003 18567 3009
rect 18690 3000 18696 3012
rect 18748 3000 18754 3052
rect 19444 3040 19472 3139
rect 19610 3136 19616 3188
rect 19668 3176 19674 3188
rect 22002 3176 22008 3188
rect 19668 3148 20300 3176
rect 21963 3148 22008 3176
rect 19668 3136 19674 3148
rect 20272 3049 20300 3148
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 22649 3111 22707 3117
rect 22649 3077 22661 3111
rect 22695 3108 22707 3111
rect 23842 3108 23848 3120
rect 22695 3080 23848 3108
rect 22695 3077 22707 3080
rect 22649 3071 22707 3077
rect 23842 3068 23848 3080
rect 23900 3068 23906 3120
rect 20073 3043 20131 3049
rect 20073 3040 20085 3043
rect 19444 3012 20085 3040
rect 20073 3009 20085 3012
rect 20119 3009 20131 3043
rect 20073 3003 20131 3009
rect 20257 3043 20315 3049
rect 20257 3009 20269 3043
rect 20303 3009 20315 3043
rect 23658 3040 23664 3052
rect 23619 3012 23664 3040
rect 20257 3003 20315 3009
rect 23658 3000 23664 3012
rect 23716 3000 23722 3052
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 19687 2975 19745 2981
rect 19687 2972 19699 2975
rect 19392 2944 19699 2972
rect 19392 2932 19398 2944
rect 19687 2941 19699 2944
rect 19733 2972 19745 2975
rect 20622 2972 20628 2984
rect 19733 2944 20628 2972
rect 19733 2941 19745 2944
rect 19687 2935 19745 2941
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 21177 2975 21235 2981
rect 21177 2941 21189 2975
rect 21223 2972 21235 2975
rect 21358 2972 21364 2984
rect 21223 2944 21364 2972
rect 21223 2941 21235 2944
rect 21177 2935 21235 2941
rect 21358 2932 21364 2944
rect 21416 2932 21422 2984
rect 21453 2975 21511 2981
rect 21453 2941 21465 2975
rect 21499 2972 21511 2975
rect 22465 2975 22523 2981
rect 22465 2972 22477 2975
rect 21499 2944 22477 2972
rect 21499 2941 21511 2944
rect 21453 2935 21511 2941
rect 22465 2941 22477 2944
rect 22511 2972 22523 2975
rect 23017 2975 23075 2981
rect 23017 2972 23029 2975
rect 22511 2944 23029 2972
rect 22511 2941 22523 2944
rect 22465 2935 22523 2941
rect 23017 2941 23029 2944
rect 23063 2941 23075 2975
rect 23017 2935 23075 2941
rect 18601 2907 18659 2913
rect 18601 2904 18613 2907
rect 17420 2876 18613 2904
rect 15166 2867 15224 2873
rect 18601 2873 18613 2876
rect 18647 2904 18659 2907
rect 20162 2904 20168 2916
rect 18647 2876 19656 2904
rect 20123 2876 20168 2904
rect 18647 2873 18659 2876
rect 18601 2867 18659 2873
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3694 2836 3700 2848
rect 2832 2808 2877 2836
rect 3655 2808 3700 2836
rect 2832 2796 2838 2808
rect 3694 2796 3700 2808
rect 3752 2796 3758 2848
rect 4338 2796 4344 2848
rect 4396 2836 4402 2848
rect 5169 2839 5227 2845
rect 5169 2836 5181 2839
rect 4396 2808 5181 2836
rect 4396 2796 4402 2808
rect 5169 2805 5181 2808
rect 5215 2805 5227 2839
rect 5169 2799 5227 2805
rect 9490 2796 9496 2848
rect 9548 2796 9554 2848
rect 10965 2839 11023 2845
rect 10965 2805 10977 2839
rect 11011 2836 11023 2839
rect 11146 2836 11152 2848
rect 11011 2808 11152 2836
rect 11011 2805 11023 2808
rect 10965 2799 11023 2805
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 11238 2796 11244 2848
rect 11296 2836 11302 2848
rect 11698 2836 11704 2848
rect 11296 2808 11704 2836
rect 11296 2796 11302 2808
rect 11698 2796 11704 2808
rect 11756 2836 11762 2848
rect 13817 2839 13875 2845
rect 13817 2836 13829 2839
rect 11756 2808 13829 2836
rect 11756 2796 11762 2808
rect 13817 2805 13829 2808
rect 13863 2805 13875 2839
rect 13817 2799 13875 2805
rect 16301 2839 16359 2845
rect 16301 2805 16313 2839
rect 16347 2836 16359 2839
rect 16482 2836 16488 2848
rect 16347 2808 16488 2836
rect 16347 2805 16359 2808
rect 16301 2799 16359 2805
rect 16482 2796 16488 2808
rect 16540 2796 16546 2848
rect 19628 2836 19656 2876
rect 20162 2864 20168 2876
rect 20220 2864 20226 2916
rect 20898 2836 20904 2848
rect 19628 2808 20904 2836
rect 20898 2796 20904 2808
rect 20956 2796 20962 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2961 2635 3019 2641
rect 2961 2632 2973 2635
rect 1995 2604 2973 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2961 2601 2973 2604
rect 3007 2632 3019 2635
rect 4890 2632 4896 2644
rect 3007 2604 4896 2632
rect 3007 2601 3019 2604
rect 2961 2595 3019 2601
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 6733 2635 6791 2641
rect 6733 2601 6745 2635
rect 6779 2632 6791 2635
rect 7282 2632 7288 2644
rect 6779 2604 7288 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 9490 2632 9496 2644
rect 9451 2604 9496 2632
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 10321 2635 10379 2641
rect 10321 2601 10333 2635
rect 10367 2632 10379 2635
rect 10686 2632 10692 2644
rect 10367 2604 10692 2632
rect 10367 2601 10379 2604
rect 10321 2595 10379 2601
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 10873 2635 10931 2641
rect 10873 2601 10885 2635
rect 10919 2632 10931 2635
rect 11146 2632 11152 2644
rect 10919 2604 11152 2632
rect 10919 2601 10931 2604
rect 10873 2595 10931 2601
rect 11146 2592 11152 2604
rect 11204 2632 11210 2644
rect 11204 2604 13308 2632
rect 11204 2592 11210 2604
rect 3053 2567 3111 2573
rect 3053 2533 3065 2567
rect 3099 2564 3111 2567
rect 3970 2564 3976 2576
rect 3099 2536 3976 2564
rect 3099 2533 3111 2536
rect 3053 2527 3111 2533
rect 3970 2524 3976 2536
rect 4028 2524 4034 2576
rect 4338 2573 4344 2576
rect 4332 2564 4344 2573
rect 4299 2536 4344 2564
rect 4332 2527 4344 2536
rect 4338 2524 4344 2527
rect 4396 2524 4402 2576
rect 6549 2567 6607 2573
rect 6549 2533 6561 2567
rect 6595 2564 6607 2567
rect 7162 2567 7220 2573
rect 7162 2564 7174 2567
rect 6595 2536 7174 2564
rect 6595 2533 6607 2536
rect 6549 2527 6607 2533
rect 7162 2533 7174 2536
rect 7208 2533 7220 2567
rect 7162 2527 7220 2533
rect 3694 2456 3700 2508
rect 3752 2496 3758 2508
rect 3881 2499 3939 2505
rect 3881 2496 3893 2499
rect 3752 2468 3893 2496
rect 3752 2456 3758 2468
rect 3881 2465 3893 2468
rect 3927 2496 3939 2499
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3927 2468 4077 2496
rect 3927 2465 3939 2468
rect 3881 2459 3939 2465
rect 4065 2465 4077 2468
rect 4111 2496 4123 2499
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 4111 2468 6929 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 6917 2465 6929 2468
rect 6963 2496 6975 2499
rect 7291 2496 7319 2592
rect 9766 2524 9772 2576
rect 9824 2564 9830 2576
rect 10137 2567 10195 2573
rect 10137 2564 10149 2567
rect 9824 2536 10149 2564
rect 9824 2524 9830 2536
rect 10137 2533 10149 2536
rect 10183 2533 10195 2567
rect 10137 2527 10195 2533
rect 10413 2567 10471 2573
rect 10413 2533 10425 2567
rect 10459 2564 10471 2567
rect 11238 2564 11244 2576
rect 10459 2536 11244 2564
rect 10459 2533 10471 2536
rect 10413 2527 10471 2533
rect 6963 2468 7319 2496
rect 9217 2499 9275 2505
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 9217 2465 9229 2499
rect 9263 2496 9275 2499
rect 10428 2496 10456 2527
rect 11238 2524 11244 2536
rect 11296 2524 11302 2576
rect 12434 2524 12440 2576
rect 12492 2564 12498 2576
rect 12710 2564 12716 2576
rect 12492 2536 12716 2564
rect 12492 2524 12498 2536
rect 12710 2524 12716 2536
rect 12768 2564 12774 2576
rect 12989 2567 13047 2573
rect 12989 2564 13001 2567
rect 12768 2536 13001 2564
rect 12768 2524 12774 2536
rect 12989 2533 13001 2536
rect 13035 2533 13047 2567
rect 13170 2564 13176 2576
rect 13131 2536 13176 2564
rect 12989 2527 13047 2533
rect 13170 2524 13176 2536
rect 13228 2524 13234 2576
rect 13280 2573 13308 2604
rect 14918 2592 14924 2644
rect 14976 2632 14982 2644
rect 15197 2635 15255 2641
rect 15197 2632 15209 2635
rect 14976 2604 15209 2632
rect 14976 2592 14982 2604
rect 15197 2601 15209 2604
rect 15243 2601 15255 2635
rect 15197 2595 15255 2601
rect 13265 2567 13323 2573
rect 13265 2533 13277 2567
rect 13311 2564 13323 2567
rect 13633 2567 13691 2573
rect 13633 2564 13645 2567
rect 13311 2536 13645 2564
rect 13311 2533 13323 2536
rect 13265 2527 13323 2533
rect 13633 2533 13645 2536
rect 13679 2533 13691 2567
rect 13633 2527 13691 2533
rect 11146 2496 11152 2508
rect 9263 2468 10456 2496
rect 11107 2468 11152 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 11146 2456 11152 2468
rect 11204 2496 11210 2508
rect 11333 2499 11391 2505
rect 11333 2496 11345 2499
rect 11204 2468 11345 2496
rect 11204 2456 11210 2468
rect 11333 2465 11345 2468
rect 11379 2465 11391 2499
rect 11333 2459 11391 2465
rect 12069 2499 12127 2505
rect 12069 2465 12081 2499
rect 12115 2496 12127 2499
rect 13188 2496 13216 2524
rect 12115 2468 13216 2496
rect 12115 2465 12127 2468
rect 12069 2459 12127 2465
rect 13446 2456 13452 2508
rect 13504 2496 13510 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 13504 2468 14197 2496
rect 13504 2456 13510 2468
rect 14185 2465 14197 2468
rect 14231 2496 14243 2499
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14231 2468 14749 2496
rect 14231 2465 14243 2468
rect 14185 2459 14243 2465
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 15212 2496 15240 2595
rect 16666 2592 16672 2644
rect 16724 2632 16730 2644
rect 16853 2635 16911 2641
rect 16853 2632 16865 2635
rect 16724 2604 16865 2632
rect 16724 2592 16730 2604
rect 16853 2601 16865 2604
rect 16899 2601 16911 2635
rect 16853 2595 16911 2601
rect 18877 2635 18935 2641
rect 18877 2601 18889 2635
rect 18923 2632 18935 2635
rect 19334 2632 19340 2644
rect 18923 2604 19340 2632
rect 18923 2601 18935 2604
rect 18877 2595 18935 2601
rect 19334 2592 19340 2604
rect 19392 2592 19398 2644
rect 19705 2635 19763 2641
rect 19705 2601 19717 2635
rect 19751 2632 19763 2635
rect 20162 2632 20168 2644
rect 19751 2604 20168 2632
rect 19751 2601 19763 2604
rect 19705 2595 19763 2601
rect 20162 2592 20168 2604
rect 20220 2592 20226 2644
rect 20622 2592 20628 2644
rect 20680 2632 20686 2644
rect 20809 2635 20867 2641
rect 20809 2632 20821 2635
rect 20680 2604 20821 2632
rect 20680 2592 20686 2604
rect 20809 2601 20821 2604
rect 20855 2601 20867 2635
rect 20809 2595 20867 2601
rect 21453 2635 21511 2641
rect 21453 2601 21465 2635
rect 21499 2632 21511 2635
rect 23290 2632 23296 2644
rect 21499 2604 23296 2632
rect 21499 2601 21511 2604
rect 21453 2595 21511 2601
rect 23290 2592 23296 2604
rect 23348 2592 23354 2644
rect 20533 2567 20591 2573
rect 20533 2564 20545 2567
rect 19904 2536 20545 2564
rect 19904 2508 19932 2536
rect 20533 2533 20545 2536
rect 20579 2533 20591 2567
rect 20533 2527 20591 2533
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15212 2468 15485 2496
rect 14737 2459 14795 2465
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15729 2499 15787 2505
rect 15729 2496 15741 2499
rect 15473 2459 15531 2465
rect 15580 2468 15741 2496
rect 1394 2428 1400 2440
rect 1355 2400 1400 2428
rect 1394 2388 1400 2400
rect 1452 2388 1458 2440
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 2961 2431 3019 2437
rect 2961 2428 2973 2431
rect 2363 2400 2973 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 2961 2397 2973 2400
rect 3007 2428 3019 2431
rect 3602 2428 3608 2440
rect 3007 2400 3608 2428
rect 3007 2397 3019 2400
rect 2961 2391 3019 2397
rect 3602 2388 3608 2400
rect 3660 2388 3666 2440
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2428 14151 2431
rect 14458 2428 14464 2440
rect 14139 2400 14464 2428
rect 14139 2397 14151 2400
rect 14093 2391 14151 2397
rect 14458 2388 14464 2400
rect 14516 2428 14522 2440
rect 15580 2428 15608 2468
rect 15729 2465 15741 2468
rect 15775 2465 15787 2499
rect 15729 2459 15787 2465
rect 16574 2456 16580 2508
rect 16632 2496 16638 2508
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 16632 2468 17693 2496
rect 16632 2456 16638 2468
rect 17681 2465 17693 2468
rect 17727 2496 17739 2499
rect 18969 2499 19027 2505
rect 18969 2496 18981 2499
rect 17727 2468 18981 2496
rect 17727 2465 17739 2468
rect 17681 2459 17739 2465
rect 18969 2465 18981 2468
rect 19015 2465 19027 2499
rect 19886 2496 19892 2508
rect 19799 2468 19892 2496
rect 18969 2459 19027 2465
rect 19886 2456 19892 2468
rect 19944 2456 19950 2508
rect 20438 2456 20444 2508
rect 20496 2496 20502 2508
rect 21269 2499 21327 2505
rect 21269 2496 21281 2499
rect 20496 2468 21281 2496
rect 20496 2456 20502 2468
rect 21269 2465 21281 2468
rect 21315 2496 21327 2499
rect 21821 2499 21879 2505
rect 21821 2496 21833 2499
rect 21315 2468 21833 2496
rect 21315 2465 21327 2468
rect 21269 2459 21327 2465
rect 21821 2465 21833 2468
rect 21867 2465 21879 2499
rect 22462 2496 22468 2508
rect 22423 2468 22468 2496
rect 21821 2459 21879 2465
rect 22462 2456 22468 2468
rect 22520 2496 22526 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22520 2468 23029 2496
rect 22520 2456 22526 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 24026 2496 24032 2508
rect 23987 2468 24032 2496
rect 23017 2459 23075 2465
rect 24026 2456 24032 2468
rect 24084 2496 24090 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 24084 2468 24593 2496
rect 24084 2456 24090 2468
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 24581 2459 24639 2465
rect 18785 2431 18843 2437
rect 18785 2428 18797 2431
rect 14516 2400 15608 2428
rect 18064 2400 18797 2428
rect 14516 2388 14522 2400
rect 5350 2320 5356 2372
rect 5408 2360 5414 2372
rect 5994 2360 6000 2372
rect 5408 2332 6000 2360
rect 5408 2320 5414 2332
rect 5994 2320 6000 2332
rect 6052 2320 6058 2372
rect 9861 2363 9919 2369
rect 9861 2329 9873 2363
rect 9907 2360 9919 2363
rect 11882 2360 11888 2372
rect 9907 2332 11888 2360
rect 9907 2329 9919 2332
rect 9861 2323 9919 2329
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 12250 2320 12256 2372
rect 12308 2360 12314 2372
rect 12713 2363 12771 2369
rect 12713 2360 12725 2363
rect 12308 2332 12725 2360
rect 12308 2320 12314 2332
rect 12713 2329 12725 2332
rect 12759 2329 12771 2363
rect 14366 2360 14372 2372
rect 14327 2332 14372 2360
rect 12713 2323 12771 2329
rect 14366 2320 14372 2332
rect 14424 2320 14430 2372
rect 18064 2304 18092 2400
rect 18785 2397 18797 2400
rect 18831 2397 18843 2431
rect 18785 2391 18843 2397
rect 18322 2320 18328 2372
rect 18380 2360 18386 2372
rect 18417 2363 18475 2369
rect 18417 2360 18429 2363
rect 18380 2332 18429 2360
rect 18380 2320 18386 2332
rect 18417 2329 18429 2332
rect 18463 2329 18475 2363
rect 18417 2323 18475 2329
rect 20073 2363 20131 2369
rect 20073 2329 20085 2363
rect 20119 2360 20131 2363
rect 20622 2360 20628 2372
rect 20119 2332 20628 2360
rect 20119 2329 20131 2332
rect 20073 2323 20131 2329
rect 20622 2320 20628 2332
rect 20680 2320 20686 2372
rect 22649 2363 22707 2369
rect 22649 2329 22661 2363
rect 22695 2360 22707 2363
rect 24118 2360 24124 2372
rect 22695 2332 24124 2360
rect 22695 2329 22707 2332
rect 22649 2323 22707 2329
rect 24118 2320 24124 2332
rect 24176 2320 24182 2372
rect 2498 2292 2504 2304
rect 2459 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2292 2562 2304
rect 2774 2292 2780 2304
rect 2556 2264 2780 2292
rect 2556 2252 2562 2264
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 4706 2292 4712 2304
rect 3559 2264 4712 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 4706 2252 4712 2264
rect 4764 2292 4770 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 4764 2264 5457 2292
rect 4764 2252 4770 2264
rect 5445 2261 5457 2264
rect 5491 2292 5503 2295
rect 6273 2295 6331 2301
rect 6273 2292 6285 2295
rect 5491 2264 6285 2292
rect 5491 2261 5503 2264
rect 5445 2255 5503 2261
rect 6273 2261 6285 2264
rect 6319 2292 6331 2295
rect 6549 2295 6607 2301
rect 6549 2292 6561 2295
rect 6319 2264 6561 2292
rect 6319 2261 6331 2264
rect 6273 2255 6331 2261
rect 6549 2261 6561 2264
rect 6595 2261 6607 2295
rect 11514 2292 11520 2304
rect 11475 2264 11520 2292
rect 6549 2255 6607 2261
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 18046 2292 18052 2304
rect 18007 2264 18052 2292
rect 18046 2252 18052 2264
rect 18104 2252 18110 2304
rect 22186 2292 22192 2304
rect 22147 2264 22192 2292
rect 22186 2252 22192 2264
rect 22244 2252 22250 2304
rect 24210 2292 24216 2304
rect 24171 2264 24216 2292
rect 24210 2252 24216 2264
rect 24268 2252 24274 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 12894 1844 12900 1896
rect 12952 1884 12958 1896
rect 14182 1884 14188 1896
rect 12952 1856 14188 1884
rect 12952 1844 12958 1856
rect 14182 1844 14188 1856
rect 14240 1844 14246 1896
rect 15470 552 15476 604
rect 15528 592 15534 604
rect 16850 592 16856 604
rect 15528 564 16856 592
rect 15528 552 15534 564
rect 16850 552 16856 564
rect 16908 552 16914 604
rect 20714 552 20720 604
rect 20772 592 20778 604
rect 21174 592 21180 604
rect 20772 564 21180 592
rect 20772 552 20778 564
rect 21174 552 21180 564
rect 21232 552 21238 604
<< via1 >>
rect 4068 26256 4120 26308
rect 12164 26256 12216 26308
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 2320 25440 2372 25492
rect 3424 25372 3476 25424
rect 5448 25440 5500 25492
rect 3516 25304 3568 25356
rect 5172 25372 5224 25424
rect 8576 25372 8628 25424
rect 11520 25372 11572 25424
rect 7012 25304 7064 25356
rect 11060 25304 11112 25356
rect 14004 25304 14056 25356
rect 8484 25236 8536 25288
rect 11888 25236 11940 25288
rect 5632 25168 5684 25220
rect 6460 25168 6512 25220
rect 7932 25168 7984 25220
rect 23480 25168 23532 25220
rect 24308 25168 24360 25220
rect 4436 25143 4488 25152
rect 4436 25109 4445 25143
rect 4445 25109 4479 25143
rect 4479 25109 4488 25143
rect 4436 25100 4488 25109
rect 7748 25100 7800 25152
rect 10784 25100 10836 25152
rect 10968 25100 11020 25152
rect 25964 25100 26016 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 2872 24896 2924 24948
rect 3608 24896 3660 24948
rect 5172 24896 5224 24948
rect 3516 24871 3568 24880
rect 3516 24837 3525 24871
rect 3525 24837 3559 24871
rect 3559 24837 3568 24871
rect 3516 24828 3568 24837
rect 4068 24828 4120 24880
rect 11980 24896 12032 24948
rect 8484 24828 8536 24880
rect 11888 24828 11940 24880
rect 1400 24760 1452 24812
rect 4436 24760 4488 24812
rect 6092 24760 6144 24812
rect 10876 24760 10928 24812
rect 3424 24692 3476 24744
rect 7656 24692 7708 24744
rect 4620 24667 4672 24676
rect 4620 24633 4629 24667
rect 4629 24633 4663 24667
rect 4663 24633 4672 24667
rect 4620 24624 4672 24633
rect 7932 24692 7984 24744
rect 4068 24599 4120 24608
rect 4068 24565 4101 24599
rect 4101 24565 4120 24599
rect 4068 24556 4120 24565
rect 4436 24556 4488 24608
rect 9864 24624 9916 24676
rect 7012 24599 7064 24608
rect 7012 24565 7021 24599
rect 7021 24565 7055 24599
rect 7055 24565 7064 24599
rect 7012 24556 7064 24565
rect 7380 24556 7432 24608
rect 8576 24556 8628 24608
rect 9956 24556 10008 24608
rect 10784 24556 10836 24608
rect 11060 24599 11112 24608
rect 11060 24565 11069 24599
rect 11069 24565 11103 24599
rect 11103 24565 11112 24599
rect 11060 24556 11112 24565
rect 11520 24599 11572 24608
rect 11520 24565 11529 24599
rect 11529 24565 11563 24599
rect 11563 24565 11572 24599
rect 11520 24556 11572 24565
rect 11888 24599 11940 24608
rect 11888 24565 11897 24599
rect 11897 24565 11931 24599
rect 11931 24565 11940 24599
rect 11888 24556 11940 24565
rect 12440 24556 12492 24608
rect 14004 24599 14056 24608
rect 14004 24565 14013 24599
rect 14013 24565 14047 24599
rect 14047 24565 14056 24599
rect 14004 24556 14056 24565
rect 15108 24556 15160 24608
rect 15568 24599 15620 24608
rect 15568 24565 15577 24599
rect 15577 24565 15611 24599
rect 15611 24565 15620 24599
rect 15568 24556 15620 24565
rect 16120 24556 16172 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 3056 24352 3108 24404
rect 3516 24352 3568 24404
rect 7932 24352 7984 24404
rect 8668 24352 8720 24404
rect 9864 24352 9916 24404
rect 16488 24352 16540 24404
rect 17500 24352 17552 24404
rect 17684 24395 17736 24404
rect 17684 24361 17693 24395
rect 17693 24361 17727 24395
rect 17727 24361 17736 24395
rect 17684 24352 17736 24361
rect 19984 24352 20036 24404
rect 1676 24284 1728 24336
rect 4896 24327 4948 24336
rect 4896 24293 4905 24327
rect 4905 24293 4939 24327
rect 4939 24293 4948 24327
rect 4896 24284 4948 24293
rect 6368 24284 6420 24336
rect 8116 24327 8168 24336
rect 8116 24293 8125 24327
rect 8125 24293 8159 24327
rect 8159 24293 8168 24327
rect 8116 24284 8168 24293
rect 2504 24216 2556 24268
rect 4620 24216 4672 24268
rect 8484 24284 8536 24336
rect 11152 24284 11204 24336
rect 15292 24259 15344 24268
rect 6276 24148 6328 24200
rect 4988 24080 5040 24132
rect 6092 24123 6144 24132
rect 6092 24089 6101 24123
rect 6101 24089 6135 24123
rect 6135 24089 6144 24123
rect 6092 24080 6144 24089
rect 6920 24080 6972 24132
rect 8300 24148 8352 24200
rect 10600 24148 10652 24200
rect 15292 24225 15301 24259
rect 15301 24225 15335 24259
rect 15335 24225 15344 24259
rect 15292 24216 15344 24225
rect 16396 24259 16448 24268
rect 16396 24225 16405 24259
rect 16405 24225 16439 24259
rect 16439 24225 16448 24259
rect 16396 24216 16448 24225
rect 17408 24216 17460 24268
rect 20168 24216 20220 24268
rect 14280 24148 14332 24200
rect 7656 24123 7708 24132
rect 7656 24089 7665 24123
rect 7665 24089 7699 24123
rect 7699 24089 7708 24123
rect 7656 24080 7708 24089
rect 4436 24055 4488 24064
rect 4436 24021 4445 24055
rect 4445 24021 4479 24055
rect 4479 24021 4488 24055
rect 4436 24012 4488 24021
rect 6000 24012 6052 24064
rect 12072 24012 12124 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1492 23851 1544 23860
rect 1492 23817 1501 23851
rect 1501 23817 1535 23851
rect 1535 23817 1544 23851
rect 1492 23808 1544 23817
rect 4620 23808 4672 23860
rect 6092 23808 6144 23860
rect 6276 23808 6328 23860
rect 8300 23851 8352 23860
rect 8300 23817 8309 23851
rect 8309 23817 8343 23851
rect 8343 23817 8352 23851
rect 8300 23808 8352 23817
rect 10600 23808 10652 23860
rect 15292 23851 15344 23860
rect 5908 23740 5960 23792
rect 6368 23740 6420 23792
rect 6920 23783 6972 23792
rect 6920 23749 6929 23783
rect 6929 23749 6963 23783
rect 6963 23749 6972 23783
rect 6920 23740 6972 23749
rect 2044 23715 2096 23724
rect 2044 23681 2053 23715
rect 2053 23681 2087 23715
rect 2087 23681 2096 23715
rect 2044 23672 2096 23681
rect 7104 23672 7156 23724
rect 10876 23715 10928 23724
rect 10876 23681 10885 23715
rect 10885 23681 10919 23715
rect 10919 23681 10928 23715
rect 10876 23672 10928 23681
rect 15292 23817 15301 23851
rect 15301 23817 15335 23851
rect 15335 23817 15344 23851
rect 15292 23808 15344 23817
rect 16396 23851 16448 23860
rect 16396 23817 16405 23851
rect 16405 23817 16439 23851
rect 16439 23817 16448 23851
rect 16396 23808 16448 23817
rect 17132 23808 17184 23860
rect 17408 23808 17460 23860
rect 18696 23851 18748 23860
rect 18696 23817 18705 23851
rect 18705 23817 18739 23851
rect 18739 23817 18748 23851
rect 18696 23808 18748 23817
rect 20996 23808 21048 23860
rect 22008 23851 22060 23860
rect 22008 23817 22017 23851
rect 22017 23817 22051 23851
rect 22051 23817 22060 23851
rect 22008 23808 22060 23817
rect 12440 23715 12492 23724
rect 12440 23681 12449 23715
rect 12449 23681 12483 23715
rect 12483 23681 12492 23715
rect 12440 23672 12492 23681
rect 22652 23740 22704 23792
rect 1400 23604 1452 23656
rect 2504 23579 2556 23588
rect 2504 23545 2513 23579
rect 2513 23545 2547 23579
rect 2547 23545 2556 23579
rect 2504 23536 2556 23545
rect 3056 23604 3108 23656
rect 4988 23647 5040 23656
rect 4988 23613 4997 23647
rect 4997 23613 5031 23647
rect 5031 23613 5040 23647
rect 4988 23604 5040 23613
rect 6000 23604 6052 23656
rect 7196 23647 7248 23656
rect 7196 23613 7205 23647
rect 7205 23613 7239 23647
rect 7239 23613 7248 23647
rect 7196 23604 7248 23613
rect 8668 23647 8720 23656
rect 8668 23613 8702 23647
rect 8702 23613 8720 23647
rect 8668 23604 8720 23613
rect 3516 23536 3568 23588
rect 7380 23579 7432 23588
rect 7380 23545 7389 23579
rect 7389 23545 7423 23579
rect 7423 23545 7432 23579
rect 7380 23536 7432 23545
rect 7472 23579 7524 23588
rect 7472 23545 7481 23579
rect 7481 23545 7515 23579
rect 7515 23545 7524 23579
rect 7472 23536 7524 23545
rect 11060 23536 11112 23588
rect 12072 23536 12124 23588
rect 1952 23511 2004 23520
rect 1952 23477 1961 23511
rect 1961 23477 1995 23511
rect 1995 23477 2004 23511
rect 1952 23468 2004 23477
rect 6276 23468 6328 23520
rect 7656 23468 7708 23520
rect 8116 23468 8168 23520
rect 9772 23511 9824 23520
rect 9772 23477 9781 23511
rect 9781 23477 9815 23511
rect 9815 23477 9824 23511
rect 9772 23468 9824 23477
rect 11152 23468 11204 23520
rect 13820 23511 13872 23520
rect 13820 23477 13829 23511
rect 13829 23477 13863 23511
rect 13863 23477 13872 23511
rect 13820 23468 13872 23477
rect 14188 23468 14240 23520
rect 14280 23468 14332 23520
rect 14740 23468 14792 23520
rect 16856 23647 16908 23656
rect 16856 23613 16865 23647
rect 16865 23613 16899 23647
rect 16899 23613 16908 23647
rect 16856 23604 16908 23613
rect 18512 23647 18564 23656
rect 18512 23613 18521 23647
rect 18521 23613 18555 23647
rect 18555 23613 18564 23647
rect 18512 23604 18564 23613
rect 20720 23647 20772 23656
rect 20720 23613 20729 23647
rect 20729 23613 20763 23647
rect 20763 23613 20772 23647
rect 20720 23604 20772 23613
rect 21824 23647 21876 23656
rect 21824 23613 21833 23647
rect 21833 23613 21867 23647
rect 21867 23613 21876 23647
rect 21824 23604 21876 23613
rect 19524 23511 19576 23520
rect 19524 23477 19533 23511
rect 19533 23477 19567 23511
rect 19567 23477 19576 23511
rect 19524 23468 19576 23477
rect 20168 23511 20220 23520
rect 20168 23477 20177 23511
rect 20177 23477 20211 23511
rect 20211 23477 20220 23511
rect 20168 23468 20220 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1676 23307 1728 23316
rect 1676 23273 1685 23307
rect 1685 23273 1719 23307
rect 1719 23273 1728 23307
rect 1676 23264 1728 23273
rect 1952 23307 2004 23316
rect 1952 23273 1961 23307
rect 1961 23273 1995 23307
rect 1995 23273 2004 23307
rect 1952 23264 2004 23273
rect 4436 23264 4488 23316
rect 5172 23264 5224 23316
rect 5540 23264 5592 23316
rect 7472 23264 7524 23316
rect 8668 23264 8720 23316
rect 10048 23264 10100 23316
rect 13820 23264 13872 23316
rect 17868 23264 17920 23316
rect 19248 23264 19300 23316
rect 22008 23307 22060 23316
rect 22008 23273 22017 23307
rect 22017 23273 22051 23307
rect 22051 23273 22060 23307
rect 22008 23264 22060 23273
rect 2872 23128 2924 23180
rect 3056 23239 3108 23248
rect 3056 23205 3065 23239
rect 3065 23205 3099 23239
rect 3099 23205 3108 23239
rect 3056 23196 3108 23205
rect 5908 23239 5960 23248
rect 5908 23205 5917 23239
rect 5917 23205 5951 23239
rect 5951 23205 5960 23239
rect 5908 23196 5960 23205
rect 12072 23196 12124 23248
rect 12716 23239 12768 23248
rect 12716 23205 12725 23239
rect 12725 23205 12759 23239
rect 12759 23205 12768 23239
rect 12716 23196 12768 23205
rect 4252 23128 4304 23180
rect 4620 23128 4672 23180
rect 7104 23171 7156 23180
rect 7104 23137 7113 23171
rect 7113 23137 7147 23171
rect 7147 23137 7156 23171
rect 7104 23128 7156 23137
rect 7380 23171 7432 23180
rect 7380 23137 7414 23171
rect 7414 23137 7432 23171
rect 7380 23128 7432 23137
rect 8116 23128 8168 23180
rect 10048 23171 10100 23180
rect 10048 23137 10057 23171
rect 10057 23137 10091 23171
rect 10091 23137 10100 23171
rect 10048 23128 10100 23137
rect 11796 23128 11848 23180
rect 2964 23103 3016 23112
rect 2964 23069 2973 23103
rect 2973 23069 3007 23103
rect 3007 23069 3016 23103
rect 2964 23060 3016 23069
rect 6276 23060 6328 23112
rect 11060 23060 11112 23112
rect 4896 22992 4948 23044
rect 10600 23035 10652 23044
rect 10600 23001 10609 23035
rect 10609 23001 10643 23035
rect 10643 23001 10652 23035
rect 10600 22992 10652 23001
rect 15936 23196 15988 23248
rect 14648 23128 14700 23180
rect 14464 23060 14516 23112
rect 15844 23103 15896 23112
rect 15844 23069 15853 23103
rect 15853 23069 15887 23103
rect 15887 23069 15896 23103
rect 15844 23060 15896 23069
rect 16764 23128 16816 23180
rect 17960 23171 18012 23180
rect 17960 23137 17969 23171
rect 17969 23137 18003 23171
rect 18003 23137 18012 23171
rect 17960 23128 18012 23137
rect 21732 23128 21784 23180
rect 6736 22924 6788 22976
rect 13728 22967 13780 22976
rect 13728 22933 13737 22967
rect 13737 22933 13771 22967
rect 13771 22933 13780 22967
rect 13728 22924 13780 22933
rect 15384 22967 15436 22976
rect 15384 22933 15393 22967
rect 15393 22933 15427 22967
rect 15427 22933 15436 22967
rect 15384 22924 15436 22933
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2964 22720 3016 22772
rect 3976 22720 4028 22772
rect 4160 22720 4212 22772
rect 5540 22720 5592 22772
rect 6000 22720 6052 22772
rect 6920 22720 6972 22772
rect 7104 22763 7156 22772
rect 7104 22729 7113 22763
rect 7113 22729 7147 22763
rect 7147 22729 7156 22763
rect 7104 22720 7156 22729
rect 7196 22720 7248 22772
rect 4896 22695 4948 22704
rect 4896 22661 4905 22695
rect 4905 22661 4939 22695
rect 4939 22661 4948 22695
rect 4896 22652 4948 22661
rect 6276 22652 6328 22704
rect 7380 22652 7432 22704
rect 3608 22584 3660 22636
rect 7012 22584 7064 22636
rect 8668 22720 8720 22772
rect 9772 22763 9824 22772
rect 9772 22729 9781 22763
rect 9781 22729 9815 22763
rect 9815 22729 9824 22763
rect 9772 22720 9824 22729
rect 10048 22763 10100 22772
rect 10048 22729 10057 22763
rect 10057 22729 10091 22763
rect 10091 22729 10100 22763
rect 10048 22720 10100 22729
rect 11060 22763 11112 22772
rect 11060 22729 11069 22763
rect 11069 22729 11103 22763
rect 11103 22729 11112 22763
rect 11060 22720 11112 22729
rect 12716 22720 12768 22772
rect 14464 22720 14516 22772
rect 14648 22720 14700 22772
rect 16028 22720 16080 22772
rect 17960 22720 18012 22772
rect 21732 22720 21784 22772
rect 11796 22695 11848 22704
rect 11796 22661 11805 22695
rect 11805 22661 11839 22695
rect 11839 22661 11848 22695
rect 11796 22652 11848 22661
rect 12072 22695 12124 22704
rect 12072 22661 12081 22695
rect 12081 22661 12115 22695
rect 12115 22661 12124 22695
rect 12072 22652 12124 22661
rect 12440 22652 12492 22704
rect 15016 22652 15068 22704
rect 3516 22516 3568 22568
rect 5172 22559 5224 22568
rect 5172 22525 5181 22559
rect 5181 22525 5215 22559
rect 5215 22525 5224 22559
rect 5172 22516 5224 22525
rect 6736 22516 6788 22568
rect 9956 22516 10008 22568
rect 12624 22516 12676 22568
rect 2688 22448 2740 22500
rect 3792 22448 3844 22500
rect 7748 22491 7800 22500
rect 7748 22457 7757 22491
rect 7757 22457 7791 22491
rect 7791 22457 7800 22491
rect 7748 22448 7800 22457
rect 16304 22516 16356 22568
rect 4160 22380 4212 22432
rect 14188 22448 14240 22500
rect 15844 22448 15896 22500
rect 10692 22380 10744 22432
rect 16028 22423 16080 22432
rect 16028 22389 16037 22423
rect 16037 22389 16071 22423
rect 16071 22389 16080 22423
rect 16028 22380 16080 22389
rect 16212 22380 16264 22432
rect 16764 22380 16816 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2044 22176 2096 22228
rect 4896 22176 4948 22228
rect 2872 22108 2924 22160
rect 3148 22108 3200 22160
rect 5540 22108 5592 22160
rect 6828 22176 6880 22228
rect 7748 22176 7800 22228
rect 9956 22219 10008 22228
rect 9956 22185 9965 22219
rect 9965 22185 9999 22219
rect 9999 22185 10008 22219
rect 9956 22176 10008 22185
rect 13820 22176 13872 22228
rect 14188 22219 14240 22228
rect 14188 22185 14197 22219
rect 14197 22185 14231 22219
rect 14231 22185 14240 22219
rect 14188 22176 14240 22185
rect 14280 22176 14332 22228
rect 15016 22219 15068 22228
rect 15016 22185 15025 22219
rect 15025 22185 15059 22219
rect 15059 22185 15068 22219
rect 15016 22176 15068 22185
rect 15844 22219 15896 22228
rect 15844 22185 15853 22219
rect 15853 22185 15887 22219
rect 15887 22185 15896 22219
rect 15844 22176 15896 22185
rect 16304 22219 16356 22228
rect 16304 22185 16313 22219
rect 16313 22185 16347 22219
rect 16347 22185 16356 22219
rect 16304 22176 16356 22185
rect 4068 22040 4120 22092
rect 8208 22108 8260 22160
rect 7012 22083 7064 22092
rect 2964 22015 3016 22024
rect 2964 21981 2973 22015
rect 2973 21981 3007 22015
rect 3007 21981 3016 22015
rect 2964 21972 3016 21981
rect 3056 22015 3108 22024
rect 3056 21981 3065 22015
rect 3065 21981 3099 22015
rect 3099 21981 3108 22015
rect 3056 21972 3108 21981
rect 2504 21947 2556 21956
rect 2504 21913 2513 21947
rect 2513 21913 2547 21947
rect 2547 21913 2556 21947
rect 2504 21904 2556 21913
rect 2596 21904 2648 21956
rect 7012 22049 7021 22083
rect 7021 22049 7055 22083
rect 7055 22049 7064 22083
rect 7012 22040 7064 22049
rect 8116 22040 8168 22092
rect 9864 22040 9916 22092
rect 10508 22083 10560 22092
rect 10508 22049 10517 22083
rect 10517 22049 10551 22083
rect 10551 22049 10560 22083
rect 10508 22040 10560 22049
rect 10784 22040 10836 22092
rect 12624 22083 12676 22092
rect 12624 22049 12633 22083
rect 12633 22049 12667 22083
rect 12667 22049 12676 22083
rect 12624 22040 12676 22049
rect 13452 22040 13504 22092
rect 14464 22040 14516 22092
rect 15384 22040 15436 22092
rect 16212 22040 16264 22092
rect 16948 22040 17000 22092
rect 5632 22015 5684 22024
rect 5632 21981 5641 22015
rect 5641 21981 5675 22015
rect 5675 21981 5684 22015
rect 5632 21972 5684 21981
rect 2688 21836 2740 21888
rect 7380 21972 7432 22024
rect 10600 21972 10652 22024
rect 11888 21904 11940 21956
rect 13084 21904 13136 21956
rect 16028 21972 16080 22024
rect 17040 21947 17092 21956
rect 17040 21913 17049 21947
rect 17049 21913 17083 21947
rect 17083 21913 17092 21947
rect 17040 21904 17092 21913
rect 6276 21836 6328 21888
rect 6736 21879 6788 21888
rect 6736 21845 6745 21879
rect 6745 21845 6779 21879
rect 6779 21845 6788 21879
rect 6736 21836 6788 21845
rect 9036 21879 9088 21888
rect 9036 21845 9045 21879
rect 9045 21845 9079 21879
rect 9079 21845 9088 21879
rect 9036 21836 9088 21845
rect 9404 21879 9456 21888
rect 9404 21845 9413 21879
rect 9413 21845 9447 21879
rect 9447 21845 9456 21879
rect 9404 21836 9456 21845
rect 10876 21836 10928 21888
rect 11428 21836 11480 21888
rect 11796 21836 11848 21888
rect 15384 21879 15436 21888
rect 15384 21845 15393 21879
rect 15393 21845 15427 21879
rect 15427 21845 15436 21879
rect 15384 21836 15436 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 5540 21675 5592 21684
rect 5540 21641 5549 21675
rect 5549 21641 5583 21675
rect 5583 21641 5592 21675
rect 5540 21632 5592 21641
rect 7012 21632 7064 21684
rect 8208 21632 8260 21684
rect 9128 21675 9180 21684
rect 9128 21641 9137 21675
rect 9137 21641 9171 21675
rect 9171 21641 9180 21675
rect 9128 21632 9180 21641
rect 10692 21675 10744 21684
rect 10692 21641 10701 21675
rect 10701 21641 10735 21675
rect 10735 21641 10744 21675
rect 10692 21632 10744 21641
rect 11888 21675 11940 21684
rect 11888 21641 11897 21675
rect 11897 21641 11931 21675
rect 11931 21641 11940 21675
rect 11888 21632 11940 21641
rect 12532 21675 12584 21684
rect 12532 21641 12541 21675
rect 12541 21641 12575 21675
rect 12575 21641 12584 21675
rect 12532 21632 12584 21641
rect 13360 21632 13412 21684
rect 13820 21675 13872 21684
rect 13820 21641 13829 21675
rect 13829 21641 13863 21675
rect 13863 21641 13872 21675
rect 13820 21632 13872 21641
rect 14464 21675 14516 21684
rect 14464 21641 14473 21675
rect 14473 21641 14507 21675
rect 14507 21641 14516 21675
rect 14464 21632 14516 21641
rect 14740 21632 14792 21684
rect 16948 21675 17000 21684
rect 16948 21641 16957 21675
rect 16957 21641 16991 21675
rect 16991 21641 17000 21675
rect 16948 21632 17000 21641
rect 18328 21675 18380 21684
rect 18328 21641 18337 21675
rect 18337 21641 18371 21675
rect 18371 21641 18380 21675
rect 18328 21632 18380 21641
rect 2964 21564 3016 21616
rect 7748 21564 7800 21616
rect 12440 21564 12492 21616
rect 13452 21607 13504 21616
rect 13452 21573 13461 21607
rect 13461 21573 13495 21607
rect 13495 21573 13504 21607
rect 13452 21564 13504 21573
rect 2504 21539 2556 21548
rect 2504 21505 2513 21539
rect 2513 21505 2547 21539
rect 2547 21505 2556 21539
rect 2504 21496 2556 21505
rect 3516 21471 3568 21480
rect 3516 21437 3525 21471
rect 3525 21437 3559 21471
rect 3559 21437 3568 21471
rect 3516 21428 3568 21437
rect 10508 21496 10560 21548
rect 3792 21471 3844 21480
rect 3792 21437 3826 21471
rect 3826 21437 3844 21471
rect 3792 21428 3844 21437
rect 7380 21428 7432 21480
rect 10048 21471 10100 21480
rect 10048 21437 10057 21471
rect 10057 21437 10091 21471
rect 10091 21437 10100 21471
rect 10048 21428 10100 21437
rect 13084 21471 13136 21480
rect 13084 21437 13093 21471
rect 13093 21437 13127 21471
rect 13127 21437 13136 21471
rect 13084 21428 13136 21437
rect 14740 21428 14792 21480
rect 18328 21428 18380 21480
rect 3056 21403 3108 21412
rect 3056 21369 3065 21403
rect 3065 21369 3099 21403
rect 3099 21369 3108 21403
rect 3056 21360 3108 21369
rect 1584 21292 1636 21344
rect 2596 21292 2648 21344
rect 9404 21403 9456 21412
rect 9404 21369 9413 21403
rect 9413 21369 9447 21403
rect 9447 21369 9456 21403
rect 9404 21360 9456 21369
rect 11244 21360 11296 21412
rect 11796 21360 11848 21412
rect 12532 21360 12584 21412
rect 15660 21360 15712 21412
rect 15752 21360 15804 21412
rect 26240 21360 26292 21412
rect 27620 21360 27672 21412
rect 5264 21292 5316 21344
rect 6000 21292 6052 21344
rect 6828 21292 6880 21344
rect 6920 21292 6972 21344
rect 9036 21292 9088 21344
rect 10692 21292 10744 21344
rect 11060 21292 11112 21344
rect 11336 21292 11388 21344
rect 15016 21292 15068 21344
rect 15384 21292 15436 21344
rect 16028 21335 16080 21344
rect 16028 21301 16037 21335
rect 16037 21301 16071 21335
rect 16071 21301 16080 21335
rect 16028 21292 16080 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 2320 21088 2372 21140
rect 3792 21088 3844 21140
rect 4252 21131 4304 21140
rect 4252 21097 4261 21131
rect 4261 21097 4295 21131
rect 4295 21097 4304 21131
rect 4252 21088 4304 21097
rect 5448 21088 5500 21140
rect 6276 21131 6328 21140
rect 6276 21097 6285 21131
rect 6285 21097 6319 21131
rect 6319 21097 6328 21131
rect 6276 21088 6328 21097
rect 6920 21131 6972 21140
rect 6920 21097 6929 21131
rect 6929 21097 6963 21131
rect 6963 21097 6972 21131
rect 6920 21088 6972 21097
rect 10048 21088 10100 21140
rect 10784 21088 10836 21140
rect 11980 21088 12032 21140
rect 12532 21131 12584 21140
rect 12532 21097 12541 21131
rect 12541 21097 12575 21131
rect 12575 21097 12584 21131
rect 12532 21088 12584 21097
rect 13084 21088 13136 21140
rect 15016 21131 15068 21140
rect 15016 21097 15025 21131
rect 15025 21097 15059 21131
rect 15059 21097 15068 21131
rect 15016 21088 15068 21097
rect 15844 21088 15896 21140
rect 5264 21020 5316 21072
rect 7748 21063 7800 21072
rect 7748 21029 7757 21063
rect 7757 21029 7791 21063
rect 7791 21029 7800 21063
rect 7748 21020 7800 21029
rect 3516 20952 3568 21004
rect 4988 20952 5040 21004
rect 6736 20952 6788 21004
rect 10692 21020 10744 21072
rect 14188 21063 14240 21072
rect 14188 21029 14197 21063
rect 14197 21029 14231 21063
rect 14231 21029 14240 21063
rect 14188 21020 14240 21029
rect 14280 21063 14332 21072
rect 14280 21029 14289 21063
rect 14289 21029 14323 21063
rect 14323 21029 14332 21063
rect 14280 21020 14332 21029
rect 15660 21020 15712 21072
rect 16488 21020 16540 21072
rect 21916 21088 21968 21140
rect 9956 20995 10008 21004
rect 9956 20961 9990 20995
rect 9990 20961 10008 20995
rect 9956 20952 10008 20961
rect 14096 20952 14148 21004
rect 15752 20952 15804 21004
rect 15936 20995 15988 21004
rect 15936 20961 15970 20995
rect 15970 20961 15988 20995
rect 15936 20952 15988 20961
rect 20904 20995 20956 21004
rect 20904 20961 20913 20995
rect 20913 20961 20947 20995
rect 20947 20961 20956 20995
rect 20904 20952 20956 20961
rect 2320 20927 2372 20936
rect 2320 20893 2329 20927
rect 2329 20893 2363 20927
rect 2363 20893 2372 20927
rect 2320 20884 2372 20893
rect 2688 20884 2740 20936
rect 8300 20884 8352 20936
rect 15660 20927 15712 20936
rect 15660 20893 15669 20927
rect 15669 20893 15703 20927
rect 15703 20893 15712 20927
rect 15660 20884 15712 20893
rect 9036 20816 9088 20868
rect 1860 20748 1912 20800
rect 2504 20748 2556 20800
rect 3700 20748 3752 20800
rect 7380 20748 7432 20800
rect 9588 20748 9640 20800
rect 12900 20791 12952 20800
rect 12900 20757 12909 20791
rect 12909 20757 12943 20791
rect 12943 20757 12952 20791
rect 12900 20748 12952 20757
rect 13636 20748 13688 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 2412 20544 2464 20596
rect 3056 20544 3108 20596
rect 4620 20544 4672 20596
rect 6276 20587 6328 20596
rect 6276 20553 6285 20587
rect 6285 20553 6319 20587
rect 6319 20553 6328 20587
rect 6276 20544 6328 20553
rect 4436 20476 4488 20528
rect 4712 20519 4764 20528
rect 4712 20485 4721 20519
rect 4721 20485 4755 20519
rect 4755 20485 4764 20519
rect 4712 20476 4764 20485
rect 3608 20451 3660 20460
rect 3608 20417 3617 20451
rect 3617 20417 3651 20451
rect 3651 20417 3660 20451
rect 3608 20408 3660 20417
rect 5448 20408 5500 20460
rect 1860 20383 1912 20392
rect 1860 20349 1869 20383
rect 1869 20349 1903 20383
rect 1903 20349 1912 20383
rect 1860 20340 1912 20349
rect 3700 20383 3752 20392
rect 3700 20349 3709 20383
rect 3709 20349 3743 20383
rect 3743 20349 3752 20383
rect 3700 20340 3752 20349
rect 4988 20340 5040 20392
rect 7104 20544 7156 20596
rect 8300 20544 8352 20596
rect 9404 20587 9456 20596
rect 9404 20553 9413 20587
rect 9413 20553 9447 20587
rect 9447 20553 9456 20587
rect 9404 20544 9456 20553
rect 10968 20544 11020 20596
rect 11244 20544 11296 20596
rect 13452 20544 13504 20596
rect 14096 20587 14148 20596
rect 14096 20553 14105 20587
rect 14105 20553 14139 20587
rect 14139 20553 14148 20587
rect 14096 20544 14148 20553
rect 14280 20544 14332 20596
rect 12532 20519 12584 20528
rect 12532 20485 12541 20519
rect 12541 20485 12575 20519
rect 12575 20485 12584 20519
rect 12532 20476 12584 20485
rect 9956 20451 10008 20460
rect 9956 20417 9965 20451
rect 9965 20417 9999 20451
rect 9999 20417 10008 20451
rect 9956 20408 10008 20417
rect 12900 20408 12952 20460
rect 13728 20408 13780 20460
rect 18328 20451 18380 20460
rect 18328 20417 18337 20451
rect 18337 20417 18371 20451
rect 18371 20417 18380 20451
rect 18328 20408 18380 20417
rect 15660 20340 15712 20392
rect 18052 20383 18104 20392
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 2688 20272 2740 20324
rect 3148 20272 3200 20324
rect 6276 20272 6328 20324
rect 9680 20315 9732 20324
rect 9680 20281 9689 20315
rect 9689 20281 9723 20315
rect 9723 20281 9732 20315
rect 9680 20272 9732 20281
rect 12900 20272 12952 20324
rect 14280 20272 14332 20324
rect 1768 20204 1820 20256
rect 4160 20247 4212 20256
rect 4160 20213 4169 20247
rect 4169 20213 4203 20247
rect 4203 20213 4212 20247
rect 4160 20204 4212 20213
rect 4620 20204 4672 20256
rect 8208 20247 8260 20256
rect 8208 20213 8217 20247
rect 8217 20213 8251 20247
rect 8251 20213 8260 20247
rect 8208 20204 8260 20213
rect 9496 20204 9548 20256
rect 10692 20204 10744 20256
rect 11244 20204 11296 20256
rect 11796 20247 11848 20256
rect 11796 20213 11805 20247
rect 11805 20213 11839 20247
rect 11839 20213 11848 20247
rect 11796 20204 11848 20213
rect 11888 20204 11940 20256
rect 13452 20204 13504 20256
rect 16028 20204 16080 20256
rect 20904 20247 20956 20256
rect 20904 20213 20913 20247
rect 20913 20213 20947 20247
rect 20947 20213 20956 20247
rect 20904 20204 20956 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2320 20043 2372 20052
rect 2320 20009 2329 20043
rect 2329 20009 2363 20043
rect 2363 20009 2372 20043
rect 2320 20000 2372 20009
rect 3608 20000 3660 20052
rect 5264 20043 5316 20052
rect 5264 20009 5273 20043
rect 5273 20009 5307 20043
rect 5307 20009 5316 20043
rect 5264 20000 5316 20009
rect 6736 20000 6788 20052
rect 6920 20043 6972 20052
rect 6920 20009 6929 20043
rect 6929 20009 6963 20043
rect 6963 20009 6972 20043
rect 6920 20000 6972 20009
rect 8300 20000 8352 20052
rect 9956 20000 10008 20052
rect 10784 20043 10836 20052
rect 10784 20009 10793 20043
rect 10793 20009 10827 20043
rect 10827 20009 10836 20043
rect 10784 20000 10836 20009
rect 11060 20000 11112 20052
rect 11796 20000 11848 20052
rect 12900 20000 12952 20052
rect 15660 20043 15712 20052
rect 15660 20009 15669 20043
rect 15669 20009 15703 20043
rect 15703 20009 15712 20043
rect 15660 20000 15712 20009
rect 2964 19932 3016 19984
rect 4712 19975 4764 19984
rect 4712 19941 4721 19975
rect 4721 19941 4755 19975
rect 4755 19941 4764 19975
rect 4712 19932 4764 19941
rect 5172 19932 5224 19984
rect 10232 19932 10284 19984
rect 12808 19932 12860 19984
rect 14188 19975 14240 19984
rect 14188 19941 14197 19975
rect 14197 19941 14231 19975
rect 14231 19941 14240 19975
rect 14188 19932 14240 19941
rect 14280 19975 14332 19984
rect 14280 19941 14289 19975
rect 14289 19941 14323 19975
rect 14323 19941 14332 19975
rect 14280 19932 14332 19941
rect 7104 19907 7156 19916
rect 7104 19873 7113 19907
rect 7113 19873 7147 19907
rect 7147 19873 7156 19907
rect 7104 19864 7156 19873
rect 7380 19907 7432 19916
rect 7380 19873 7414 19907
rect 7414 19873 7432 19907
rect 7380 19864 7432 19873
rect 8208 19864 8260 19916
rect 11244 19864 11296 19916
rect 11428 19907 11480 19916
rect 11428 19873 11462 19907
rect 11462 19873 11480 19907
rect 11428 19864 11480 19873
rect 13820 19864 13872 19916
rect 16488 19975 16540 19984
rect 16488 19941 16522 19975
rect 16522 19941 16540 19975
rect 16488 19932 16540 19941
rect 20904 19932 20956 19984
rect 16304 19864 16356 19916
rect 19156 19907 19208 19916
rect 19156 19873 19165 19907
rect 19165 19873 19199 19907
rect 19199 19873 19208 19907
rect 19156 19864 19208 19873
rect 4804 19839 4856 19848
rect 4804 19805 4813 19839
rect 4813 19805 4847 19839
rect 4847 19805 4856 19839
rect 4804 19796 4856 19805
rect 9772 19796 9824 19848
rect 5448 19728 5500 19780
rect 15844 19728 15896 19780
rect 16120 19728 16172 19780
rect 17592 19771 17644 19780
rect 17592 19737 17601 19771
rect 17601 19737 17635 19771
rect 17635 19737 17644 19771
rect 17592 19728 17644 19737
rect 1768 19660 1820 19712
rect 2688 19703 2740 19712
rect 2688 19669 2697 19703
rect 2697 19669 2731 19703
rect 2731 19669 2740 19703
rect 2688 19660 2740 19669
rect 3792 19703 3844 19712
rect 3792 19669 3801 19703
rect 3801 19669 3835 19703
rect 3835 19669 3844 19703
rect 3792 19660 3844 19669
rect 4252 19703 4304 19712
rect 4252 19669 4261 19703
rect 4261 19669 4295 19703
rect 4295 19669 4304 19703
rect 4252 19660 4304 19669
rect 9496 19660 9548 19712
rect 9864 19660 9916 19712
rect 12900 19660 12952 19712
rect 13728 19703 13780 19712
rect 13728 19669 13737 19703
rect 13737 19669 13771 19703
rect 13771 19669 13780 19703
rect 13728 19660 13780 19669
rect 15568 19660 15620 19712
rect 16028 19703 16080 19712
rect 16028 19669 16037 19703
rect 16037 19669 16071 19703
rect 16071 19669 16080 19703
rect 16028 19660 16080 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2688 19456 2740 19508
rect 5172 19499 5224 19508
rect 5172 19465 5181 19499
rect 5181 19465 5215 19499
rect 5215 19465 5224 19499
rect 5172 19456 5224 19465
rect 7104 19456 7156 19508
rect 9680 19456 9732 19508
rect 11796 19456 11848 19508
rect 13360 19456 13412 19508
rect 13820 19456 13872 19508
rect 14740 19456 14792 19508
rect 16304 19499 16356 19508
rect 16304 19465 16313 19499
rect 16313 19465 16347 19499
rect 16347 19465 16356 19499
rect 16304 19456 16356 19465
rect 16488 19456 16540 19508
rect 14464 19388 14516 19440
rect 2780 19320 2832 19372
rect 3792 19320 3844 19372
rect 2412 19252 2464 19304
rect 4344 19320 4396 19372
rect 4804 19363 4856 19372
rect 4804 19329 4813 19363
rect 4813 19329 4847 19363
rect 4847 19329 4856 19363
rect 4804 19320 4856 19329
rect 5632 19295 5684 19304
rect 5632 19261 5641 19295
rect 5641 19261 5675 19295
rect 5675 19261 5684 19295
rect 5632 19252 5684 19261
rect 8208 19320 8260 19372
rect 6920 19252 6972 19304
rect 9036 19252 9088 19304
rect 9772 19320 9824 19372
rect 13452 19320 13504 19372
rect 10600 19295 10652 19304
rect 10600 19261 10609 19295
rect 10609 19261 10643 19295
rect 10643 19261 10652 19295
rect 10600 19252 10652 19261
rect 11244 19252 11296 19304
rect 12348 19252 12400 19304
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 21548 19252 21600 19304
rect 2320 19184 2372 19236
rect 4068 19184 4120 19236
rect 4252 19184 4304 19236
rect 2964 19116 3016 19168
rect 3332 19159 3384 19168
rect 3332 19125 3341 19159
rect 3341 19125 3375 19159
rect 3375 19125 3384 19159
rect 3332 19116 3384 19125
rect 6000 19184 6052 19236
rect 7564 19184 7616 19236
rect 8208 19184 8260 19236
rect 10048 19184 10100 19236
rect 10232 19184 10284 19236
rect 11152 19227 11204 19236
rect 11152 19193 11161 19227
rect 11161 19193 11195 19227
rect 11195 19193 11204 19227
rect 11152 19184 11204 19193
rect 11428 19227 11480 19236
rect 11428 19193 11437 19227
rect 11437 19193 11471 19227
rect 11471 19193 11480 19227
rect 11428 19184 11480 19193
rect 12900 19184 12952 19236
rect 15476 19227 15528 19236
rect 15476 19193 15485 19227
rect 15485 19193 15519 19227
rect 15519 19193 15528 19227
rect 15476 19184 15528 19193
rect 15568 19227 15620 19236
rect 15568 19193 15577 19227
rect 15577 19193 15611 19227
rect 15611 19193 15620 19227
rect 15568 19184 15620 19193
rect 5448 19116 5500 19168
rect 7104 19116 7156 19168
rect 8760 19159 8812 19168
rect 8760 19125 8769 19159
rect 8769 19125 8803 19159
rect 8803 19125 8812 19159
rect 8760 19116 8812 19125
rect 9772 19116 9824 19168
rect 11060 19116 11112 19168
rect 12348 19116 12400 19168
rect 12624 19116 12676 19168
rect 13820 19159 13872 19168
rect 13820 19125 13829 19159
rect 13829 19125 13863 19159
rect 13863 19125 13872 19159
rect 13820 19116 13872 19125
rect 14280 19116 14332 19168
rect 15016 19116 15068 19168
rect 19156 19159 19208 19168
rect 19156 19125 19165 19159
rect 19165 19125 19199 19159
rect 19199 19125 19208 19159
rect 19156 19116 19208 19125
rect 23388 19116 23440 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2320 18955 2372 18964
rect 2320 18921 2329 18955
rect 2329 18921 2363 18955
rect 2363 18921 2372 18955
rect 2320 18912 2372 18921
rect 4252 18912 4304 18964
rect 5448 18955 5500 18964
rect 5448 18921 5457 18955
rect 5457 18921 5491 18955
rect 5491 18921 5500 18955
rect 5448 18912 5500 18921
rect 7564 18955 7616 18964
rect 7564 18921 7573 18955
rect 7573 18921 7607 18955
rect 7607 18921 7616 18955
rect 7564 18912 7616 18921
rect 9036 18955 9088 18964
rect 9036 18921 9045 18955
rect 9045 18921 9079 18955
rect 9079 18921 9088 18955
rect 9036 18912 9088 18921
rect 11428 18912 11480 18964
rect 15016 18955 15068 18964
rect 15016 18921 15025 18955
rect 15025 18921 15059 18955
rect 15059 18921 15068 18955
rect 15016 18912 15068 18921
rect 15476 18912 15528 18964
rect 2504 18844 2556 18896
rect 3332 18844 3384 18896
rect 4160 18844 4212 18896
rect 7104 18887 7156 18896
rect 7104 18853 7113 18887
rect 7113 18853 7147 18887
rect 7147 18853 7156 18887
rect 7104 18844 7156 18853
rect 10692 18844 10744 18896
rect 11244 18887 11296 18896
rect 11244 18853 11253 18887
rect 11253 18853 11287 18887
rect 11287 18853 11296 18887
rect 11244 18844 11296 18853
rect 14740 18844 14792 18896
rect 15936 18887 15988 18896
rect 15936 18853 15945 18887
rect 15945 18853 15979 18887
rect 15979 18853 15988 18887
rect 15936 18844 15988 18853
rect 2412 18776 2464 18828
rect 4344 18819 4396 18828
rect 4344 18785 4367 18819
rect 4367 18785 4396 18819
rect 4344 18776 4396 18785
rect 6920 18819 6972 18828
rect 6920 18785 6929 18819
rect 6929 18785 6963 18819
rect 6963 18785 6972 18819
rect 6920 18776 6972 18785
rect 10048 18776 10100 18828
rect 11888 18776 11940 18828
rect 13820 18776 13872 18828
rect 15660 18819 15712 18828
rect 15660 18785 15669 18819
rect 15669 18785 15703 18819
rect 15703 18785 15712 18819
rect 15660 18776 15712 18785
rect 3056 18751 3108 18760
rect 3056 18717 3065 18751
rect 3065 18717 3099 18751
rect 3099 18717 3108 18751
rect 3056 18708 3108 18717
rect 3516 18708 3568 18760
rect 7380 18708 7432 18760
rect 10232 18751 10284 18760
rect 10232 18717 10241 18751
rect 10241 18717 10275 18751
rect 10275 18717 10284 18751
rect 10232 18708 10284 18717
rect 12716 18751 12768 18760
rect 12716 18717 12725 18751
rect 12725 18717 12759 18751
rect 12759 18717 12768 18751
rect 12716 18708 12768 18717
rect 2780 18640 2832 18692
rect 9864 18640 9916 18692
rect 2964 18572 3016 18624
rect 4252 18572 4304 18624
rect 6828 18572 6880 18624
rect 11336 18572 11388 18624
rect 12900 18572 12952 18624
rect 13084 18572 13136 18624
rect 15384 18615 15436 18624
rect 15384 18581 15393 18615
rect 15393 18581 15427 18615
rect 15427 18581 15436 18615
rect 15384 18572 15436 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 3056 18368 3108 18420
rect 3516 18368 3568 18420
rect 4344 18368 4396 18420
rect 7104 18368 7156 18420
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 12532 18411 12584 18420
rect 12532 18377 12541 18411
rect 12541 18377 12575 18411
rect 12575 18377 12584 18411
rect 12532 18368 12584 18377
rect 12716 18368 12768 18420
rect 13452 18368 13504 18420
rect 13912 18368 13964 18420
rect 14740 18368 14792 18420
rect 15752 18368 15804 18420
rect 2320 18232 2372 18284
rect 4160 18300 4212 18352
rect 6368 18300 6420 18352
rect 7932 18300 7984 18352
rect 9588 18300 9640 18352
rect 10876 18343 10928 18352
rect 10876 18309 10885 18343
rect 10885 18309 10919 18343
rect 10919 18309 10928 18343
rect 10876 18300 10928 18309
rect 3056 18164 3108 18216
rect 7380 18232 7432 18284
rect 9220 18232 9272 18284
rect 10968 18232 11020 18284
rect 11336 18275 11388 18284
rect 11336 18241 11345 18275
rect 11345 18241 11379 18275
rect 11379 18241 11388 18275
rect 11336 18232 11388 18241
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 15384 18232 15436 18284
rect 5448 18164 5500 18216
rect 2504 18096 2556 18148
rect 8116 18164 8168 18216
rect 9680 18096 9732 18148
rect 10232 18139 10284 18148
rect 10232 18105 10241 18139
rect 10241 18105 10275 18139
rect 10275 18105 10284 18139
rect 10232 18096 10284 18105
rect 12256 18096 12308 18148
rect 14096 18164 14148 18216
rect 15936 18232 15988 18284
rect 21548 18275 21600 18284
rect 21548 18241 21557 18275
rect 21557 18241 21591 18275
rect 21591 18241 21600 18275
rect 21548 18232 21600 18241
rect 2688 18028 2740 18080
rect 9772 18071 9824 18080
rect 9772 18037 9781 18071
rect 9781 18037 9815 18071
rect 9815 18037 9824 18071
rect 9772 18028 9824 18037
rect 11336 18071 11388 18080
rect 11336 18037 11345 18071
rect 11345 18037 11379 18071
rect 11379 18037 11388 18071
rect 11336 18028 11388 18037
rect 12072 18028 12124 18080
rect 12900 18096 12952 18148
rect 12992 18071 13044 18080
rect 12992 18037 13001 18071
rect 13001 18037 13035 18071
rect 13035 18037 13044 18071
rect 12992 18028 13044 18037
rect 13452 18071 13504 18080
rect 13452 18037 13461 18071
rect 13461 18037 13495 18071
rect 13495 18037 13504 18071
rect 13452 18028 13504 18037
rect 14188 18096 14240 18148
rect 21272 18207 21324 18216
rect 21272 18173 21281 18207
rect 21281 18173 21315 18207
rect 21315 18173 21324 18207
rect 21272 18164 21324 18173
rect 15384 18139 15436 18148
rect 15384 18105 15393 18139
rect 15393 18105 15427 18139
rect 15427 18105 15436 18139
rect 15384 18096 15436 18105
rect 16120 18139 16172 18148
rect 16120 18105 16129 18139
rect 16129 18105 16163 18139
rect 16163 18105 16172 18139
rect 16120 18096 16172 18105
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2412 17824 2464 17876
rect 3516 17824 3568 17876
rect 4436 17824 4488 17876
rect 7380 17867 7432 17876
rect 2780 17756 2832 17808
rect 3056 17799 3108 17808
rect 3056 17765 3065 17799
rect 3065 17765 3099 17799
rect 3099 17765 3108 17799
rect 5356 17799 5408 17808
rect 3056 17756 3108 17765
rect 5356 17765 5390 17799
rect 5390 17765 5408 17799
rect 5356 17756 5408 17765
rect 6276 17756 6328 17808
rect 7380 17833 7389 17867
rect 7389 17833 7423 17867
rect 7423 17833 7432 17867
rect 7380 17824 7432 17833
rect 9220 17867 9272 17876
rect 9220 17833 9229 17867
rect 9229 17833 9263 17867
rect 9263 17833 9272 17867
rect 9220 17824 9272 17833
rect 10048 17824 10100 17876
rect 11336 17824 11388 17876
rect 11888 17824 11940 17876
rect 12256 17824 12308 17876
rect 13360 17824 13412 17876
rect 14188 17867 14240 17876
rect 14188 17833 14197 17867
rect 14197 17833 14231 17867
rect 14231 17833 14240 17867
rect 14188 17824 14240 17833
rect 14556 17867 14608 17876
rect 14556 17833 14565 17867
rect 14565 17833 14599 17867
rect 14599 17833 14608 17867
rect 14556 17824 14608 17833
rect 7564 17756 7616 17808
rect 7932 17799 7984 17808
rect 7932 17765 7941 17799
rect 7941 17765 7975 17799
rect 7975 17765 7984 17799
rect 7932 17756 7984 17765
rect 6828 17688 6880 17740
rect 10232 17756 10284 17808
rect 12440 17756 12492 17808
rect 12992 17756 13044 17808
rect 13268 17799 13320 17808
rect 13268 17765 13277 17799
rect 13277 17765 13311 17799
rect 13311 17765 13320 17799
rect 13268 17756 13320 17765
rect 15844 17799 15896 17808
rect 15844 17765 15853 17799
rect 15853 17765 15887 17799
rect 15887 17765 15896 17799
rect 15844 17756 15896 17765
rect 15936 17799 15988 17808
rect 15936 17765 15945 17799
rect 15945 17765 15979 17799
rect 15979 17765 15988 17799
rect 15936 17756 15988 17765
rect 16396 17756 16448 17808
rect 9128 17688 9180 17740
rect 13084 17688 13136 17740
rect 15384 17688 15436 17740
rect 15752 17688 15804 17740
rect 2872 17663 2924 17672
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 2872 17620 2924 17629
rect 4436 17620 4488 17672
rect 8208 17663 8260 17672
rect 8208 17629 8217 17663
rect 8217 17629 8251 17663
rect 8251 17629 8260 17663
rect 8208 17620 8260 17629
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 11428 17620 11480 17672
rect 13176 17663 13228 17672
rect 13176 17629 13185 17663
rect 13185 17629 13219 17663
rect 13219 17629 13228 17663
rect 13176 17620 13228 17629
rect 2504 17595 2556 17604
rect 2504 17561 2513 17595
rect 2513 17561 2547 17595
rect 2547 17561 2556 17595
rect 2504 17552 2556 17561
rect 7656 17595 7708 17604
rect 7656 17561 7665 17595
rect 7665 17561 7699 17595
rect 7699 17561 7708 17595
rect 7656 17552 7708 17561
rect 15292 17552 15344 17604
rect 10692 17484 10744 17536
rect 12808 17527 12860 17536
rect 12808 17493 12817 17527
rect 12817 17493 12851 17527
rect 12851 17493 12860 17527
rect 12808 17484 12860 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2780 17280 2832 17332
rect 2872 17323 2924 17332
rect 2872 17289 2881 17323
rect 2881 17289 2915 17323
rect 2915 17289 2924 17323
rect 2872 17280 2924 17289
rect 3056 17280 3108 17332
rect 3884 17280 3936 17332
rect 5448 17280 5500 17332
rect 6276 17323 6328 17332
rect 6276 17289 6285 17323
rect 6285 17289 6319 17323
rect 6319 17289 6328 17323
rect 6276 17280 6328 17289
rect 8208 17280 8260 17332
rect 9128 17323 9180 17332
rect 9128 17289 9137 17323
rect 9137 17289 9171 17323
rect 9171 17289 9180 17323
rect 9128 17280 9180 17289
rect 10968 17280 11020 17332
rect 13084 17280 13136 17332
rect 15844 17280 15896 17332
rect 16396 17323 16448 17332
rect 16396 17289 16405 17323
rect 16405 17289 16439 17323
rect 16439 17289 16448 17323
rect 16396 17280 16448 17289
rect 5356 17212 5408 17264
rect 4436 17144 4488 17196
rect 5448 17144 5500 17196
rect 11244 17212 11296 17264
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 9772 17144 9824 17196
rect 10140 17144 10192 17196
rect 7104 17119 7156 17128
rect 7104 17085 7127 17119
rect 7127 17085 7156 17119
rect 7104 17076 7156 17085
rect 11152 17051 11204 17060
rect 1860 16940 1912 16992
rect 5724 16983 5776 16992
rect 5724 16949 5733 16983
rect 5733 16949 5767 16983
rect 5767 16949 5776 16983
rect 5724 16940 5776 16949
rect 11152 17017 11161 17051
rect 11161 17017 11195 17051
rect 11195 17017 11204 17051
rect 11152 17008 11204 17017
rect 11428 17051 11480 17060
rect 11428 17017 11437 17051
rect 11437 17017 11471 17051
rect 11471 17017 11480 17051
rect 11428 17008 11480 17017
rect 13360 17119 13412 17128
rect 13360 17085 13394 17119
rect 13394 17085 13412 17119
rect 13360 17076 13412 17085
rect 13452 17008 13504 17060
rect 7012 16940 7064 16992
rect 7380 16940 7432 16992
rect 10140 16940 10192 16992
rect 10876 16940 10928 16992
rect 11980 16940 12032 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 15292 16983 15344 16992
rect 15292 16949 15301 16983
rect 15301 16949 15335 16983
rect 15335 16949 15344 16983
rect 15292 16940 15344 16949
rect 15844 16940 15896 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 4160 16736 4212 16788
rect 4988 16736 5040 16788
rect 5724 16736 5776 16788
rect 8208 16736 8260 16788
rect 8760 16736 8812 16788
rect 9864 16736 9916 16788
rect 10876 16779 10928 16788
rect 6184 16668 6236 16720
rect 7380 16711 7432 16720
rect 7380 16677 7414 16711
rect 7414 16677 7432 16711
rect 7380 16668 7432 16677
rect 10048 16668 10100 16720
rect 10876 16745 10885 16779
rect 10885 16745 10919 16779
rect 10919 16745 10928 16779
rect 10876 16736 10928 16745
rect 11152 16779 11204 16788
rect 11152 16745 11161 16779
rect 11161 16745 11195 16779
rect 11195 16745 11204 16779
rect 11152 16736 11204 16745
rect 12440 16736 12492 16788
rect 13360 16736 13412 16788
rect 15476 16736 15528 16788
rect 11428 16668 11480 16720
rect 12716 16668 12768 16720
rect 13084 16668 13136 16720
rect 14004 16668 14056 16720
rect 2412 16643 2464 16652
rect 2412 16609 2421 16643
rect 2421 16609 2455 16643
rect 2455 16609 2464 16643
rect 2412 16600 2464 16609
rect 6828 16600 6880 16652
rect 11060 16600 11112 16652
rect 15568 16600 15620 16652
rect 1400 16464 1452 16516
rect 9404 16532 9456 16584
rect 10600 16532 10652 16584
rect 11888 16575 11940 16584
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 11888 16532 11940 16541
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 1308 16396 1360 16448
rect 5356 16396 5408 16448
rect 5540 16396 5592 16448
rect 7380 16396 7432 16448
rect 15292 16396 15344 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2228 16192 2280 16244
rect 4988 16235 5040 16244
rect 4988 16201 4997 16235
rect 4997 16201 5031 16235
rect 5031 16201 5040 16235
rect 4988 16192 5040 16201
rect 6920 16235 6972 16244
rect 6920 16201 6929 16235
rect 6929 16201 6963 16235
rect 6963 16201 6972 16235
rect 6920 16192 6972 16201
rect 10048 16192 10100 16244
rect 13268 16192 13320 16244
rect 15844 16192 15896 16244
rect 2504 16124 2556 16176
rect 5264 16167 5316 16176
rect 5264 16133 5273 16167
rect 5273 16133 5307 16167
rect 5307 16133 5316 16167
rect 5264 16124 5316 16133
rect 6368 16124 6420 16176
rect 6644 16124 6696 16176
rect 6828 16124 6880 16176
rect 10600 16167 10652 16176
rect 10600 16133 10609 16167
rect 10609 16133 10643 16167
rect 10643 16133 10652 16167
rect 10600 16124 10652 16133
rect 13176 16124 13228 16176
rect 2228 16056 2280 16108
rect 6000 16056 6052 16108
rect 7104 16056 7156 16108
rect 8668 16099 8720 16108
rect 8668 16065 8677 16099
rect 8677 16065 8711 16099
rect 8711 16065 8720 16099
rect 8668 16056 8720 16065
rect 11152 16099 11204 16108
rect 11152 16065 11161 16099
rect 11161 16065 11195 16099
rect 11195 16065 11204 16099
rect 11152 16056 11204 16065
rect 15476 16056 15528 16108
rect 1400 15988 1452 16040
rect 3700 15920 3752 15972
rect 6460 15988 6512 16040
rect 6644 15988 6696 16040
rect 8760 15988 8812 16040
rect 5816 15963 5868 15972
rect 5816 15929 5825 15963
rect 5825 15929 5859 15963
rect 5859 15929 5868 15963
rect 5816 15920 5868 15929
rect 1952 15852 2004 15904
rect 3240 15852 3292 15904
rect 3516 15895 3568 15904
rect 3516 15861 3525 15895
rect 3525 15861 3559 15895
rect 3559 15861 3568 15895
rect 3516 15852 3568 15861
rect 3884 15852 3936 15904
rect 6184 15895 6236 15904
rect 6184 15861 6193 15895
rect 6193 15861 6227 15895
rect 6227 15861 6236 15895
rect 7380 15963 7432 15972
rect 7380 15929 7389 15963
rect 7389 15929 7423 15963
rect 7423 15929 7432 15963
rect 7380 15920 7432 15929
rect 11888 15920 11940 15972
rect 12900 15920 12952 15972
rect 14004 15988 14056 16040
rect 16672 16031 16724 16040
rect 16672 15997 16681 16031
rect 16681 15997 16715 16031
rect 16715 15997 16724 16031
rect 16672 15988 16724 15997
rect 6184 15852 6236 15861
rect 9956 15852 10008 15904
rect 12716 15895 12768 15904
rect 12716 15861 12725 15895
rect 12725 15861 12759 15895
rect 12759 15861 12768 15895
rect 12716 15852 12768 15861
rect 18420 15920 18472 15972
rect 14556 15852 14608 15904
rect 15476 15852 15528 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 6000 15648 6052 15700
rect 7104 15648 7156 15700
rect 8760 15648 8812 15700
rect 11060 15648 11112 15700
rect 13820 15648 13872 15700
rect 14004 15648 14056 15700
rect 5816 15580 5868 15632
rect 7472 15580 7524 15632
rect 8116 15580 8168 15632
rect 8668 15580 8720 15632
rect 2044 15512 2096 15564
rect 2596 15512 2648 15564
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 6000 15512 6052 15564
rect 3332 15376 3384 15428
rect 8024 15512 8076 15564
rect 8300 15555 8352 15564
rect 8300 15521 8309 15555
rect 8309 15521 8343 15555
rect 8343 15521 8352 15555
rect 8300 15512 8352 15521
rect 10324 15580 10376 15632
rect 15936 15580 15988 15632
rect 17224 15623 17276 15632
rect 17224 15589 17233 15623
rect 17233 15589 17267 15623
rect 17267 15589 17276 15623
rect 17224 15580 17276 15589
rect 17408 15623 17460 15632
rect 17408 15589 17417 15623
rect 17417 15589 17451 15623
rect 17451 15589 17460 15623
rect 17408 15580 17460 15589
rect 9956 15555 10008 15564
rect 9956 15521 9990 15555
rect 9990 15521 10008 15555
rect 9956 15512 10008 15521
rect 12716 15512 12768 15564
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 2320 15351 2372 15360
rect 2320 15317 2329 15351
rect 2329 15317 2363 15351
rect 2363 15317 2372 15351
rect 2320 15308 2372 15317
rect 2688 15351 2740 15360
rect 2688 15317 2697 15351
rect 2697 15317 2731 15351
rect 2731 15317 2740 15351
rect 2688 15308 2740 15317
rect 3424 15351 3476 15360
rect 3424 15317 3433 15351
rect 3433 15317 3467 15351
rect 3467 15317 3476 15351
rect 3424 15308 3476 15317
rect 3792 15351 3844 15360
rect 3792 15317 3801 15351
rect 3801 15317 3835 15351
rect 3835 15317 3844 15351
rect 3792 15308 3844 15317
rect 7656 15308 7708 15360
rect 8760 15444 8812 15496
rect 13912 15487 13964 15496
rect 13912 15453 13921 15487
rect 13921 15453 13955 15487
rect 13955 15453 13964 15487
rect 13912 15444 13964 15453
rect 15292 15512 15344 15564
rect 18420 15555 18472 15564
rect 18420 15521 18429 15555
rect 18429 15521 18463 15555
rect 18463 15521 18472 15555
rect 18420 15512 18472 15521
rect 14556 15444 14608 15496
rect 16120 15444 16172 15496
rect 14372 15376 14424 15428
rect 15568 15376 15620 15428
rect 18236 15444 18288 15496
rect 8024 15351 8076 15360
rect 8024 15317 8033 15351
rect 8033 15317 8067 15351
rect 8067 15317 8076 15351
rect 8024 15308 8076 15317
rect 9864 15308 9916 15360
rect 11152 15308 11204 15360
rect 13084 15308 13136 15360
rect 15384 15351 15436 15360
rect 15384 15317 15393 15351
rect 15393 15317 15427 15351
rect 15427 15317 15436 15351
rect 15384 15308 15436 15317
rect 20260 15308 20312 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2044 15147 2096 15156
rect 2044 15113 2053 15147
rect 2053 15113 2087 15147
rect 2087 15113 2096 15147
rect 2044 15104 2096 15113
rect 2596 15147 2648 15156
rect 2596 15113 2605 15147
rect 2605 15113 2639 15147
rect 2639 15113 2648 15147
rect 2596 15104 2648 15113
rect 3516 15104 3568 15156
rect 5448 15147 5500 15156
rect 3240 15036 3292 15088
rect 4068 14968 4120 15020
rect 4252 15011 4304 15020
rect 4252 14977 4261 15011
rect 4261 14977 4295 15011
rect 4295 14977 4304 15011
rect 4252 14968 4304 14977
rect 5448 15113 5457 15147
rect 5457 15113 5491 15147
rect 5491 15113 5500 15147
rect 5448 15104 5500 15113
rect 6000 15104 6052 15156
rect 7012 15104 7064 15156
rect 8116 15104 8168 15156
rect 8300 15147 8352 15156
rect 8300 15113 8309 15147
rect 8309 15113 8343 15147
rect 8343 15113 8352 15147
rect 8300 15104 8352 15113
rect 6920 15079 6972 15088
rect 6920 15045 6929 15079
rect 6929 15045 6963 15079
rect 6963 15045 6972 15079
rect 6920 15036 6972 15045
rect 7472 15036 7524 15088
rect 9128 15036 9180 15088
rect 6184 14968 6236 15020
rect 8024 14968 8076 15020
rect 9956 15104 10008 15156
rect 10324 15147 10376 15156
rect 10324 15113 10333 15147
rect 10333 15113 10367 15147
rect 10367 15113 10376 15147
rect 10324 15104 10376 15113
rect 11888 15104 11940 15156
rect 13268 15104 13320 15156
rect 13728 15104 13780 15156
rect 14004 15147 14056 15156
rect 14004 15113 14013 15147
rect 14013 15113 14047 15147
rect 14047 15113 14056 15147
rect 14004 15104 14056 15113
rect 16120 15104 16172 15156
rect 17224 15147 17276 15156
rect 17224 15113 17233 15147
rect 17233 15113 17267 15147
rect 17267 15113 17276 15147
rect 17224 15104 17276 15113
rect 17408 15104 17460 15156
rect 18236 15147 18288 15156
rect 18236 15113 18245 15147
rect 18245 15113 18279 15147
rect 18279 15113 18288 15147
rect 18236 15104 18288 15113
rect 18420 15104 18472 15156
rect 11152 15036 11204 15088
rect 12440 15036 12492 15088
rect 1676 14900 1728 14952
rect 1952 14900 2004 14952
rect 3240 14943 3292 14952
rect 3240 14909 3249 14943
rect 3249 14909 3283 14943
rect 3283 14909 3292 14943
rect 3240 14900 3292 14909
rect 3332 14900 3384 14952
rect 14648 14900 14700 14952
rect 3424 14875 3476 14884
rect 3424 14841 3433 14875
rect 3433 14841 3467 14875
rect 3467 14841 3476 14875
rect 3424 14832 3476 14841
rect 3608 14832 3660 14884
rect 8392 14832 8444 14884
rect 9956 14832 10008 14884
rect 12532 14832 12584 14884
rect 12900 14875 12952 14884
rect 12900 14841 12909 14875
rect 12909 14841 12943 14875
rect 12943 14841 12952 14875
rect 12900 14832 12952 14841
rect 13084 14875 13136 14884
rect 13084 14841 13093 14875
rect 13093 14841 13127 14875
rect 13127 14841 13136 14875
rect 13084 14832 13136 14841
rect 1492 14764 1544 14816
rect 2596 14764 2648 14816
rect 2780 14764 2832 14816
rect 4252 14764 4304 14816
rect 6736 14764 6788 14816
rect 7380 14807 7432 14816
rect 7380 14773 7389 14807
rect 7389 14773 7423 14807
rect 7423 14773 7432 14807
rect 7380 14764 7432 14773
rect 9036 14807 9088 14816
rect 9036 14773 9045 14807
rect 9045 14773 9079 14807
rect 9079 14773 9088 14807
rect 9036 14764 9088 14773
rect 9404 14764 9456 14816
rect 11060 14764 11112 14816
rect 12440 14764 12492 14816
rect 15568 14832 15620 14884
rect 14556 14764 14608 14816
rect 15660 14764 15712 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2044 14560 2096 14612
rect 2596 14560 2648 14612
rect 2872 14492 2924 14544
rect 3240 14560 3292 14612
rect 3608 14560 3660 14612
rect 4804 14560 4856 14612
rect 6000 14560 6052 14612
rect 6184 14603 6236 14612
rect 6184 14569 6193 14603
rect 6193 14569 6227 14603
rect 6227 14569 6236 14603
rect 6184 14560 6236 14569
rect 8392 14603 8444 14612
rect 8392 14569 8401 14603
rect 8401 14569 8435 14603
rect 8435 14569 8444 14603
rect 8392 14560 8444 14569
rect 9956 14560 10008 14612
rect 10048 14560 10100 14612
rect 12900 14560 12952 14612
rect 15108 14603 15160 14612
rect 3332 14492 3384 14544
rect 4528 14492 4580 14544
rect 5540 14492 5592 14544
rect 7380 14492 7432 14544
rect 3516 14424 3568 14476
rect 5448 14424 5500 14476
rect 7656 14424 7708 14476
rect 9956 14424 10008 14476
rect 15108 14569 15117 14603
rect 15117 14569 15151 14603
rect 15151 14569 15160 14603
rect 15108 14560 15160 14569
rect 15936 14603 15988 14612
rect 15936 14569 15945 14603
rect 15945 14569 15979 14603
rect 15979 14569 15988 14603
rect 15936 14560 15988 14569
rect 17500 14603 17552 14612
rect 17500 14569 17509 14603
rect 17509 14569 17543 14603
rect 17543 14569 17552 14603
rect 17500 14560 17552 14569
rect 15476 14492 15528 14544
rect 16120 14492 16172 14544
rect 14648 14424 14700 14476
rect 16396 14467 16448 14476
rect 16396 14433 16430 14467
rect 16430 14433 16448 14467
rect 16396 14424 16448 14433
rect 3424 14356 3476 14408
rect 10600 14356 10652 14408
rect 13176 14356 13228 14408
rect 14280 14356 14332 14408
rect 15660 14356 15712 14408
rect 11888 14288 11940 14340
rect 1952 14220 2004 14272
rect 2136 14220 2188 14272
rect 4068 14220 4120 14272
rect 5356 14220 5408 14272
rect 9404 14220 9456 14272
rect 11152 14220 11204 14272
rect 12532 14220 12584 14272
rect 13820 14220 13872 14272
rect 14096 14220 14148 14272
rect 14648 14263 14700 14272
rect 14648 14229 14657 14263
rect 14657 14229 14691 14263
rect 14691 14229 14700 14263
rect 14648 14220 14700 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2596 14059 2648 14068
rect 2596 14025 2605 14059
rect 2605 14025 2639 14059
rect 2639 14025 2648 14059
rect 2596 14016 2648 14025
rect 2872 14016 2924 14068
rect 1676 13991 1728 14000
rect 1676 13957 1685 13991
rect 1685 13957 1719 13991
rect 1719 13957 1728 13991
rect 1676 13948 1728 13957
rect 2320 13880 2372 13932
rect 3516 14016 3568 14068
rect 4528 14059 4580 14068
rect 4528 14025 4537 14059
rect 4537 14025 4571 14059
rect 4571 14025 4580 14059
rect 4528 14016 4580 14025
rect 5540 13948 5592 14000
rect 5448 13880 5500 13932
rect 6000 13880 6052 13932
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 10600 14059 10652 14068
rect 10600 14025 10609 14059
rect 10609 14025 10643 14059
rect 10643 14025 10652 14059
rect 10600 14016 10652 14025
rect 14280 14016 14332 14068
rect 14740 14059 14792 14068
rect 14740 14025 14749 14059
rect 14749 14025 14783 14059
rect 14783 14025 14792 14059
rect 14740 14016 14792 14025
rect 10876 13991 10928 14000
rect 10876 13957 10885 13991
rect 10885 13957 10919 13991
rect 10919 13957 10928 13991
rect 10876 13948 10928 13957
rect 14924 13948 14976 14000
rect 15108 13880 15160 13932
rect 15384 13923 15436 13932
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 15384 13880 15436 13889
rect 3240 13812 3292 13864
rect 5080 13812 5132 13864
rect 2228 13787 2280 13796
rect 2228 13753 2237 13787
rect 2237 13753 2271 13787
rect 2271 13753 2280 13787
rect 2228 13744 2280 13753
rect 6736 13744 6788 13796
rect 11152 13855 11204 13864
rect 11152 13821 11161 13855
rect 11161 13821 11195 13855
rect 11195 13821 11204 13855
rect 11152 13812 11204 13821
rect 12348 13744 12400 13796
rect 12532 13744 12584 13796
rect 12808 13744 12860 13796
rect 14648 13744 14700 13796
rect 2136 13719 2188 13728
rect 2136 13685 2145 13719
rect 2145 13685 2179 13719
rect 2179 13685 2188 13719
rect 2136 13676 2188 13685
rect 8208 13719 8260 13728
rect 8208 13685 8217 13719
rect 8217 13685 8251 13719
rect 8251 13685 8260 13719
rect 8208 13676 8260 13685
rect 11336 13719 11388 13728
rect 11336 13685 11345 13719
rect 11345 13685 11379 13719
rect 11379 13685 11388 13719
rect 11336 13676 11388 13685
rect 13728 13676 13780 13728
rect 15016 13744 15068 13796
rect 16396 13812 16448 13864
rect 17040 13812 17092 13864
rect 15660 13676 15712 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2228 13472 2280 13524
rect 3240 13472 3292 13524
rect 3516 13515 3568 13524
rect 3516 13481 3525 13515
rect 3525 13481 3559 13515
rect 3559 13481 3568 13515
rect 3516 13472 3568 13481
rect 6736 13515 6788 13524
rect 6736 13481 6745 13515
rect 6745 13481 6779 13515
rect 6779 13481 6788 13515
rect 6736 13472 6788 13481
rect 7472 13515 7524 13524
rect 7472 13481 7481 13515
rect 7481 13481 7515 13515
rect 7515 13481 7524 13515
rect 7472 13472 7524 13481
rect 9956 13472 10008 13524
rect 10876 13472 10928 13524
rect 11888 13472 11940 13524
rect 15108 13472 15160 13524
rect 17040 13515 17092 13524
rect 17040 13481 17049 13515
rect 17049 13481 17083 13515
rect 17083 13481 17092 13515
rect 17040 13472 17092 13481
rect 2872 13404 2924 13456
rect 3884 13404 3936 13456
rect 4068 13404 4120 13456
rect 4620 13447 4672 13456
rect 4620 13413 4629 13447
rect 4629 13413 4663 13447
rect 4663 13413 4672 13447
rect 4620 13404 4672 13413
rect 6920 13404 6972 13456
rect 12348 13404 12400 13456
rect 13728 13404 13780 13456
rect 14096 13404 14148 13456
rect 15016 13447 15068 13456
rect 15016 13413 15025 13447
rect 15025 13413 15059 13447
rect 15059 13413 15068 13447
rect 15016 13404 15068 13413
rect 16120 13404 16172 13456
rect 2044 13336 2096 13388
rect 4804 13336 4856 13388
rect 6276 13336 6328 13388
rect 11888 13336 11940 13388
rect 12716 13336 12768 13388
rect 18512 13379 18564 13388
rect 18512 13345 18521 13379
rect 18521 13345 18555 13379
rect 18555 13345 18564 13379
rect 18512 13336 18564 13345
rect 8208 13268 8260 13320
rect 4160 13243 4212 13252
rect 4160 13209 4169 13243
rect 4169 13209 4203 13243
rect 4203 13209 4212 13243
rect 4160 13200 4212 13209
rect 11704 13311 11756 13320
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 12532 13268 12584 13320
rect 15660 13311 15712 13320
rect 15660 13277 15669 13311
rect 15669 13277 15703 13311
rect 15703 13277 15712 13311
rect 15660 13268 15712 13277
rect 19432 13268 19484 13320
rect 11336 13200 11388 13252
rect 3056 13132 3108 13184
rect 4068 13132 4120 13184
rect 5080 13175 5132 13184
rect 5080 13141 5089 13175
rect 5089 13141 5123 13175
rect 5123 13141 5132 13175
rect 5080 13132 5132 13141
rect 6092 13132 6144 13184
rect 7012 13175 7064 13184
rect 7012 13141 7021 13175
rect 7021 13141 7055 13175
rect 7055 13141 7064 13175
rect 7012 13132 7064 13141
rect 7564 13132 7616 13184
rect 8484 13132 8536 13184
rect 10324 13175 10376 13184
rect 10324 13141 10333 13175
rect 10333 13141 10367 13175
rect 10367 13141 10376 13175
rect 10324 13132 10376 13141
rect 11060 13132 11112 13184
rect 11428 13132 11480 13184
rect 11520 13132 11572 13184
rect 15476 13175 15528 13184
rect 15476 13141 15485 13175
rect 15485 13141 15519 13175
rect 15519 13141 15528 13175
rect 15476 13132 15528 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2044 12971 2096 12980
rect 2044 12937 2053 12971
rect 2053 12937 2087 12971
rect 2087 12937 2096 12971
rect 2044 12928 2096 12937
rect 2320 12928 2372 12980
rect 2780 12928 2832 12980
rect 3884 12971 3936 12980
rect 1676 12860 1728 12912
rect 2872 12860 2924 12912
rect 3884 12937 3893 12971
rect 3893 12937 3927 12971
rect 3927 12937 3936 12971
rect 3884 12928 3936 12937
rect 4620 12928 4672 12980
rect 4804 12928 4856 12980
rect 6276 12928 6328 12980
rect 8208 12971 8260 12980
rect 8208 12937 8217 12971
rect 8217 12937 8251 12971
rect 8251 12937 8260 12971
rect 8208 12928 8260 12937
rect 10324 12928 10376 12980
rect 10784 12971 10836 12980
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 12900 12971 12952 12980
rect 12900 12937 12909 12971
rect 12909 12937 12943 12971
rect 12943 12937 12952 12971
rect 12900 12928 12952 12937
rect 14096 12971 14148 12980
rect 14096 12937 14105 12971
rect 14105 12937 14139 12971
rect 14139 12937 14148 12971
rect 14096 12928 14148 12937
rect 14648 12928 14700 12980
rect 16120 12971 16172 12980
rect 16120 12937 16129 12971
rect 16129 12937 16163 12971
rect 16163 12937 16172 12971
rect 16120 12928 16172 12937
rect 18512 12971 18564 12980
rect 18512 12937 18521 12971
rect 18521 12937 18555 12971
rect 18555 12937 18564 12971
rect 18512 12928 18564 12937
rect 5356 12860 5408 12912
rect 6920 12903 6972 12912
rect 6920 12869 6929 12903
rect 6929 12869 6963 12903
rect 6963 12869 6972 12903
rect 6920 12860 6972 12869
rect 10876 12860 10928 12912
rect 12716 12860 12768 12912
rect 13084 12860 13136 12912
rect 4344 12792 4396 12844
rect 5080 12792 5132 12844
rect 1308 12724 1360 12776
rect 1768 12724 1820 12776
rect 3884 12724 3936 12776
rect 4436 12724 4488 12776
rect 6460 12792 6512 12844
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 9956 12792 10008 12844
rect 11060 12792 11112 12844
rect 11428 12792 11480 12844
rect 6552 12724 6604 12776
rect 3976 12656 4028 12708
rect 4068 12656 4120 12708
rect 4528 12656 4580 12708
rect 12900 12724 12952 12776
rect 8116 12656 8168 12708
rect 9404 12656 9456 12708
rect 11060 12699 11112 12708
rect 11060 12665 11069 12699
rect 11069 12665 11103 12699
rect 11103 12665 11112 12699
rect 11060 12656 11112 12665
rect 16120 12724 16172 12776
rect 14004 12656 14056 12708
rect 1768 12588 1820 12640
rect 3056 12631 3108 12640
rect 3056 12597 3065 12631
rect 3065 12597 3099 12631
rect 3099 12597 3108 12631
rect 3056 12588 3108 12597
rect 4896 12588 4948 12640
rect 8024 12588 8076 12640
rect 9036 12588 9088 12640
rect 9956 12588 10008 12640
rect 11244 12631 11296 12640
rect 11244 12597 11253 12631
rect 11253 12597 11287 12631
rect 11287 12597 11296 12631
rect 11244 12588 11296 12597
rect 15476 12588 15528 12640
rect 15660 12588 15712 12640
rect 16488 12588 16540 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1400 12384 1452 12436
rect 3056 12384 3108 12436
rect 3884 12427 3936 12436
rect 3884 12393 3893 12427
rect 3893 12393 3927 12427
rect 3927 12393 3936 12427
rect 3884 12384 3936 12393
rect 5448 12384 5500 12436
rect 6920 12384 6972 12436
rect 7472 12384 7524 12436
rect 11704 12384 11756 12436
rect 12440 12384 12492 12436
rect 12808 12384 12860 12436
rect 14188 12427 14240 12436
rect 14188 12393 14197 12427
rect 14197 12393 14231 12427
rect 14231 12393 14240 12427
rect 14188 12384 14240 12393
rect 1952 12316 2004 12368
rect 2964 12359 3016 12368
rect 2964 12325 2973 12359
rect 2973 12325 3007 12359
rect 3007 12325 3016 12359
rect 2964 12316 3016 12325
rect 4436 12316 4488 12368
rect 2228 12248 2280 12300
rect 3240 12248 3292 12300
rect 6000 12316 6052 12368
rect 7104 12316 7156 12368
rect 7932 12316 7984 12368
rect 9036 12316 9088 12368
rect 11428 12316 11480 12368
rect 11796 12359 11848 12368
rect 11796 12325 11805 12359
rect 11805 12325 11839 12359
rect 11839 12325 11848 12359
rect 11796 12316 11848 12325
rect 13360 12359 13412 12368
rect 13360 12325 13369 12359
rect 13369 12325 13403 12359
rect 13403 12325 13412 12359
rect 13360 12316 13412 12325
rect 13820 12316 13872 12368
rect 14832 12316 14884 12368
rect 2964 12180 3016 12232
rect 4804 12180 4856 12232
rect 6368 12248 6420 12300
rect 8116 12248 8168 12300
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 10692 12291 10744 12300
rect 10692 12257 10701 12291
rect 10701 12257 10735 12291
rect 10735 12257 10744 12291
rect 10692 12248 10744 12257
rect 11060 12248 11112 12300
rect 13176 12291 13228 12300
rect 13176 12257 13185 12291
rect 13185 12257 13219 12291
rect 13219 12257 13228 12291
rect 13176 12248 13228 12257
rect 14004 12248 14056 12300
rect 15568 12248 15620 12300
rect 16764 12248 16816 12300
rect 19432 12248 19484 12300
rect 8668 12180 8720 12232
rect 9128 12180 9180 12232
rect 9588 12180 9640 12232
rect 2780 12112 2832 12164
rect 4344 12155 4396 12164
rect 4344 12121 4353 12155
rect 4353 12121 4387 12155
rect 4387 12121 4396 12155
rect 4344 12112 4396 12121
rect 8300 12112 8352 12164
rect 9220 12112 9272 12164
rect 10784 12112 10836 12164
rect 13268 12180 13320 12232
rect 13452 12223 13504 12232
rect 13452 12189 13461 12223
rect 13461 12189 13495 12223
rect 13495 12189 13504 12223
rect 13452 12180 13504 12189
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 12900 12155 12952 12164
rect 12900 12121 12909 12155
rect 12909 12121 12943 12155
rect 12943 12121 12952 12155
rect 12900 12112 12952 12121
rect 13360 12112 13412 12164
rect 15016 12112 15068 12164
rect 15476 12112 15528 12164
rect 2044 12044 2096 12096
rect 2872 12044 2924 12096
rect 3148 12044 3200 12096
rect 6920 12044 6972 12096
rect 8024 12044 8076 12096
rect 8576 12044 8628 12096
rect 9404 12044 9456 12096
rect 9588 12044 9640 12096
rect 11152 12044 11204 12096
rect 12624 12044 12676 12096
rect 12992 12044 13044 12096
rect 14832 12044 14884 12096
rect 15292 12044 15344 12096
rect 20628 12044 20680 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1952 11883 2004 11892
rect 1952 11849 1961 11883
rect 1961 11849 1995 11883
rect 1995 11849 2004 11883
rect 1952 11840 2004 11849
rect 4528 11840 4580 11892
rect 6000 11840 6052 11892
rect 4804 11815 4856 11824
rect 4804 11781 4813 11815
rect 4813 11781 4847 11815
rect 4847 11781 4856 11815
rect 4804 11772 4856 11781
rect 8116 11840 8168 11892
rect 9496 11840 9548 11892
rect 10048 11840 10100 11892
rect 10692 11840 10744 11892
rect 11796 11840 11848 11892
rect 13452 11883 13504 11892
rect 13452 11849 13461 11883
rect 13461 11849 13495 11883
rect 13495 11849 13504 11883
rect 13452 11840 13504 11849
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 15752 11840 15804 11892
rect 16764 11883 16816 11892
rect 16764 11849 16773 11883
rect 16773 11849 16807 11883
rect 16807 11849 16816 11883
rect 16764 11840 16816 11849
rect 19432 11840 19484 11892
rect 9036 11772 9088 11824
rect 9680 11815 9732 11824
rect 9680 11781 9689 11815
rect 9689 11781 9723 11815
rect 9723 11781 9732 11815
rect 9680 11772 9732 11781
rect 12532 11815 12584 11824
rect 12532 11781 12541 11815
rect 12541 11781 12575 11815
rect 12575 11781 12584 11815
rect 12532 11772 12584 11781
rect 10048 11704 10100 11756
rect 11244 11704 11296 11756
rect 3424 11636 3476 11688
rect 3608 11636 3660 11688
rect 3792 11636 3844 11688
rect 5172 11636 5224 11688
rect 6920 11636 6972 11688
rect 8208 11636 8260 11688
rect 2228 11568 2280 11620
rect 5540 11611 5592 11620
rect 5540 11577 5549 11611
rect 5549 11577 5583 11611
rect 5583 11577 5592 11611
rect 5540 11568 5592 11577
rect 10140 11611 10192 11620
rect 10140 11577 10149 11611
rect 10149 11577 10183 11611
rect 10183 11577 10192 11611
rect 10140 11568 10192 11577
rect 14188 11636 14240 11688
rect 15200 11636 15252 11688
rect 12992 11611 13044 11620
rect 12992 11577 13001 11611
rect 13001 11577 13035 11611
rect 13035 11577 13044 11611
rect 12992 11568 13044 11577
rect 13268 11568 13320 11620
rect 14280 11611 14332 11620
rect 14280 11577 14289 11611
rect 14289 11577 14323 11611
rect 14323 11577 14332 11611
rect 14280 11568 14332 11577
rect 15292 11568 15344 11620
rect 1400 11543 1452 11552
rect 1400 11509 1409 11543
rect 1409 11509 1443 11543
rect 1443 11509 1452 11543
rect 1400 11500 1452 11509
rect 3056 11500 3108 11552
rect 3792 11543 3844 11552
rect 3792 11509 3801 11543
rect 3801 11509 3835 11543
rect 3835 11509 3844 11543
rect 3792 11500 3844 11509
rect 4344 11543 4396 11552
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 5448 11500 5500 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2228 11296 2280 11348
rect 2780 11339 2832 11348
rect 2780 11305 2789 11339
rect 2789 11305 2823 11339
rect 2823 11305 2832 11339
rect 2780 11296 2832 11305
rect 3516 11296 3568 11348
rect 5540 11339 5592 11348
rect 5540 11305 5549 11339
rect 5549 11305 5583 11339
rect 5583 11305 5592 11339
rect 5540 11296 5592 11305
rect 6460 11296 6512 11348
rect 8208 11296 8260 11348
rect 9220 11296 9272 11348
rect 10140 11296 10192 11348
rect 10784 11296 10836 11348
rect 13176 11296 13228 11348
rect 15292 11296 15344 11348
rect 1400 11228 1452 11280
rect 2504 11228 2556 11280
rect 3332 11228 3384 11280
rect 3792 11228 3844 11280
rect 4620 11228 4672 11280
rect 4804 11271 4856 11280
rect 4804 11237 4813 11271
rect 4813 11237 4847 11271
rect 4847 11237 4856 11271
rect 4804 11228 4856 11237
rect 6368 11271 6420 11280
rect 6368 11237 6377 11271
rect 6377 11237 6411 11271
rect 6411 11237 6420 11271
rect 6368 11228 6420 11237
rect 9036 11228 9088 11280
rect 9680 11228 9732 11280
rect 2228 11160 2280 11212
rect 3148 11160 3200 11212
rect 3240 11160 3292 11212
rect 5172 11203 5224 11212
rect 5172 11169 5181 11203
rect 5181 11169 5215 11203
rect 5215 11169 5224 11203
rect 5172 11160 5224 11169
rect 5448 11160 5500 11212
rect 9588 11160 9640 11212
rect 15660 11228 15712 11280
rect 3424 11092 3476 11144
rect 1952 10956 2004 11008
rect 5080 11024 5132 11076
rect 5356 11024 5408 11076
rect 6920 11024 6972 11076
rect 8576 11092 8628 11144
rect 11060 11160 11112 11212
rect 11336 11160 11388 11212
rect 13728 11203 13780 11212
rect 13728 11169 13737 11203
rect 13737 11169 13771 11203
rect 13771 11169 13780 11203
rect 13728 11160 13780 11169
rect 14648 11160 14700 11212
rect 10784 11092 10836 11144
rect 11244 11135 11296 11144
rect 11244 11101 11253 11135
rect 11253 11101 11287 11135
rect 11287 11101 11296 11135
rect 11244 11092 11296 11101
rect 14004 11135 14056 11144
rect 14004 11101 14013 11135
rect 14013 11101 14047 11135
rect 14047 11101 14056 11135
rect 14004 11092 14056 11101
rect 15200 11092 15252 11144
rect 9772 11067 9824 11076
rect 9772 11033 9781 11067
rect 9781 11033 9815 11067
rect 9815 11033 9824 11067
rect 9772 11024 9824 11033
rect 13268 11067 13320 11076
rect 13268 11033 13277 11067
rect 13277 11033 13311 11067
rect 13311 11033 13320 11067
rect 13268 11024 13320 11033
rect 2872 10956 2924 11008
rect 4620 10956 4672 11008
rect 6000 10956 6052 11008
rect 7380 10999 7432 11008
rect 7380 10965 7389 10999
rect 7389 10965 7423 10999
rect 7423 10965 7432 10999
rect 7380 10956 7432 10965
rect 8760 10956 8812 11008
rect 10048 10956 10100 11008
rect 12624 10999 12676 11008
rect 12624 10965 12633 10999
rect 12633 10965 12667 10999
rect 12667 10965 12676 10999
rect 12624 10956 12676 10965
rect 16488 10956 16540 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2504 10795 2556 10804
rect 2504 10761 2513 10795
rect 2513 10761 2547 10795
rect 2547 10761 2556 10795
rect 2504 10752 2556 10761
rect 2964 10684 3016 10736
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 3424 10752 3476 10804
rect 5448 10795 5500 10804
rect 5448 10761 5457 10795
rect 5457 10761 5491 10795
rect 5491 10761 5500 10795
rect 5448 10752 5500 10761
rect 6460 10752 6512 10804
rect 8944 10752 8996 10804
rect 10048 10752 10100 10804
rect 11336 10752 11388 10804
rect 13176 10752 13228 10804
rect 14648 10752 14700 10804
rect 14832 10752 14884 10804
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 8300 10684 8352 10736
rect 7656 10616 7708 10625
rect 2228 10548 2280 10600
rect 3332 10591 3384 10600
rect 3332 10557 3366 10591
rect 3366 10557 3384 10591
rect 3332 10548 3384 10557
rect 1952 10480 2004 10532
rect 5356 10548 5408 10600
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 7288 10548 7340 10600
rect 8300 10548 8352 10600
rect 15292 10616 15344 10668
rect 12624 10548 12676 10600
rect 16580 10591 16632 10600
rect 16580 10557 16589 10591
rect 16589 10557 16623 10591
rect 16623 10557 16632 10591
rect 16580 10548 16632 10557
rect 11244 10480 11296 10532
rect 2136 10412 2188 10464
rect 3424 10412 3476 10464
rect 4528 10412 4580 10464
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 5080 10412 5132 10421
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 6920 10412 6972 10464
rect 8300 10412 8352 10464
rect 10784 10412 10836 10464
rect 11428 10412 11480 10464
rect 13544 10480 13596 10532
rect 15660 10480 15712 10532
rect 16856 10523 16908 10532
rect 16856 10489 16865 10523
rect 16865 10489 16899 10523
rect 16899 10489 16908 10523
rect 16856 10480 16908 10489
rect 13636 10412 13688 10464
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 16488 10412 16540 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2228 10251 2280 10260
rect 2228 10217 2237 10251
rect 2237 10217 2271 10251
rect 2271 10217 2280 10251
rect 2228 10208 2280 10217
rect 2412 10208 2464 10260
rect 2688 10208 2740 10260
rect 3332 10208 3384 10260
rect 3516 10208 3568 10260
rect 4620 10251 4672 10260
rect 4620 10217 4629 10251
rect 4629 10217 4663 10251
rect 4663 10217 4672 10251
rect 4620 10208 4672 10217
rect 4804 10208 4856 10260
rect 7472 10208 7524 10260
rect 7656 10208 7708 10260
rect 9036 10251 9088 10260
rect 9036 10217 9045 10251
rect 9045 10217 9079 10251
rect 9079 10217 9088 10251
rect 9036 10208 9088 10217
rect 9588 10208 9640 10260
rect 9680 10208 9732 10260
rect 11060 10208 11112 10260
rect 13728 10208 13780 10260
rect 2964 10183 3016 10192
rect 2964 10149 2973 10183
rect 2973 10149 3007 10183
rect 3007 10149 3016 10183
rect 2964 10140 3016 10149
rect 5540 10140 5592 10192
rect 10692 10183 10744 10192
rect 2688 10072 2740 10124
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 4528 10004 4580 10056
rect 5632 9936 5684 9988
rect 6092 10004 6144 10056
rect 6644 10072 6696 10124
rect 10692 10149 10701 10183
rect 10701 10149 10735 10183
rect 10735 10149 10744 10183
rect 10692 10140 10744 10149
rect 12440 10140 12492 10192
rect 13176 10183 13228 10192
rect 13176 10149 13185 10183
rect 13185 10149 13219 10183
rect 13219 10149 13228 10183
rect 13176 10140 13228 10149
rect 15476 10140 15528 10192
rect 16120 10140 16172 10192
rect 10508 10115 10560 10124
rect 6828 9936 6880 9988
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 12716 10072 12768 10124
rect 14280 10072 14332 10124
rect 14648 10072 14700 10124
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 8760 10004 8812 10056
rect 9036 10004 9088 10056
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 12624 10004 12676 10056
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 14188 9936 14240 9988
rect 15384 9979 15436 9988
rect 3884 9868 3936 9920
rect 5264 9911 5316 9920
rect 5264 9877 5273 9911
rect 5273 9877 5307 9911
rect 5307 9877 5316 9911
rect 5264 9868 5316 9877
rect 8760 9868 8812 9920
rect 11060 9868 11112 9920
rect 11888 9911 11940 9920
rect 11888 9877 11897 9911
rect 11897 9877 11931 9911
rect 11931 9877 11940 9911
rect 11888 9868 11940 9877
rect 13912 9911 13964 9920
rect 13912 9877 13921 9911
rect 13921 9877 13955 9911
rect 13955 9877 13964 9911
rect 13912 9868 13964 9877
rect 14280 9911 14332 9920
rect 14280 9877 14289 9911
rect 14289 9877 14323 9911
rect 14323 9877 14332 9911
rect 14280 9868 14332 9877
rect 15384 9945 15393 9979
rect 15393 9945 15427 9979
rect 15427 9945 15436 9979
rect 15384 9936 15436 9945
rect 15568 9868 15620 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2964 9664 3016 9716
rect 9036 9707 9088 9716
rect 9036 9673 9045 9707
rect 9045 9673 9079 9707
rect 9079 9673 9088 9707
rect 9036 9664 9088 9673
rect 10508 9664 10560 9716
rect 10784 9664 10836 9716
rect 2688 9596 2740 9648
rect 6276 9596 6328 9648
rect 6828 9596 6880 9648
rect 11060 9596 11112 9648
rect 11796 9639 11848 9648
rect 11796 9605 11805 9639
rect 11805 9605 11839 9639
rect 11839 9605 11848 9639
rect 11796 9596 11848 9605
rect 2596 9528 2648 9580
rect 8760 9528 8812 9580
rect 1584 9503 1636 9512
rect 1584 9469 1593 9503
rect 1593 9469 1627 9503
rect 1627 9469 1636 9503
rect 1584 9460 1636 9469
rect 1860 9435 1912 9444
rect 1860 9401 1869 9435
rect 1869 9401 1903 9435
rect 1903 9401 1912 9435
rect 1860 9392 1912 9401
rect 4160 9460 4212 9512
rect 4528 9503 4580 9512
rect 4528 9469 4562 9503
rect 4562 9469 4580 9503
rect 4528 9460 4580 9469
rect 8392 9503 8444 9512
rect 3700 9392 3752 9444
rect 4344 9392 4396 9444
rect 2780 9324 2832 9376
rect 3240 9324 3292 9376
rect 4160 9367 4212 9376
rect 4160 9333 4169 9367
rect 4169 9333 4203 9367
rect 4203 9333 4212 9367
rect 4160 9324 4212 9333
rect 4896 9324 4948 9376
rect 6920 9392 6972 9444
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 9496 9528 9548 9580
rect 11152 9528 11204 9580
rect 13176 9664 13228 9716
rect 15476 9664 15528 9716
rect 16856 9707 16908 9716
rect 16856 9673 16865 9707
rect 16865 9673 16899 9707
rect 16899 9673 16908 9707
rect 16856 9664 16908 9673
rect 12900 9639 12952 9648
rect 12900 9605 12909 9639
rect 12909 9605 12943 9639
rect 12943 9605 12952 9639
rect 12900 9596 12952 9605
rect 13360 9639 13412 9648
rect 13360 9605 13369 9639
rect 13369 9605 13403 9639
rect 13403 9605 13412 9639
rect 13360 9596 13412 9605
rect 13636 9460 13688 9512
rect 13912 9460 13964 9512
rect 14372 9460 14424 9512
rect 14464 9460 14516 9512
rect 7564 9392 7616 9444
rect 10876 9392 10928 9444
rect 18052 9528 18104 9580
rect 16856 9460 16908 9512
rect 16120 9435 16172 9444
rect 16120 9401 16129 9435
rect 16129 9401 16163 9435
rect 16163 9401 16172 9435
rect 16120 9392 16172 9401
rect 8392 9324 8444 9376
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 11152 9367 11204 9376
rect 11152 9333 11161 9367
rect 11161 9333 11195 9367
rect 11195 9333 11204 9367
rect 11152 9324 11204 9333
rect 11244 9324 11296 9376
rect 13636 9367 13688 9376
rect 13636 9333 13645 9367
rect 13645 9333 13679 9367
rect 13679 9333 13688 9367
rect 13636 9324 13688 9333
rect 15200 9367 15252 9376
rect 15200 9333 15209 9367
rect 15209 9333 15243 9367
rect 15243 9333 15252 9367
rect 15200 9324 15252 9333
rect 17500 9324 17552 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2044 9120 2096 9172
rect 2872 9120 2924 9172
rect 4528 9120 4580 9172
rect 8300 9120 8352 9172
rect 8576 9120 8628 9172
rect 9496 9163 9548 9172
rect 9496 9129 9505 9163
rect 9505 9129 9539 9163
rect 9539 9129 9548 9163
rect 9496 9120 9548 9129
rect 9864 9163 9916 9172
rect 9864 9129 9873 9163
rect 9873 9129 9907 9163
rect 9907 9129 9916 9163
rect 9864 9120 9916 9129
rect 10692 9163 10744 9172
rect 10692 9129 10701 9163
rect 10701 9129 10735 9163
rect 10735 9129 10744 9163
rect 10692 9120 10744 9129
rect 12440 9163 12492 9172
rect 12440 9129 12449 9163
rect 12449 9129 12483 9163
rect 12483 9129 12492 9163
rect 12440 9120 12492 9129
rect 12716 9120 12768 9172
rect 14648 9163 14700 9172
rect 14648 9129 14657 9163
rect 14657 9129 14691 9163
rect 14691 9129 14700 9163
rect 14648 9120 14700 9129
rect 15936 9163 15988 9172
rect 15936 9129 15945 9163
rect 15945 9129 15979 9163
rect 15979 9129 15988 9163
rect 15936 9120 15988 9129
rect 2780 9052 2832 9104
rect 3976 9052 4028 9104
rect 4160 9052 4212 9104
rect 5264 9052 5316 9104
rect 6368 9052 6420 9104
rect 6736 9052 6788 9104
rect 3056 9027 3108 9036
rect 3056 8993 3065 9027
rect 3065 8993 3099 9027
rect 3099 8993 3108 9027
rect 3056 8984 3108 8993
rect 3516 9027 3568 9036
rect 3516 8993 3525 9027
rect 3525 8993 3559 9027
rect 3559 8993 3568 9027
rect 3516 8984 3568 8993
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 5264 8959 5316 8968
rect 5264 8925 5273 8959
rect 5273 8925 5307 8959
rect 5307 8925 5316 8959
rect 5264 8916 5316 8925
rect 5448 8916 5500 8968
rect 5172 8848 5224 8900
rect 2688 8780 2740 8832
rect 5356 8780 5408 8832
rect 6092 8780 6144 8832
rect 6828 8984 6880 9036
rect 13544 9052 13596 9104
rect 13820 9052 13872 9104
rect 7564 8984 7616 9036
rect 8944 8984 8996 9036
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 10048 8984 10100 9036
rect 11336 9027 11388 9036
rect 11336 8993 11370 9027
rect 11370 8993 11388 9027
rect 11336 8984 11388 8993
rect 12348 8984 12400 9036
rect 15384 8984 15436 9036
rect 16396 9027 16448 9036
rect 16396 8993 16405 9027
rect 16405 8993 16439 9027
rect 16439 8993 16448 9027
rect 16396 8984 16448 8993
rect 11060 8959 11112 8968
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 14188 8959 14240 8968
rect 14188 8925 14197 8959
rect 14197 8925 14231 8959
rect 14231 8925 14240 8959
rect 14188 8916 14240 8925
rect 14648 8916 14700 8968
rect 6736 8780 6788 8832
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 8116 8780 8168 8832
rect 10508 8780 10560 8832
rect 13636 8780 13688 8832
rect 15292 8780 15344 8832
rect 16304 8780 16356 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1860 8440 1912 8492
rect 2872 8576 2924 8628
rect 3700 8619 3752 8628
rect 3700 8585 3709 8619
rect 3709 8585 3743 8619
rect 3743 8585 3752 8619
rect 3700 8576 3752 8585
rect 3976 8576 4028 8628
rect 6644 8619 6696 8628
rect 3516 8551 3568 8560
rect 3516 8517 3525 8551
rect 3525 8517 3559 8551
rect 3559 8517 3568 8551
rect 3516 8508 3568 8517
rect 5540 8508 5592 8560
rect 6644 8585 6653 8619
rect 6653 8585 6687 8619
rect 6687 8585 6696 8619
rect 6644 8576 6696 8585
rect 7564 8576 7616 8628
rect 8208 8576 8260 8628
rect 8576 8576 8628 8628
rect 10876 8576 10928 8628
rect 11060 8619 11112 8628
rect 11060 8585 11069 8619
rect 11069 8585 11103 8619
rect 11103 8585 11112 8619
rect 11060 8576 11112 8585
rect 11336 8576 11388 8628
rect 11704 8576 11756 8628
rect 8300 8508 8352 8560
rect 9680 8508 9732 8560
rect 3056 8440 3108 8492
rect 6092 8440 6144 8492
rect 7104 8440 7156 8492
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 8484 8440 8536 8492
rect 8852 8440 8904 8492
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 10324 8483 10376 8492
rect 9312 8440 9364 8449
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 13912 8576 13964 8628
rect 12440 8508 12492 8560
rect 13728 8508 13780 8560
rect 15384 8576 15436 8628
rect 16396 8576 16448 8628
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 1952 8372 2004 8424
rect 2780 8372 2832 8424
rect 3148 8372 3200 8424
rect 3240 8372 3292 8424
rect 3700 8372 3752 8424
rect 4896 8372 4948 8424
rect 7012 8415 7064 8424
rect 7012 8381 7021 8415
rect 7021 8381 7055 8415
rect 7055 8381 7064 8415
rect 7012 8372 7064 8381
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 4528 8347 4580 8356
rect 3424 8236 3476 8288
rect 4528 8313 4562 8347
rect 4562 8313 4580 8347
rect 4528 8304 4580 8313
rect 9496 8372 9548 8424
rect 8944 8347 8996 8356
rect 8944 8313 8953 8347
rect 8953 8313 8987 8347
rect 8987 8313 8996 8347
rect 12072 8372 12124 8424
rect 12900 8372 12952 8424
rect 16120 8372 16172 8424
rect 8944 8304 8996 8313
rect 13544 8304 13596 8356
rect 14648 8304 14700 8356
rect 16488 8304 16540 8356
rect 9864 8236 9916 8288
rect 10968 8236 11020 8288
rect 13452 8236 13504 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2320 8075 2372 8084
rect 2320 8041 2329 8075
rect 2329 8041 2363 8075
rect 2363 8041 2372 8075
rect 2320 8032 2372 8041
rect 3056 8032 3108 8084
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 4160 8032 4212 8084
rect 4528 8032 4580 8084
rect 5264 8032 5316 8084
rect 8668 8032 8720 8084
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 10048 8032 10100 8084
rect 11152 8032 11204 8084
rect 12348 8032 12400 8084
rect 14188 8075 14240 8084
rect 14188 8041 14197 8075
rect 14197 8041 14231 8075
rect 14231 8041 14240 8075
rect 14188 8032 14240 8041
rect 3240 7964 3292 8016
rect 3608 7964 3660 8016
rect 8300 7964 8352 8016
rect 9588 7964 9640 8016
rect 11428 8007 11480 8016
rect 11428 7973 11437 8007
rect 11437 7973 11471 8007
rect 11471 7973 11480 8007
rect 11428 7964 11480 7973
rect 11612 8007 11664 8016
rect 11612 7973 11621 8007
rect 11621 7973 11655 8007
rect 11655 7973 11664 8007
rect 11612 7964 11664 7973
rect 11704 8007 11756 8016
rect 11704 7973 11713 8007
rect 11713 7973 11747 8007
rect 11747 7973 11756 8007
rect 11704 7964 11756 7973
rect 13728 8007 13780 8016
rect 13728 7973 13737 8007
rect 13737 7973 13771 8007
rect 13771 7973 13780 8007
rect 13728 7964 13780 7973
rect 13912 7964 13964 8016
rect 14648 8007 14700 8016
rect 14648 7973 14657 8007
rect 14657 7973 14691 8007
rect 14691 7973 14700 8007
rect 14648 7964 14700 7973
rect 4620 7896 4672 7948
rect 5172 7939 5224 7948
rect 5172 7905 5195 7939
rect 5195 7905 5224 7939
rect 5172 7896 5224 7905
rect 8208 7896 8260 7948
rect 9772 7896 9824 7948
rect 12992 7896 13044 7948
rect 15384 7896 15436 7948
rect 16120 7896 16172 7948
rect 16396 7896 16448 7948
rect 16580 7939 16632 7948
rect 16580 7905 16614 7939
rect 16614 7905 16632 7939
rect 16580 7896 16632 7905
rect 2964 7871 3016 7880
rect 2964 7837 2973 7871
rect 2973 7837 3007 7871
rect 3007 7837 3016 7871
rect 2964 7828 3016 7837
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 4896 7871 4948 7880
rect 3056 7828 3108 7837
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 10048 7828 10100 7880
rect 13636 7871 13688 7880
rect 13636 7837 13645 7871
rect 13645 7837 13679 7871
rect 13679 7837 13688 7871
rect 13636 7828 13688 7837
rect 14924 7871 14976 7880
rect 14924 7837 14933 7871
rect 14933 7837 14967 7871
rect 14967 7837 14976 7871
rect 14924 7828 14976 7837
rect 6736 7760 6788 7812
rect 13452 7760 13504 7812
rect 2136 7692 2188 7744
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 5264 7692 5316 7744
rect 7012 7692 7064 7744
rect 7472 7692 7524 7744
rect 9312 7735 9364 7744
rect 9312 7701 9321 7735
rect 9321 7701 9355 7735
rect 9355 7701 9364 7735
rect 9312 7692 9364 7701
rect 11244 7692 11296 7744
rect 13268 7735 13320 7744
rect 13268 7701 13277 7735
rect 13277 7701 13311 7735
rect 13311 7701 13320 7735
rect 13268 7692 13320 7701
rect 15844 7735 15896 7744
rect 15844 7701 15853 7735
rect 15853 7701 15887 7735
rect 15887 7701 15896 7735
rect 15844 7692 15896 7701
rect 16120 7735 16172 7744
rect 16120 7701 16129 7735
rect 16129 7701 16163 7735
rect 16163 7701 16172 7735
rect 16120 7692 16172 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2964 7488 3016 7540
rect 4620 7488 4672 7540
rect 4712 7488 4764 7540
rect 5448 7488 5500 7540
rect 6276 7488 6328 7540
rect 6828 7488 6880 7540
rect 7104 7488 7156 7540
rect 8116 7488 8168 7540
rect 8300 7531 8352 7540
rect 8300 7497 8309 7531
rect 8309 7497 8343 7531
rect 8343 7497 8352 7531
rect 8300 7488 8352 7497
rect 11428 7488 11480 7540
rect 11704 7488 11756 7540
rect 13728 7488 13780 7540
rect 17592 7531 17644 7540
rect 17592 7497 17601 7531
rect 17601 7497 17635 7531
rect 17635 7497 17644 7531
rect 17592 7488 17644 7497
rect 3332 7463 3384 7472
rect 3332 7429 3341 7463
rect 3341 7429 3375 7463
rect 3375 7429 3384 7463
rect 3332 7420 3384 7429
rect 4068 7352 4120 7404
rect 6184 7420 6236 7472
rect 6460 7420 6512 7472
rect 7564 7420 7616 7472
rect 9588 7420 9640 7472
rect 10784 7463 10836 7472
rect 10784 7429 10793 7463
rect 10793 7429 10827 7463
rect 10827 7429 10836 7463
rect 10784 7420 10836 7429
rect 11612 7420 11664 7472
rect 13912 7420 13964 7472
rect 15568 7463 15620 7472
rect 15568 7429 15577 7463
rect 15577 7429 15611 7463
rect 15611 7429 15620 7463
rect 15568 7420 15620 7429
rect 6092 7352 6144 7404
rect 6644 7352 6696 7404
rect 7472 7395 7524 7404
rect 7472 7361 7481 7395
rect 7481 7361 7515 7395
rect 7515 7361 7524 7395
rect 7472 7352 7524 7361
rect 11244 7395 11296 7404
rect 11244 7361 11253 7395
rect 11253 7361 11287 7395
rect 11287 7361 11296 7395
rect 11244 7352 11296 7361
rect 2320 7327 2372 7336
rect 2320 7293 2329 7327
rect 2329 7293 2363 7327
rect 2363 7293 2372 7327
rect 2320 7284 2372 7293
rect 3976 7284 4028 7336
rect 4896 7284 4948 7336
rect 6184 7284 6236 7336
rect 7012 7284 7064 7336
rect 2044 7259 2096 7268
rect 2044 7225 2053 7259
rect 2053 7225 2087 7259
rect 2087 7225 2096 7259
rect 2044 7216 2096 7225
rect 2136 7216 2188 7268
rect 7104 7216 7156 7268
rect 9496 7259 9548 7268
rect 9496 7225 9505 7259
rect 9505 7225 9539 7259
rect 9539 7225 9548 7259
rect 9496 7216 9548 7225
rect 12256 7352 12308 7404
rect 12532 7352 12584 7404
rect 12348 7284 12400 7336
rect 13268 7284 13320 7336
rect 14464 7352 14516 7404
rect 14648 7352 14700 7404
rect 16120 7352 16172 7404
rect 10692 7216 10744 7268
rect 11152 7216 11204 7268
rect 19064 7284 19116 7336
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 2780 7148 2832 7157
rect 4068 7148 4120 7200
rect 4712 7148 4764 7200
rect 6276 7148 6328 7200
rect 7932 7148 7984 7200
rect 9864 7148 9916 7200
rect 13176 7148 13228 7200
rect 14832 7148 14884 7200
rect 15844 7216 15896 7268
rect 16580 7216 16632 7268
rect 18052 7259 18104 7268
rect 18052 7225 18061 7259
rect 18061 7225 18095 7259
rect 18095 7225 18104 7259
rect 18052 7216 18104 7225
rect 16396 7148 16448 7200
rect 16764 7148 16816 7200
rect 16948 7191 17000 7200
rect 16948 7157 16957 7191
rect 16957 7157 16991 7191
rect 16991 7157 17000 7191
rect 16948 7148 17000 7157
rect 17224 7191 17276 7200
rect 17224 7157 17233 7191
rect 17233 7157 17267 7191
rect 17267 7157 17276 7191
rect 17224 7148 17276 7157
rect 18512 7191 18564 7200
rect 18512 7157 18521 7191
rect 18521 7157 18555 7191
rect 18555 7157 18564 7191
rect 18512 7148 18564 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 2872 6944 2924 6996
rect 3608 6944 3660 6996
rect 3976 6944 4028 6996
rect 6092 6987 6144 6996
rect 3240 6876 3292 6928
rect 6092 6953 6101 6987
rect 6101 6953 6135 6987
rect 6135 6953 6144 6987
rect 6092 6944 6144 6953
rect 7380 6987 7432 6996
rect 7380 6953 7389 6987
rect 7389 6953 7423 6987
rect 7423 6953 7432 6987
rect 7380 6944 7432 6953
rect 8208 6944 8260 6996
rect 9496 6944 9548 6996
rect 9772 6944 9824 6996
rect 14648 6987 14700 6996
rect 14648 6953 14657 6987
rect 14657 6953 14691 6987
rect 14691 6953 14700 6987
rect 14648 6944 14700 6953
rect 16948 6944 17000 6996
rect 3056 6851 3108 6860
rect 3056 6817 3065 6851
rect 3065 6817 3099 6851
rect 3099 6817 3108 6851
rect 3056 6808 3108 6817
rect 3608 6808 3660 6860
rect 8852 6876 8904 6928
rect 2228 6740 2280 6792
rect 3148 6740 3200 6792
rect 6828 6808 6880 6860
rect 9036 6808 9088 6860
rect 10968 6851 11020 6860
rect 8300 6783 8352 6792
rect 3608 6672 3660 6724
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 2044 6604 2096 6656
rect 3976 6604 4028 6656
rect 4068 6604 4120 6656
rect 9496 6672 9548 6724
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 11428 6851 11480 6860
rect 11428 6817 11437 6851
rect 11437 6817 11471 6851
rect 11471 6817 11480 6851
rect 11428 6808 11480 6817
rect 13636 6876 13688 6928
rect 11980 6808 12032 6860
rect 12348 6808 12400 6860
rect 12716 6808 12768 6860
rect 14188 6876 14240 6928
rect 15384 6808 15436 6860
rect 16488 6808 16540 6860
rect 16672 6851 16724 6860
rect 16672 6817 16706 6851
rect 16706 6817 16724 6851
rect 16672 6808 16724 6817
rect 11060 6740 11112 6792
rect 11888 6740 11940 6792
rect 14004 6740 14056 6792
rect 14372 6740 14424 6792
rect 16396 6783 16448 6792
rect 16396 6749 16405 6783
rect 16405 6749 16439 6783
rect 16439 6749 16448 6783
rect 16396 6740 16448 6749
rect 18880 6783 18932 6792
rect 18880 6749 18889 6783
rect 18889 6749 18923 6783
rect 18923 6749 18932 6783
rect 18880 6740 18932 6749
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 8392 6604 8444 6656
rect 12440 6647 12492 6656
rect 12440 6613 12449 6647
rect 12449 6613 12483 6647
rect 12483 6613 12492 6647
rect 12440 6604 12492 6613
rect 14004 6647 14056 6656
rect 14004 6613 14013 6647
rect 14013 6613 14047 6647
rect 14047 6613 14056 6647
rect 14004 6604 14056 6613
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 16396 6604 16448 6656
rect 16672 6604 16724 6656
rect 18328 6647 18380 6656
rect 18328 6613 18337 6647
rect 18337 6613 18371 6647
rect 18371 6613 18380 6647
rect 18328 6604 18380 6613
rect 18696 6647 18748 6656
rect 18696 6613 18705 6647
rect 18705 6613 18739 6647
rect 18739 6613 18748 6647
rect 18696 6604 18748 6613
rect 19340 6647 19392 6656
rect 19340 6613 19349 6647
rect 19349 6613 19383 6647
rect 19383 6613 19392 6647
rect 19340 6604 19392 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 3700 6400 3752 6452
rect 4252 6400 4304 6452
rect 2596 6332 2648 6384
rect 3608 6332 3660 6384
rect 4896 6400 4948 6452
rect 5172 6443 5224 6452
rect 5172 6409 5181 6443
rect 5181 6409 5215 6443
rect 5215 6409 5224 6443
rect 5172 6400 5224 6409
rect 8024 6332 8076 6384
rect 5540 6264 5592 6316
rect 8208 6264 8260 6316
rect 8576 6400 8628 6452
rect 9680 6400 9732 6452
rect 11428 6400 11480 6452
rect 12716 6400 12768 6452
rect 15384 6443 15436 6452
rect 15384 6409 15393 6443
rect 15393 6409 15427 6443
rect 15427 6409 15436 6443
rect 15384 6400 15436 6409
rect 15752 6443 15804 6452
rect 15752 6409 15761 6443
rect 15761 6409 15795 6443
rect 15795 6409 15804 6443
rect 15752 6400 15804 6409
rect 16120 6400 16172 6452
rect 16764 6400 16816 6452
rect 11980 6332 12032 6384
rect 11244 6307 11296 6316
rect 11244 6273 11253 6307
rect 11253 6273 11287 6307
rect 11287 6273 11296 6307
rect 11244 6264 11296 6273
rect 16488 6264 16540 6316
rect 18052 6307 18104 6316
rect 18052 6273 18061 6307
rect 18061 6273 18095 6307
rect 18095 6273 18104 6307
rect 18052 6264 18104 6273
rect 4896 6196 4948 6248
rect 7748 6196 7800 6248
rect 10968 6196 11020 6248
rect 12440 6239 12492 6248
rect 3608 6128 3660 6180
rect 5080 6128 5132 6180
rect 6828 6128 6880 6180
rect 7196 6171 7248 6180
rect 7196 6137 7205 6171
rect 7205 6137 7239 6171
rect 7239 6137 7248 6171
rect 7196 6128 7248 6137
rect 7380 6171 7432 6180
rect 7380 6137 7389 6171
rect 7389 6137 7423 6171
rect 7423 6137 7432 6171
rect 7380 6128 7432 6137
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 3976 6103 4028 6112
rect 3976 6069 3985 6103
rect 3985 6069 4019 6103
rect 4019 6069 4028 6103
rect 3976 6060 4028 6069
rect 6460 6060 6512 6112
rect 6644 6060 6696 6112
rect 7288 6060 7340 6112
rect 10876 6128 10928 6180
rect 12440 6205 12449 6239
rect 12449 6205 12483 6239
rect 12483 6205 12492 6239
rect 12440 6196 12492 6205
rect 12348 6128 12400 6180
rect 16488 6171 16540 6180
rect 16488 6137 16497 6171
rect 16497 6137 16531 6171
rect 16531 6137 16540 6171
rect 16488 6128 16540 6137
rect 18972 6128 19024 6180
rect 9680 6060 9732 6112
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 11888 6060 11940 6069
rect 15752 6060 15804 6112
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 19432 6103 19484 6112
rect 19432 6069 19441 6103
rect 19441 6069 19475 6103
rect 19475 6069 19484 6103
rect 19432 6060 19484 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 3516 5899 3568 5908
rect 3516 5865 3525 5899
rect 3525 5865 3559 5899
rect 3559 5865 3568 5899
rect 3516 5856 3568 5865
rect 3608 5856 3660 5908
rect 5080 5899 5132 5908
rect 5080 5865 5089 5899
rect 5089 5865 5123 5899
rect 5123 5865 5132 5899
rect 5080 5856 5132 5865
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 7288 5899 7340 5908
rect 7288 5865 7297 5899
rect 7297 5865 7331 5899
rect 7331 5865 7340 5899
rect 7288 5856 7340 5865
rect 9496 5899 9548 5908
rect 9496 5865 9505 5899
rect 9505 5865 9539 5899
rect 9539 5865 9548 5899
rect 9496 5856 9548 5865
rect 12716 5856 12768 5908
rect 4068 5788 4120 5840
rect 4620 5831 4672 5840
rect 4620 5797 4629 5831
rect 4629 5797 4663 5831
rect 4663 5797 4672 5831
rect 4620 5788 4672 5797
rect 4712 5831 4764 5840
rect 4712 5797 4721 5831
rect 4721 5797 4755 5831
rect 4755 5797 4764 5831
rect 4712 5788 4764 5797
rect 1860 5720 1912 5772
rect 2780 5720 2832 5772
rect 3976 5720 4028 5772
rect 4436 5763 4488 5772
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 4252 5652 4304 5704
rect 5448 5720 5500 5772
rect 6184 5763 6236 5772
rect 6184 5729 6218 5763
rect 6218 5729 6236 5763
rect 6184 5720 6236 5729
rect 11428 5788 11480 5840
rect 14004 5831 14056 5840
rect 14004 5797 14013 5831
rect 14013 5797 14047 5831
rect 14047 5797 14056 5831
rect 14004 5788 14056 5797
rect 18972 5899 19024 5908
rect 18972 5865 18981 5899
rect 18981 5865 19015 5899
rect 19015 5865 19024 5899
rect 18972 5856 19024 5865
rect 19524 5856 19576 5908
rect 15936 5788 15988 5840
rect 16396 5831 16448 5840
rect 16396 5797 16405 5831
rect 16405 5797 16439 5831
rect 16439 5797 16448 5831
rect 16396 5788 16448 5797
rect 16488 5831 16540 5840
rect 16488 5797 16497 5831
rect 16497 5797 16531 5831
rect 16531 5797 16540 5831
rect 16488 5788 16540 5797
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 9956 5763 10008 5772
rect 9956 5729 9965 5763
rect 9965 5729 9999 5763
rect 9999 5729 10008 5763
rect 9956 5720 10008 5729
rect 10876 5720 10928 5772
rect 13820 5720 13872 5772
rect 15660 5720 15712 5772
rect 17868 5763 17920 5772
rect 17868 5729 17902 5763
rect 17902 5729 17920 5763
rect 17868 5720 17920 5729
rect 13912 5695 13964 5704
rect 3056 5584 3108 5636
rect 4160 5627 4212 5636
rect 4160 5593 4169 5627
rect 4169 5593 4203 5627
rect 4203 5593 4212 5627
rect 4160 5584 4212 5593
rect 1952 5559 2004 5568
rect 1952 5525 1961 5559
rect 1961 5525 1995 5559
rect 1995 5525 2004 5559
rect 1952 5516 2004 5525
rect 2688 5516 2740 5568
rect 5540 5516 5592 5568
rect 13912 5661 13921 5695
rect 13921 5661 13955 5695
rect 13955 5661 13964 5695
rect 13912 5652 13964 5661
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20352 5652 20404 5661
rect 7840 5627 7892 5636
rect 7840 5593 7849 5627
rect 7849 5593 7883 5627
rect 7883 5593 7892 5627
rect 7840 5584 7892 5593
rect 11980 5584 12032 5636
rect 14280 5584 14332 5636
rect 15752 5584 15804 5636
rect 15844 5584 15896 5636
rect 6092 5516 6144 5568
rect 8300 5559 8352 5568
rect 8300 5525 8309 5559
rect 8309 5525 8343 5559
rect 8343 5525 8352 5559
rect 8300 5516 8352 5525
rect 8576 5559 8628 5568
rect 8576 5525 8585 5559
rect 8585 5525 8619 5559
rect 8619 5525 8628 5559
rect 8576 5516 8628 5525
rect 9036 5559 9088 5568
rect 9036 5525 9045 5559
rect 9045 5525 9079 5559
rect 9079 5525 9088 5559
rect 9036 5516 9088 5525
rect 9772 5516 9824 5568
rect 10876 5559 10928 5568
rect 10876 5525 10885 5559
rect 10885 5525 10919 5559
rect 10919 5525 10928 5559
rect 10876 5516 10928 5525
rect 12348 5559 12400 5568
rect 12348 5525 12357 5559
rect 12357 5525 12391 5559
rect 12391 5525 12400 5559
rect 12348 5516 12400 5525
rect 13820 5516 13872 5568
rect 20076 5559 20128 5568
rect 20076 5525 20085 5559
rect 20085 5525 20119 5559
rect 20119 5525 20128 5559
rect 20076 5516 20128 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1860 5355 1912 5364
rect 1860 5321 1869 5355
rect 1869 5321 1903 5355
rect 1903 5321 1912 5355
rect 1860 5312 1912 5321
rect 4068 5355 4120 5364
rect 4068 5321 4077 5355
rect 4077 5321 4111 5355
rect 4111 5321 4120 5355
rect 4068 5312 4120 5321
rect 4528 5312 4580 5364
rect 7012 5355 7064 5364
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 7288 5312 7340 5364
rect 2596 5244 2648 5296
rect 4620 5244 4672 5296
rect 5080 5244 5132 5296
rect 2780 5176 2832 5228
rect 4068 5176 4120 5228
rect 3608 5108 3660 5160
rect 5448 5176 5500 5228
rect 8484 5355 8536 5364
rect 8484 5321 8493 5355
rect 8493 5321 8527 5355
rect 8527 5321 8536 5355
rect 8484 5312 8536 5321
rect 9864 5312 9916 5364
rect 10968 5355 11020 5364
rect 10968 5321 10977 5355
rect 10977 5321 11011 5355
rect 11011 5321 11020 5355
rect 10968 5312 11020 5321
rect 12440 5312 12492 5364
rect 14464 5312 14516 5364
rect 15384 5312 15436 5364
rect 15936 5355 15988 5364
rect 15936 5321 15945 5355
rect 15945 5321 15979 5355
rect 15979 5321 15988 5355
rect 15936 5312 15988 5321
rect 16396 5312 16448 5364
rect 18880 5312 18932 5364
rect 19432 5355 19484 5364
rect 19432 5321 19441 5355
rect 19441 5321 19475 5355
rect 19475 5321 19484 5355
rect 19432 5312 19484 5321
rect 19984 5312 20036 5364
rect 20996 5355 21048 5364
rect 20996 5321 21005 5355
rect 21005 5321 21039 5355
rect 21039 5321 21048 5355
rect 20996 5312 21048 5321
rect 16488 5287 16540 5296
rect 16488 5253 16497 5287
rect 16497 5253 16531 5287
rect 16531 5253 16540 5287
rect 16488 5244 16540 5253
rect 13360 5176 13412 5228
rect 17224 5176 17276 5228
rect 19524 5244 19576 5296
rect 20076 5176 20128 5228
rect 4712 5108 4764 5160
rect 6092 5108 6144 5160
rect 11152 5151 11204 5160
rect 3332 5040 3384 5092
rect 3792 5040 3844 5092
rect 4160 5040 4212 5092
rect 6736 5040 6788 5092
rect 11152 5117 11161 5151
rect 11161 5117 11195 5151
rect 11195 5117 11204 5151
rect 11152 5108 11204 5117
rect 12440 5151 12492 5160
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 12440 5108 12492 5117
rect 14096 5108 14148 5160
rect 17408 5108 17460 5160
rect 17960 5108 18012 5160
rect 18512 5108 18564 5160
rect 20720 5151 20772 5160
rect 20720 5117 20729 5151
rect 20729 5117 20763 5151
rect 20763 5117 20772 5151
rect 20720 5108 20772 5117
rect 7656 5040 7708 5092
rect 8760 5040 8812 5092
rect 9588 5040 9640 5092
rect 12716 5040 12768 5092
rect 4436 4972 4488 5024
rect 5448 5015 5500 5024
rect 5448 4981 5457 5015
rect 5457 4981 5491 5015
rect 5491 4981 5500 5015
rect 5448 4972 5500 4981
rect 6092 4972 6144 5024
rect 8668 4972 8720 5024
rect 9128 4972 9180 5024
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 11428 4972 11480 5024
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 12624 5015 12676 5024
rect 12624 4981 12633 5015
rect 12633 4981 12667 5015
rect 12667 4981 12676 5015
rect 12624 4972 12676 4981
rect 14280 5040 14332 5092
rect 18604 5083 18656 5092
rect 18604 5049 18613 5083
rect 18613 5049 18647 5083
rect 18647 5049 18656 5083
rect 18604 5040 18656 5049
rect 19616 5040 19668 5092
rect 19984 5083 20036 5092
rect 19984 5049 19993 5083
rect 19993 5049 20027 5083
rect 20027 5049 20036 5083
rect 19984 5040 20036 5049
rect 13912 4972 13964 5024
rect 14832 4972 14884 5024
rect 16948 5015 17000 5024
rect 16948 4981 16957 5015
rect 16957 4981 16991 5015
rect 16991 4981 17000 5015
rect 16948 4972 17000 4981
rect 17224 4972 17276 5024
rect 17592 4972 17644 5024
rect 20444 4972 20496 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 4620 4811 4672 4820
rect 4620 4777 4629 4811
rect 4629 4777 4663 4811
rect 4663 4777 4672 4811
rect 4620 4768 4672 4777
rect 5540 4768 5592 4820
rect 2964 4743 3016 4752
rect 2964 4709 2973 4743
rect 2973 4709 3007 4743
rect 3007 4709 3016 4743
rect 2964 4700 3016 4709
rect 4712 4743 4764 4752
rect 4712 4709 4721 4743
rect 4721 4709 4755 4743
rect 4755 4709 4764 4743
rect 4712 4700 4764 4709
rect 4068 4632 4120 4684
rect 6184 4768 6236 4820
rect 8760 4811 8812 4820
rect 8760 4777 8769 4811
rect 8769 4777 8803 4811
rect 8803 4777 8812 4811
rect 8760 4768 8812 4777
rect 10140 4768 10192 4820
rect 12164 4768 12216 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 14096 4811 14148 4820
rect 14096 4777 14105 4811
rect 14105 4777 14139 4811
rect 14139 4777 14148 4811
rect 14096 4768 14148 4777
rect 15568 4768 15620 4820
rect 16948 4768 17000 4820
rect 19524 4768 19576 4820
rect 6828 4743 6880 4752
rect 6828 4709 6862 4743
rect 6862 4709 6880 4743
rect 6828 4700 6880 4709
rect 13544 4700 13596 4752
rect 6552 4675 6604 4684
rect 6552 4641 6561 4675
rect 6561 4641 6595 4675
rect 6595 4641 6604 4675
rect 6552 4632 6604 4641
rect 9956 4632 10008 4684
rect 12348 4632 12400 4684
rect 13268 4632 13320 4684
rect 16672 4632 16724 4684
rect 17224 4632 17276 4684
rect 17408 4675 17460 4684
rect 17408 4641 17442 4675
rect 17442 4641 17460 4675
rect 17408 4632 17460 4641
rect 19616 4675 19668 4684
rect 19616 4641 19625 4675
rect 19625 4641 19659 4675
rect 19659 4641 19668 4675
rect 19616 4632 19668 4641
rect 20904 4675 20956 4684
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 2504 4539 2556 4548
rect 2504 4505 2513 4539
rect 2513 4505 2547 4539
rect 2547 4505 2556 4539
rect 2504 4496 2556 4505
rect 1768 4428 1820 4480
rect 2872 4428 2924 4480
rect 3884 4564 3936 4616
rect 9864 4564 9916 4616
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 4804 4496 4856 4548
rect 9772 4539 9824 4548
rect 9772 4505 9781 4539
rect 9781 4505 9815 4539
rect 9815 4505 9824 4539
rect 9772 4496 9824 4505
rect 12348 4496 12400 4548
rect 3516 4471 3568 4480
rect 3516 4437 3525 4471
rect 3525 4437 3559 4471
rect 3559 4437 3568 4471
rect 3516 4428 3568 4437
rect 4344 4428 4396 4480
rect 6736 4428 6788 4480
rect 8944 4428 8996 4480
rect 10968 4428 11020 4480
rect 14004 4496 14056 4548
rect 16212 4496 16264 4548
rect 16580 4496 16632 4548
rect 20536 4564 20588 4616
rect 18512 4539 18564 4548
rect 18512 4505 18521 4539
rect 18521 4505 18555 4539
rect 18555 4505 18564 4539
rect 18512 4496 18564 4505
rect 20720 4496 20772 4548
rect 13728 4428 13780 4480
rect 15660 4471 15712 4480
rect 15660 4437 15669 4471
rect 15669 4437 15703 4471
rect 15703 4437 15712 4471
rect 15660 4428 15712 4437
rect 16856 4428 16908 4480
rect 19432 4471 19484 4480
rect 19432 4437 19441 4471
rect 19441 4437 19475 4471
rect 19475 4437 19484 4471
rect 19432 4428 19484 4437
rect 19892 4428 19944 4480
rect 21088 4471 21140 4480
rect 21088 4437 21097 4471
rect 21097 4437 21131 4471
rect 21131 4437 21140 4471
rect 21088 4428 21140 4437
rect 21456 4471 21508 4480
rect 21456 4437 21465 4471
rect 21465 4437 21499 4471
rect 21499 4437 21508 4471
rect 21456 4428 21508 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2964 4224 3016 4276
rect 4620 4267 4672 4276
rect 4620 4233 4629 4267
rect 4629 4233 4663 4267
rect 4663 4233 4672 4267
rect 4620 4224 4672 4233
rect 6828 4224 6880 4276
rect 10140 4267 10192 4276
rect 10140 4233 10149 4267
rect 10149 4233 10183 4267
rect 10183 4233 10192 4267
rect 10140 4224 10192 4233
rect 12072 4224 12124 4276
rect 13636 4224 13688 4276
rect 6552 4199 6604 4208
rect 6552 4165 6561 4199
rect 6561 4165 6595 4199
rect 6595 4165 6604 4199
rect 6552 4156 6604 4165
rect 7288 4156 7340 4208
rect 10692 4199 10744 4208
rect 2136 4088 2188 4140
rect 2228 4088 2280 4140
rect 4068 4088 4120 4140
rect 5724 4131 5776 4140
rect 5724 4097 5733 4131
rect 5733 4097 5767 4131
rect 5767 4097 5776 4131
rect 5724 4088 5776 4097
rect 7380 4088 7432 4140
rect 10692 4165 10701 4199
rect 10701 4165 10735 4199
rect 10735 4165 10744 4199
rect 10692 4156 10744 4165
rect 11980 4156 12032 4208
rect 14464 4224 14516 4276
rect 15568 4224 15620 4276
rect 16580 4224 16632 4276
rect 19524 4224 19576 4276
rect 20260 4224 20312 4276
rect 20904 4224 20956 4276
rect 15660 4156 15712 4208
rect 19616 4199 19668 4208
rect 12164 4088 12216 4140
rect 13360 4088 13412 4140
rect 19616 4165 19625 4199
rect 19625 4165 19659 4199
rect 19659 4165 19668 4199
rect 19616 4156 19668 4165
rect 2872 4020 2924 4072
rect 3976 4063 4028 4072
rect 3976 4029 3985 4063
rect 3985 4029 4019 4063
rect 4019 4029 4028 4063
rect 3976 4020 4028 4029
rect 6460 4020 6512 4072
rect 2228 3952 2280 4004
rect 2780 3952 2832 4004
rect 4344 3952 4396 4004
rect 5540 3952 5592 4004
rect 6276 3952 6328 4004
rect 9864 4020 9916 4072
rect 11888 4020 11940 4072
rect 12348 4020 12400 4072
rect 20168 4063 20220 4072
rect 20168 4029 20177 4063
rect 20177 4029 20211 4063
rect 20211 4029 20220 4063
rect 20168 4020 20220 4029
rect 21272 4063 21324 4072
rect 21272 4029 21281 4063
rect 21281 4029 21315 4063
rect 21315 4029 21324 4063
rect 21272 4020 21324 4029
rect 7104 3995 7156 4004
rect 7104 3961 7113 3995
rect 7113 3961 7147 3995
rect 7147 3961 7156 3995
rect 7104 3952 7156 3961
rect 8944 3952 8996 4004
rect 2596 3927 2648 3936
rect 2596 3893 2605 3927
rect 2605 3893 2639 3927
rect 2639 3893 2648 3927
rect 2596 3884 2648 3893
rect 4068 3884 4120 3936
rect 4160 3927 4212 3936
rect 4160 3893 4169 3927
rect 4169 3893 4203 3927
rect 4203 3893 4212 3927
rect 4160 3884 4212 3893
rect 5632 3884 5684 3936
rect 8208 3884 8260 3936
rect 9496 3927 9548 3936
rect 9496 3893 9505 3927
rect 9505 3893 9539 3927
rect 9539 3893 9548 3927
rect 9496 3884 9548 3893
rect 10140 3884 10192 3936
rect 11060 3884 11112 3936
rect 12256 3952 12308 4004
rect 12716 3995 12768 4004
rect 12716 3961 12725 3995
rect 12725 3961 12759 3995
rect 12759 3961 12768 3995
rect 12716 3952 12768 3961
rect 13544 3952 13596 4004
rect 14372 3952 14424 4004
rect 16948 3995 17000 4004
rect 16948 3961 16957 3995
rect 16957 3961 16991 3995
rect 16991 3961 17000 3995
rect 16948 3952 17000 3961
rect 17408 3952 17460 4004
rect 18328 3995 18380 4004
rect 18328 3961 18337 3995
rect 18337 3961 18371 3995
rect 18371 3961 18380 3995
rect 18328 3952 18380 3961
rect 19432 3952 19484 4004
rect 20076 3952 20128 4004
rect 13176 3884 13228 3936
rect 13636 3884 13688 3936
rect 14464 3884 14516 3936
rect 16212 3927 16264 3936
rect 16212 3893 16221 3927
rect 16221 3893 16255 3927
rect 16255 3893 16264 3927
rect 16212 3884 16264 3893
rect 16856 3927 16908 3936
rect 16856 3893 16865 3927
rect 16865 3893 16899 3927
rect 16899 3893 16908 3927
rect 16856 3884 16908 3893
rect 20352 3927 20404 3936
rect 20352 3893 20361 3927
rect 20361 3893 20395 3927
rect 20395 3893 20404 3927
rect 20352 3884 20404 3893
rect 22376 3927 22428 3936
rect 22376 3893 22385 3927
rect 22385 3893 22419 3927
rect 22419 3893 22428 3927
rect 22376 3884 22428 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2136 3723 2188 3732
rect 2136 3689 2145 3723
rect 2145 3689 2179 3723
rect 2179 3689 2188 3723
rect 2136 3680 2188 3689
rect 3240 3680 3292 3732
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 5540 3680 5592 3732
rect 6000 3680 6052 3732
rect 6460 3723 6512 3732
rect 6460 3689 6469 3723
rect 6469 3689 6503 3723
rect 6503 3689 6512 3723
rect 6460 3680 6512 3689
rect 2596 3612 2648 3664
rect 3608 3612 3660 3664
rect 4068 3612 4120 3664
rect 4620 3655 4672 3664
rect 4620 3621 4629 3655
rect 4629 3621 4663 3655
rect 4663 3621 4672 3655
rect 4620 3612 4672 3621
rect 6092 3612 6144 3664
rect 7288 3612 7340 3664
rect 8484 3680 8536 3732
rect 8944 3723 8996 3732
rect 8944 3689 8953 3723
rect 8953 3689 8987 3723
rect 8987 3689 8996 3723
rect 8944 3680 8996 3689
rect 9956 3680 10008 3732
rect 10784 3680 10836 3732
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 3516 3587 3568 3596
rect 3516 3553 3525 3587
rect 3525 3553 3559 3587
rect 3559 3553 3568 3587
rect 3516 3544 3568 3553
rect 3976 3544 4028 3596
rect 6736 3544 6788 3596
rect 7840 3587 7892 3596
rect 7840 3553 7849 3587
rect 7849 3553 7883 3587
rect 7883 3553 7892 3587
rect 7840 3544 7892 3553
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 6552 3476 6604 3528
rect 7472 3476 7524 3528
rect 9864 3612 9916 3664
rect 12624 3680 12676 3732
rect 13820 3723 13872 3732
rect 13820 3689 13829 3723
rect 13829 3689 13863 3723
rect 13863 3689 13872 3723
rect 13820 3680 13872 3689
rect 14832 3680 14884 3732
rect 16948 3680 17000 3732
rect 21364 3680 21416 3732
rect 13268 3612 13320 3664
rect 13728 3612 13780 3664
rect 16028 3612 16080 3664
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 10876 3544 10928 3596
rect 11060 3587 11112 3596
rect 11060 3553 11094 3587
rect 11094 3553 11112 3587
rect 11060 3544 11112 3553
rect 16488 3612 16540 3664
rect 16672 3544 16724 3596
rect 18696 3544 18748 3596
rect 19064 3587 19116 3596
rect 19064 3553 19073 3587
rect 19073 3553 19107 3587
rect 19107 3553 19116 3587
rect 19064 3544 19116 3553
rect 20904 3587 20956 3596
rect 20904 3553 20913 3587
rect 20913 3553 20947 3587
rect 20947 3553 20956 3587
rect 20904 3544 20956 3553
rect 22008 3587 22060 3596
rect 22008 3553 22017 3587
rect 22017 3553 22051 3587
rect 22051 3553 22060 3587
rect 22008 3544 22060 3553
rect 14464 3476 14516 3528
rect 16580 3519 16632 3528
rect 16580 3485 16589 3519
rect 16589 3485 16623 3519
rect 16623 3485 16632 3519
rect 16580 3476 16632 3485
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 3700 3408 3752 3460
rect 3884 3408 3936 3460
rect 4252 3408 4304 3460
rect 5632 3408 5684 3460
rect 6184 3408 6236 3460
rect 7380 3408 7432 3460
rect 8300 3408 8352 3460
rect 13360 3451 13412 3460
rect 13360 3417 13369 3451
rect 13369 3417 13403 3451
rect 13403 3417 13412 3451
rect 13360 3408 13412 3417
rect 14372 3451 14424 3460
rect 14372 3417 14381 3451
rect 14381 3417 14415 3451
rect 14415 3417 14424 3451
rect 14372 3408 14424 3417
rect 16488 3408 16540 3460
rect 22744 3408 22796 3460
rect 2504 3383 2556 3392
rect 2504 3349 2513 3383
rect 2513 3349 2547 3383
rect 2547 3349 2556 3383
rect 2504 3340 2556 3349
rect 6368 3340 6420 3392
rect 7196 3340 7248 3392
rect 9680 3340 9732 3392
rect 19248 3383 19300 3392
rect 19248 3349 19257 3383
rect 19257 3349 19291 3383
rect 19291 3349 19300 3383
rect 19248 3340 19300 3349
rect 19984 3383 20036 3392
rect 19984 3349 19993 3383
rect 19993 3349 20027 3383
rect 20027 3349 20036 3383
rect 19984 3340 20036 3349
rect 20260 3340 20312 3392
rect 21824 3383 21876 3392
rect 21824 3349 21833 3383
rect 21833 3349 21867 3383
rect 21867 3349 21876 3383
rect 21824 3340 21876 3349
rect 22192 3383 22244 3392
rect 22192 3349 22201 3383
rect 22201 3349 22235 3383
rect 22235 3349 22244 3383
rect 22192 3340 22244 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1768 3179 1820 3188
rect 1768 3145 1777 3179
rect 1777 3145 1811 3179
rect 1811 3145 1820 3179
rect 1768 3136 1820 3145
rect 2596 3136 2648 3188
rect 3240 3179 3292 3188
rect 3240 3145 3249 3179
rect 3249 3145 3283 3179
rect 3283 3145 3292 3179
rect 3240 3136 3292 3145
rect 6092 3136 6144 3188
rect 2320 3111 2372 3120
rect 2320 3077 2329 3111
rect 2329 3077 2363 3111
rect 2363 3077 2372 3111
rect 2320 3068 2372 3077
rect 2780 3000 2832 3052
rect 7288 3136 7340 3188
rect 8484 3179 8536 3188
rect 8484 3145 8493 3179
rect 8493 3145 8527 3179
rect 8527 3145 8536 3179
rect 8484 3136 8536 3145
rect 10876 3136 10928 3188
rect 14464 3179 14516 3188
rect 14464 3145 14473 3179
rect 14473 3145 14507 3179
rect 14507 3145 14516 3179
rect 14464 3136 14516 3145
rect 16856 3136 16908 3188
rect 19064 3179 19116 3188
rect 19064 3145 19073 3179
rect 19073 3145 19107 3179
rect 19107 3145 19116 3179
rect 19064 3136 19116 3145
rect 19340 3136 19392 3188
rect 17132 3068 17184 3120
rect 2228 2932 2280 2984
rect 2596 2975 2648 2984
rect 2596 2941 2605 2975
rect 2605 2941 2639 2975
rect 2639 2941 2648 2975
rect 2596 2932 2648 2941
rect 6552 2975 6604 2984
rect 6552 2941 6561 2975
rect 6561 2941 6595 2975
rect 6595 2941 6604 2975
rect 6552 2932 6604 2941
rect 7380 2975 7432 2984
rect 7380 2941 7414 2975
rect 7414 2941 7432 2975
rect 7380 2932 7432 2941
rect 7840 2932 7892 2984
rect 10876 2932 10928 2984
rect 14924 2975 14976 2984
rect 14924 2941 14933 2975
rect 14933 2941 14967 2975
rect 14967 2941 14976 2975
rect 14924 2932 14976 2941
rect 16580 2932 16632 2984
rect 3976 2864 4028 2916
rect 9956 2864 10008 2916
rect 12072 2864 12124 2916
rect 12624 2864 12676 2916
rect 14832 2864 14884 2916
rect 18144 3000 18196 3052
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 18696 3000 18748 3009
rect 19616 3136 19668 3188
rect 22008 3179 22060 3188
rect 22008 3145 22017 3179
rect 22017 3145 22051 3179
rect 22051 3145 22060 3179
rect 22008 3136 22060 3145
rect 23848 3068 23900 3120
rect 23664 3043 23716 3052
rect 23664 3009 23673 3043
rect 23673 3009 23707 3043
rect 23707 3009 23716 3043
rect 23664 3000 23716 3009
rect 19340 2932 19392 2984
rect 20628 2932 20680 2984
rect 21364 2932 21416 2984
rect 20168 2907 20220 2916
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 3700 2839 3752 2848
rect 2780 2796 2832 2805
rect 3700 2805 3709 2839
rect 3709 2805 3743 2839
rect 3743 2805 3752 2839
rect 3700 2796 3752 2805
rect 4344 2796 4396 2848
rect 9496 2796 9548 2848
rect 11152 2796 11204 2848
rect 11244 2796 11296 2848
rect 11704 2796 11756 2848
rect 16488 2796 16540 2848
rect 20168 2873 20177 2907
rect 20177 2873 20211 2907
rect 20211 2873 20220 2907
rect 20168 2864 20220 2873
rect 20904 2839 20956 2848
rect 20904 2805 20913 2839
rect 20913 2805 20947 2839
rect 20947 2805 20956 2839
rect 20904 2796 20956 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 4896 2592 4948 2644
rect 7288 2592 7340 2644
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 10692 2592 10744 2644
rect 11152 2592 11204 2644
rect 3976 2524 4028 2576
rect 4344 2567 4396 2576
rect 4344 2533 4378 2567
rect 4378 2533 4396 2567
rect 4344 2524 4396 2533
rect 3700 2456 3752 2508
rect 9772 2524 9824 2576
rect 11244 2524 11296 2576
rect 12440 2567 12492 2576
rect 12440 2533 12449 2567
rect 12449 2533 12483 2567
rect 12483 2533 12492 2567
rect 12440 2524 12492 2533
rect 12716 2524 12768 2576
rect 13176 2567 13228 2576
rect 13176 2533 13185 2567
rect 13185 2533 13219 2567
rect 13219 2533 13228 2567
rect 13176 2524 13228 2533
rect 14924 2592 14976 2644
rect 11152 2499 11204 2508
rect 11152 2465 11161 2499
rect 11161 2465 11195 2499
rect 11195 2465 11204 2499
rect 11152 2456 11204 2465
rect 13452 2456 13504 2508
rect 16672 2592 16724 2644
rect 19340 2592 19392 2644
rect 20168 2592 20220 2644
rect 20628 2592 20680 2644
rect 23296 2592 23348 2644
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 3608 2388 3660 2440
rect 14464 2388 14516 2440
rect 16580 2456 16632 2508
rect 19892 2499 19944 2508
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 20444 2456 20496 2508
rect 22468 2499 22520 2508
rect 22468 2465 22477 2499
rect 22477 2465 22511 2499
rect 22511 2465 22520 2499
rect 22468 2456 22520 2465
rect 24032 2499 24084 2508
rect 24032 2465 24041 2499
rect 24041 2465 24075 2499
rect 24075 2465 24084 2499
rect 24032 2456 24084 2465
rect 5356 2320 5408 2372
rect 6000 2320 6052 2372
rect 11888 2320 11940 2372
rect 12256 2320 12308 2372
rect 14372 2363 14424 2372
rect 14372 2329 14381 2363
rect 14381 2329 14415 2363
rect 14415 2329 14424 2363
rect 14372 2320 14424 2329
rect 18328 2320 18380 2372
rect 20628 2320 20680 2372
rect 24124 2320 24176 2372
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 2780 2252 2832 2304
rect 4712 2252 4764 2304
rect 11520 2295 11572 2304
rect 11520 2261 11529 2295
rect 11529 2261 11563 2295
rect 11563 2261 11572 2295
rect 11520 2252 11572 2261
rect 18052 2295 18104 2304
rect 18052 2261 18061 2295
rect 18061 2261 18095 2295
rect 18095 2261 18104 2295
rect 18052 2252 18104 2261
rect 22192 2295 22244 2304
rect 22192 2261 22201 2295
rect 22201 2261 22235 2295
rect 22235 2261 22244 2295
rect 22192 2252 22244 2261
rect 24216 2295 24268 2304
rect 24216 2261 24225 2295
rect 24225 2261 24259 2295
rect 24259 2261 24268 2295
rect 24216 2252 24268 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 12900 1844 12952 1896
rect 14188 1844 14240 1896
rect 15476 552 15528 604
rect 16856 552 16908 604
rect 20720 552 20772 604
rect 21180 552 21232 604
<< metal2 >>
rect 202 27520 258 28000
rect 662 27520 718 28000
rect 1214 27520 1270 28000
rect 1766 27520 1822 28000
rect 2318 27520 2374 28000
rect 2870 27520 2926 28000
rect 3238 27704 3294 27713
rect 3238 27639 3294 27648
rect 216 23633 244 27520
rect 676 24313 704 27520
rect 1228 24834 1256 27520
rect 1674 25800 1730 25809
rect 1674 25735 1730 25744
rect 1228 24818 1440 24834
rect 1228 24812 1452 24818
rect 1228 24806 1400 24812
rect 1400 24754 1452 24760
rect 662 24304 718 24313
rect 662 24239 718 24248
rect 1412 23769 1440 24754
rect 1490 24576 1546 24585
rect 1490 24511 1546 24520
rect 1504 23866 1532 24511
rect 1688 24342 1716 25735
rect 1780 24721 1808 27520
rect 2226 27024 2282 27033
rect 2226 26959 2282 26968
rect 1766 24712 1822 24721
rect 1766 24647 1822 24656
rect 1676 24336 1728 24342
rect 1676 24278 1728 24284
rect 1492 23860 1544 23866
rect 1492 23802 1544 23808
rect 1398 23760 1454 23769
rect 1398 23695 1454 23704
rect 1412 23662 1440 23695
rect 1400 23656 1452 23662
rect 202 23624 258 23633
rect 1400 23598 1452 23604
rect 202 23559 258 23568
rect 1688 23322 1716 24278
rect 2044 23724 2096 23730
rect 2044 23666 2096 23672
rect 1950 23624 2006 23633
rect 1950 23559 2006 23568
rect 1964 23526 1992 23559
rect 1952 23520 2004 23526
rect 1952 23462 2004 23468
rect 1964 23322 1992 23462
rect 1676 23316 1728 23322
rect 1676 23258 1728 23264
rect 1952 23316 2004 23322
rect 1952 23258 2004 23264
rect 1964 23089 1992 23258
rect 1950 23080 2006 23089
rect 1950 23015 2006 23024
rect 2056 22234 2084 23666
rect 2044 22228 2096 22234
rect 2044 22170 2096 22176
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1596 20602 1624 21286
rect 2240 21026 2268 26959
rect 2332 25498 2360 27520
rect 2320 25492 2372 25498
rect 2320 25434 2372 25440
rect 2884 24954 2912 27520
rect 2872 24948 2924 24954
rect 2872 24890 2924 24896
rect 3056 24404 3108 24410
rect 3056 24346 3108 24352
rect 2504 24268 2556 24274
rect 2504 24210 2556 24216
rect 2516 23594 2544 24210
rect 3068 23662 3096 24346
rect 3146 24304 3202 24313
rect 3146 24239 3202 24248
rect 3056 23656 3108 23662
rect 3056 23598 3108 23604
rect 2504 23588 2556 23594
rect 2504 23530 2556 23536
rect 3068 23254 3096 23598
rect 3056 23248 3108 23254
rect 2778 23216 2834 23225
rect 3056 23190 3108 23196
rect 2778 23151 2834 23160
rect 2872 23180 2924 23186
rect 2688 22500 2740 22506
rect 2688 22442 2740 22448
rect 2318 21992 2374 22001
rect 2318 21927 2374 21936
rect 2502 21992 2558 22001
rect 2502 21927 2504 21936
rect 2332 21146 2360 21927
rect 2556 21927 2558 21936
rect 2596 21956 2648 21962
rect 2504 21898 2556 21904
rect 2596 21898 2648 21904
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 2516 21457 2544 21490
rect 2502 21448 2558 21457
rect 2502 21383 2558 21392
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 1688 20998 2268 21026
rect 2332 21026 2360 21082
rect 2332 20998 2452 21026
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1400 16516 1452 16522
rect 1400 16458 1452 16464
rect 1308 16448 1360 16454
rect 1308 16390 1360 16396
rect 1320 12782 1348 16390
rect 1412 16046 1440 16458
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1308 12776 1360 12782
rect 1308 12718 1360 12724
rect 1412 12442 1440 15982
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1400 12436 1452 12442
rect 1400 12378 1452 12384
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1412 11286 1440 11494
rect 1400 11280 1452 11286
rect 570 11248 626 11257
rect 1400 11222 1452 11228
rect 570 11183 626 11192
rect 584 4978 612 11183
rect 1504 8537 1532 14758
rect 1596 10441 1624 15302
rect 1688 14958 1716 20998
rect 2320 20936 2372 20942
rect 2320 20878 2372 20884
rect 1860 20800 1912 20806
rect 1860 20742 1912 20748
rect 1872 20398 1900 20742
rect 1860 20392 1912 20398
rect 1860 20334 1912 20340
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1780 19718 1808 20198
rect 1768 19712 1820 19718
rect 1768 19654 1820 19660
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1676 14000 1728 14006
rect 1676 13942 1728 13948
rect 1688 13569 1716 13942
rect 1674 13560 1730 13569
rect 1674 13495 1730 13504
rect 1780 13025 1808 19654
rect 1872 17513 1900 20334
rect 2332 20058 2360 20878
rect 2424 20602 2452 20998
rect 2516 20806 2544 21383
rect 2608 21350 2636 21898
rect 2700 21894 2728 22442
rect 2688 21888 2740 21894
rect 2688 21830 2740 21836
rect 2596 21344 2648 21350
rect 2596 21286 2648 21292
rect 2700 20942 2728 21830
rect 2688 20936 2740 20942
rect 2688 20878 2740 20884
rect 2504 20800 2556 20806
rect 2504 20742 2556 20748
rect 2412 20596 2464 20602
rect 2412 20538 2464 20544
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2424 19394 2452 20538
rect 2700 20330 2728 20878
rect 2688 20324 2740 20330
rect 2688 20266 2740 20272
rect 2700 19718 2728 20266
rect 2688 19712 2740 19718
rect 2688 19654 2740 19660
rect 2700 19514 2728 19654
rect 2688 19508 2740 19514
rect 2792 19496 2820 23151
rect 2872 23122 2924 23128
rect 2884 22166 2912 23122
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 2976 22778 3004 23054
rect 2964 22772 3016 22778
rect 2964 22714 3016 22720
rect 3160 22166 3188 24239
rect 2872 22160 2924 22166
rect 2870 22128 2872 22137
rect 3148 22160 3200 22166
rect 2924 22128 2926 22137
rect 3148 22102 3200 22108
rect 2870 22063 2926 22072
rect 2964 22024 3016 22030
rect 2964 21966 3016 21972
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 2976 21622 3004 21966
rect 2964 21616 3016 21622
rect 2964 21558 3016 21564
rect 2976 19990 3004 21558
rect 3068 21418 3096 21966
rect 3056 21412 3108 21418
rect 3056 21354 3108 21360
rect 3056 20596 3108 20602
rect 3160 20584 3188 22102
rect 3108 20556 3188 20584
rect 3056 20538 3108 20544
rect 3160 20330 3188 20556
rect 3148 20324 3200 20330
rect 3148 20266 3200 20272
rect 2964 19984 3016 19990
rect 2964 19926 3016 19932
rect 2792 19468 3004 19496
rect 2688 19450 2740 19456
rect 2240 19366 2452 19394
rect 2686 19408 2742 19417
rect 1858 17504 1914 17513
rect 1914 17462 1992 17490
rect 1858 17439 1914 17448
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1766 13016 1822 13025
rect 1766 12951 1822 12960
rect 1676 12912 1728 12918
rect 1676 12854 1728 12860
rect 1582 10432 1638 10441
rect 1582 10367 1638 10376
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1490 8528 1546 8537
rect 1490 8463 1546 8472
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1214 7712 1270 7721
rect 1214 7647 1270 7656
rect 216 4950 612 4978
rect 216 480 244 4950
rect 662 3768 718 3777
rect 662 3703 718 3712
rect 676 480 704 3703
rect 1228 480 1256 7647
rect 1412 6225 1440 8366
rect 1596 7177 1624 9454
rect 1582 7168 1638 7177
rect 1582 7103 1638 7112
rect 1398 6216 1454 6225
rect 1398 6151 1454 6160
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1398 3632 1454 3641
rect 1398 3567 1400 3576
rect 1452 3567 1454 3576
rect 1400 3538 1452 3544
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1412 1601 1440 2382
rect 1596 2281 1624 6054
rect 1688 3074 1716 12854
rect 1768 12776 1820 12782
rect 1766 12744 1768 12753
rect 1820 12744 1822 12753
rect 1766 12679 1822 12688
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1780 6089 1808 12582
rect 1872 9602 1900 16934
rect 1964 15910 1992 17462
rect 2240 16250 2268 19366
rect 2686 19343 2742 19352
rect 2780 19372 2832 19378
rect 2412 19304 2464 19310
rect 2412 19246 2464 19252
rect 2320 19236 2372 19242
rect 2320 19178 2372 19184
rect 2332 18970 2360 19178
rect 2320 18964 2372 18970
rect 2320 18906 2372 18912
rect 2332 18290 2360 18906
rect 2424 18834 2452 19246
rect 2504 18896 2556 18902
rect 2504 18838 2556 18844
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2424 17882 2452 18770
rect 2516 18154 2544 18838
rect 2594 18320 2650 18329
rect 2594 18255 2650 18264
rect 2504 18148 2556 18154
rect 2504 18090 2556 18096
rect 2412 17876 2464 17882
rect 2412 17818 2464 17824
rect 2516 17610 2544 18090
rect 2504 17604 2556 17610
rect 2504 17546 2556 17552
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 2240 16114 2268 16186
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 1964 15706 1992 15846
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 2056 15337 2084 15506
rect 2320 15360 2372 15366
rect 2042 15328 2098 15337
rect 2320 15302 2372 15308
rect 2042 15263 2098 15272
rect 2056 15162 2084 15263
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 1964 14278 1992 14894
rect 2044 14612 2096 14618
rect 2044 14554 2096 14560
rect 2056 14385 2084 14554
rect 2042 14376 2098 14385
rect 2042 14311 2098 14320
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 2136 14272 2188 14278
rect 2136 14214 2188 14220
rect 1964 13546 1992 14214
rect 2148 13734 2176 14214
rect 2332 13938 2360 15302
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2226 13832 2282 13841
rect 2226 13767 2228 13776
rect 2280 13767 2282 13776
rect 2228 13738 2280 13744
rect 2136 13728 2188 13734
rect 2134 13696 2136 13705
rect 2188 13696 2190 13705
rect 2134 13631 2190 13640
rect 1964 13518 2176 13546
rect 2240 13530 2268 13738
rect 2148 13410 2176 13518
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2044 13388 2096 13394
rect 2148 13382 2268 13410
rect 2044 13330 2096 13336
rect 1950 13016 2006 13025
rect 2056 12986 2084 13330
rect 1950 12951 2006 12960
rect 2044 12980 2096 12986
rect 1964 12374 1992 12951
rect 2096 12940 2176 12968
rect 2044 12922 2096 12928
rect 1952 12368 2004 12374
rect 1952 12310 2004 12316
rect 1964 11898 1992 12310
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1964 10538 1992 10950
rect 2056 10674 2084 12038
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 1952 10532 2004 10538
rect 1952 10474 2004 10480
rect 1872 9574 1992 9602
rect 1858 9480 1914 9489
rect 1858 9415 1860 9424
rect 1912 9415 1914 9424
rect 1860 9386 1912 9392
rect 1858 8664 1914 8673
rect 1858 8599 1914 8608
rect 1872 8498 1900 8599
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1964 8430 1992 9574
rect 2056 9178 2084 10610
rect 2148 10470 2176 12940
rect 2240 12866 2268 13382
rect 2332 12986 2360 13874
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2240 12838 2360 12866
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2240 11626 2268 12242
rect 2228 11620 2280 11626
rect 2228 11562 2280 11568
rect 2240 11354 2268 11562
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2240 11218 2268 11290
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2240 10266 2268 10542
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2332 8922 2360 12838
rect 2424 11540 2452 16594
rect 2504 16176 2556 16182
rect 2504 16118 2556 16124
rect 2516 11642 2544 16118
rect 2608 15570 2636 18255
rect 2700 18086 2728 19343
rect 2780 19314 2832 19320
rect 2792 18698 2820 19314
rect 2976 19174 3004 19468
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2870 18728 2926 18737
rect 2780 18692 2832 18698
rect 2870 18663 2926 18672
rect 2780 18634 2832 18640
rect 2688 18080 2740 18086
rect 2688 18022 2740 18028
rect 2780 17808 2832 17814
rect 2780 17750 2832 17756
rect 2792 17338 2820 17750
rect 2884 17678 2912 18663
rect 2976 18630 3004 19110
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 3068 18426 3096 18702
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 3068 17814 3096 18158
rect 3056 17808 3108 17814
rect 3056 17750 3108 17756
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2884 17338 2912 17614
rect 3068 17338 3096 17750
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2608 15162 2636 15506
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 14618 2636 14758
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2608 14074 2636 14554
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2700 11801 2728 15302
rect 2792 14822 2820 17274
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2884 14550 2912 17274
rect 3252 17252 3280 27639
rect 3422 27520 3478 28000
rect 3974 27520 4030 28000
rect 4526 27520 4582 28000
rect 5078 27520 5134 28000
rect 5630 27520 5686 28000
rect 6182 27520 6238 28000
rect 6734 27520 6790 28000
rect 7286 27520 7342 28000
rect 7838 27520 7894 28000
rect 8390 27520 8446 28000
rect 8942 27520 8998 28000
rect 9494 27520 9550 28000
rect 10046 27520 10102 28000
rect 10598 27520 10654 28000
rect 11150 27520 11206 28000
rect 11702 27520 11758 28000
rect 12254 27520 12310 28000
rect 12806 27520 12862 28000
rect 13358 27520 13414 28000
rect 13910 27520 13966 28000
rect 14370 27520 14426 28000
rect 14922 27520 14978 28000
rect 15474 27520 15530 28000
rect 16026 27520 16082 28000
rect 16578 27520 16634 28000
rect 17130 27520 17186 28000
rect 17682 27520 17738 28000
rect 18234 27520 18290 28000
rect 18786 27520 18842 28000
rect 19338 27520 19394 28000
rect 19890 27520 19946 28000
rect 20442 27520 20498 28000
rect 20994 27520 21050 28000
rect 21546 27520 21602 28000
rect 22098 27520 22154 28000
rect 22650 27520 22706 28000
rect 23202 27520 23258 28000
rect 23754 27520 23810 28000
rect 24306 27520 24362 28000
rect 24858 27520 24914 28000
rect 25410 27520 25466 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 3436 25430 3464 27520
rect 3424 25424 3476 25430
rect 3424 25366 3476 25372
rect 3436 24750 3464 25366
rect 3516 25356 3568 25362
rect 3516 25298 3568 25304
rect 3528 24886 3556 25298
rect 3608 24948 3660 24954
rect 3608 24890 3660 24896
rect 3516 24880 3568 24886
rect 3516 24822 3568 24828
rect 3424 24744 3476 24750
rect 3424 24686 3476 24692
rect 3330 24440 3386 24449
rect 3528 24410 3556 24822
rect 3330 24375 3386 24384
rect 3516 24404 3568 24410
rect 3344 21049 3372 24375
rect 3516 24346 3568 24352
rect 3516 23588 3568 23594
rect 3516 23530 3568 23536
rect 3528 22574 3556 23530
rect 3620 22642 3648 24890
rect 3698 23896 3754 23905
rect 3698 23831 3754 23840
rect 3712 23089 3740 23831
rect 3988 23361 4016 27520
rect 4066 26344 4122 26353
rect 4066 26279 4068 26288
rect 4120 26279 4122 26288
rect 4068 26250 4120 26256
rect 4436 25152 4488 25158
rect 4066 25120 4122 25129
rect 4436 25094 4488 25100
rect 4066 25055 4122 25064
rect 4080 24886 4108 25055
rect 4068 24880 4120 24886
rect 4068 24822 4120 24828
rect 4448 24818 4476 25094
rect 4436 24812 4488 24818
rect 4436 24754 4488 24760
rect 4068 24608 4120 24614
rect 4436 24608 4488 24614
rect 4068 24550 4120 24556
rect 4434 24576 4436 24585
rect 4488 24576 4490 24585
rect 3974 23352 4030 23361
rect 3974 23287 4030 23296
rect 3698 23080 3754 23089
rect 3698 23015 3754 23024
rect 3976 22772 4028 22778
rect 4080 22760 4108 24550
rect 4434 24511 4490 24520
rect 4436 24064 4488 24070
rect 4436 24006 4488 24012
rect 4448 23322 4476 24006
rect 4436 23316 4488 23322
rect 4436 23258 4488 23264
rect 4252 23180 4304 23186
rect 4252 23122 4304 23128
rect 4160 22772 4212 22778
rect 4080 22732 4160 22760
rect 3976 22714 4028 22720
rect 4160 22714 4212 22720
rect 3988 22681 4016 22714
rect 3974 22672 4030 22681
rect 3608 22636 3660 22642
rect 3974 22607 4030 22616
rect 3608 22578 3660 22584
rect 3516 22568 3568 22574
rect 3516 22510 3568 22516
rect 3528 21486 3556 22510
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3330 21040 3386 21049
rect 3528 21010 3556 21422
rect 3330 20975 3386 20984
rect 3516 21004 3568 21010
rect 3516 20946 3568 20952
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3344 18902 3372 19110
rect 3332 18896 3384 18902
rect 3332 18838 3384 18844
rect 3528 18766 3556 20946
rect 3620 20466 3648 22578
rect 3882 22536 3938 22545
rect 3792 22500 3844 22506
rect 3882 22471 3938 22480
rect 3792 22442 3844 22448
rect 3804 21486 3832 22442
rect 3792 21480 3844 21486
rect 3792 21422 3844 21428
rect 3804 21146 3832 21422
rect 3792 21140 3844 21146
rect 3792 21082 3844 21088
rect 3700 20800 3752 20806
rect 3700 20742 3752 20748
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3620 20058 3648 20402
rect 3712 20398 3740 20742
rect 3700 20392 3752 20398
rect 3700 20334 3752 20340
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3712 19825 3740 20334
rect 3698 19816 3754 19825
rect 3698 19751 3754 19760
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3804 19378 3832 19654
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3528 18426 3556 18702
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3528 17882 3556 18362
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3896 17338 3924 22471
rect 4172 22438 4200 22714
rect 4160 22432 4212 22438
rect 4160 22374 4212 22380
rect 4264 22250 4292 23122
rect 4080 22222 4292 22250
rect 4080 22098 4108 22222
rect 4068 22092 4120 22098
rect 4068 22034 4120 22040
rect 4250 21448 4306 21457
rect 4250 21383 4306 21392
rect 3974 21312 4030 21321
rect 3974 21247 4030 21256
rect 3988 17921 4016 21247
rect 4264 21146 4292 21383
rect 4252 21140 4304 21146
rect 4252 21082 4304 21088
rect 4436 20528 4488 20534
rect 4436 20470 4488 20476
rect 4448 20369 4476 20470
rect 4434 20360 4490 20369
rect 4434 20295 4490 20304
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 4080 18737 4108 19178
rect 4172 18902 4200 20198
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4264 19242 4292 19654
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4252 19236 4304 19242
rect 4252 19178 4304 19184
rect 4264 18970 4292 19178
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4160 18896 4212 18902
rect 4160 18838 4212 18844
rect 4066 18728 4122 18737
rect 4066 18663 4122 18672
rect 4172 18358 4200 18838
rect 4356 18834 4384 19314
rect 4344 18828 4396 18834
rect 4344 18770 4396 18776
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 4066 18184 4122 18193
rect 4066 18119 4122 18128
rect 3974 17912 4030 17921
rect 3974 17847 4030 17856
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 3160 17224 3280 17252
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2884 14074 2912 14486
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2792 12170 2820 12922
rect 2884 12918 2912 13398
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 2872 12912 2924 12918
rect 2870 12880 2872 12889
rect 2924 12880 2926 12889
rect 2870 12815 2926 12824
rect 3068 12646 3096 13126
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3068 12442 3096 12582
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 2976 12238 3004 12310
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2686 11792 2742 11801
rect 2686 11727 2742 11736
rect 2516 11614 2820 11642
rect 2424 11512 2636 11540
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2516 10810 2544 11222
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2240 8894 2360 8922
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 2148 7274 2176 7686
rect 2044 7268 2096 7274
rect 2044 7210 2096 7216
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 2056 6662 2084 7210
rect 2240 6882 2268 8894
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2332 7342 2360 8026
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2332 7002 2360 7278
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2148 6854 2268 6882
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 1766 6080 1822 6089
rect 1766 6015 1822 6024
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1872 5370 1900 5714
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1964 5137 1992 5510
rect 1950 5128 2006 5137
rect 1950 5063 2006 5072
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1780 3194 1808 4422
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1688 3046 1900 3074
rect 1872 2666 1900 3046
rect 2056 2961 2084 6598
rect 2148 6497 2176 6854
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2134 6488 2190 6497
rect 2134 6423 2190 6432
rect 2148 4146 2176 6423
rect 2240 4146 2268 6734
rect 2332 5953 2360 6938
rect 2318 5944 2374 5953
rect 2318 5879 2374 5888
rect 2424 5794 2452 10202
rect 2608 9586 2636 11512
rect 2686 11520 2742 11529
rect 2686 11455 2742 11464
rect 2700 10266 2728 11455
rect 2792 11354 2820 11614
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2884 11098 2912 12038
rect 2976 11540 3004 12174
rect 3160 12102 3188 17224
rect 4080 16810 4108 18119
rect 4080 16794 4200 16810
rect 4080 16788 4212 16794
rect 4080 16782 4160 16788
rect 4160 16730 4212 16736
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3252 15094 3280 15846
rect 3332 15428 3384 15434
rect 3332 15370 3384 15376
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 3252 14958 3280 15030
rect 3344 14958 3372 15370
rect 3424 15360 3476 15366
rect 3424 15302 3476 15308
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3252 13870 3280 14554
rect 3344 14550 3372 14894
rect 3436 14890 3464 15302
rect 3528 15162 3556 15846
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3424 14884 3476 14890
rect 3424 14826 3476 14832
rect 3608 14884 3660 14890
rect 3608 14826 3660 14832
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 3436 14414 3464 14826
rect 3620 14618 3648 14826
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3528 14074 3556 14418
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3252 13530 3280 13806
rect 3528 13530 3556 14010
rect 3240 13524 3292 13530
rect 3516 13524 3568 13530
rect 3240 13466 3292 13472
rect 3436 13484 3516 13512
rect 3252 12306 3280 13466
rect 3240 12300 3292 12306
rect 3240 12242 3292 12248
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3146 11656 3202 11665
rect 3146 11591 3202 11600
rect 3056 11552 3108 11558
rect 2976 11512 3056 11540
rect 3056 11494 3108 11500
rect 2792 11070 2912 11098
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2700 9654 2728 10066
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 7041 2544 7686
rect 2502 7032 2558 7041
rect 2502 6967 2558 6976
rect 2608 6390 2636 9522
rect 2792 9382 2820 11070
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2884 10062 2912 10950
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 2976 10198 3004 10678
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 3068 10146 3096 11494
rect 3160 11218 3188 11591
rect 3252 11218 3280 12242
rect 3436 11694 3464 13484
rect 3516 13466 3568 13472
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3344 10606 3372 11222
rect 3436 11150 3464 11630
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3436 10810 3464 11086
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3344 10266 3372 10542
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2884 9178 2912 9998
rect 2976 9722 3004 10134
rect 3068 10118 3372 10146
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2700 7834 2728 8774
rect 2792 8430 2820 9046
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2962 8936 3018 8945
rect 2884 8634 2912 8910
rect 2962 8871 3018 8880
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2976 7886 3004 8871
rect 3068 8498 3096 8978
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3068 8090 3096 8434
rect 3252 8430 3280 9318
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2964 7880 3016 7886
rect 2870 7848 2926 7857
rect 2700 7806 2870 7834
rect 2964 7822 3016 7828
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2870 7783 2926 7792
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2596 6384 2648 6390
rect 2596 6326 2648 6332
rect 2332 5766 2452 5794
rect 2792 5778 2820 7142
rect 2884 7002 2912 7783
rect 2976 7546 3004 7822
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 3068 6866 3096 7822
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2962 6080 3018 6089
rect 2962 6015 3018 6024
rect 2780 5772 2832 5778
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2148 3738 2176 4082
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 2240 2990 2268 3946
rect 2332 3346 2360 5766
rect 2780 5714 2832 5720
rect 2976 5710 3004 6015
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 3068 5642 3096 6802
rect 3160 6798 3188 8366
rect 3240 8016 3292 8022
rect 3240 7958 3292 7964
rect 3344 7970 3372 10118
rect 3436 8401 3464 10406
rect 3528 10266 3556 11290
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3514 9072 3570 9081
rect 3514 9007 3516 9016
rect 3568 9007 3570 9016
rect 3516 8978 3568 8984
rect 3528 8566 3556 8978
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 3422 8392 3478 8401
rect 3422 8327 3478 8336
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 8090 3464 8230
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3620 8022 3648 11630
rect 3712 9450 3740 15914
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3974 15872 4030 15881
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 11694 3832 15302
rect 3896 13462 3924 15846
rect 3974 15807 4030 15816
rect 3884 13456 3936 13462
rect 3988 13433 4016 15807
rect 4264 15026 4292 18566
rect 4356 18426 4384 18770
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 4436 17876 4488 17882
rect 4436 17818 4488 17824
rect 4448 17678 4476 17818
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4448 17202 4476 17614
rect 4540 17252 4568 27520
rect 4620 24676 4672 24682
rect 4620 24618 4672 24624
rect 4632 24274 4660 24618
rect 4896 24336 4948 24342
rect 4896 24278 4948 24284
rect 4620 24268 4672 24274
rect 4620 24210 4672 24216
rect 4632 23866 4660 24210
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 4632 23186 4660 23802
rect 4710 23760 4766 23769
rect 4710 23695 4766 23704
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4724 23066 4752 23695
rect 4632 23038 4752 23066
rect 4908 23050 4936 24278
rect 4988 24132 5040 24138
rect 4988 24074 5040 24080
rect 5000 23662 5028 24074
rect 4988 23656 5040 23662
rect 4986 23624 4988 23633
rect 5040 23624 5042 23633
rect 4986 23559 5042 23568
rect 4896 23044 4948 23050
rect 4632 20602 4660 23038
rect 4896 22986 4948 22992
rect 4896 22704 4948 22710
rect 4896 22646 4948 22652
rect 4908 22234 4936 22646
rect 4986 22536 5042 22545
rect 4986 22471 5042 22480
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 5000 22114 5028 22471
rect 4908 22086 5028 22114
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 4632 20262 4660 20538
rect 4712 20528 4764 20534
rect 4712 20470 4764 20476
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 4724 19990 4752 20470
rect 4712 19984 4764 19990
rect 4712 19926 4764 19932
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4816 19378 4844 19790
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4540 17224 4752 17252
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 4434 15600 4490 15609
rect 4434 15535 4436 15544
rect 4488 15535 4490 15544
rect 4436 15506 4488 15512
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4080 14278 4108 14962
rect 4264 14822 4292 14962
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4528 14544 4580 14550
rect 4528 14486 4580 14492
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 4080 13462 4108 14214
rect 4540 14074 4568 14486
rect 4528 14068 4580 14074
rect 4448 14028 4528 14056
rect 4068 13456 4120 13462
rect 3884 13398 3936 13404
rect 3974 13424 4030 13433
rect 3896 12986 3924 13398
rect 4068 13398 4120 13404
rect 3974 13359 4030 13368
rect 4158 13288 4214 13297
rect 4158 13223 4160 13232
rect 4212 13223 4214 13232
rect 4160 13194 4212 13200
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3896 12442 3924 12718
rect 4080 12714 4108 13126
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3988 12209 4016 12650
rect 3974 12200 4030 12209
rect 4356 12170 4384 12786
rect 4448 12782 4476 14028
rect 4528 14010 4580 14016
rect 4620 13456 4672 13462
rect 4620 13398 4672 13404
rect 4632 12986 4660 13398
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4436 12368 4488 12374
rect 4434 12336 4436 12345
rect 4488 12336 4490 12345
rect 4434 12271 4490 12280
rect 3974 12135 4030 12144
rect 4344 12164 4396 12170
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3804 11286 3832 11494
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3988 10792 4016 12135
rect 4344 12106 4396 12112
rect 4344 11552 4396 11558
rect 4342 11520 4344 11529
rect 4448 11540 4476 12271
rect 4540 11898 4568 12650
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4396 11520 4476 11540
rect 4398 11512 4476 11520
rect 4342 11455 4398 11464
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 4632 11014 4660 11222
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 3988 10764 4108 10792
rect 3974 10704 4030 10713
rect 3974 10639 4030 10648
rect 3790 10296 3846 10305
rect 3790 10231 3846 10240
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3712 8537 3740 8570
rect 3698 8528 3754 8537
rect 3698 8463 3754 8472
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3608 8016 3660 8022
rect 3252 7041 3280 7958
rect 3344 7942 3464 7970
rect 3608 7958 3660 7964
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3238 7032 3294 7041
rect 3238 6967 3294 6976
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 2688 5568 2740 5574
rect 2778 5536 2834 5545
rect 2740 5516 2778 5522
rect 2688 5510 2778 5516
rect 2700 5494 2778 5510
rect 2778 5471 2834 5480
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2502 4584 2558 4593
rect 2502 4519 2504 4528
rect 2556 4519 2558 4528
rect 2504 4490 2556 4496
rect 2608 4321 2636 5238
rect 2792 5234 2820 5471
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2686 5128 2742 5137
rect 2686 5063 2742 5072
rect 2700 4706 2728 5063
rect 2964 4752 3016 4758
rect 2700 4678 2820 4706
rect 2964 4694 3016 4700
rect 2594 4312 2650 4321
rect 2594 4247 2650 4256
rect 2792 4010 2820 4678
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2884 4078 2912 4422
rect 2976 4282 3004 4694
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2596 3936 2648 3942
rect 2594 3904 2596 3913
rect 2648 3904 2650 3913
rect 2594 3839 2650 3848
rect 2596 3664 2648 3670
rect 2596 3606 2648 3612
rect 2504 3392 2556 3398
rect 2502 3360 2504 3369
rect 2556 3360 2558 3369
rect 2332 3318 2452 3346
rect 2424 3210 2452 3318
rect 2502 3295 2558 3304
rect 2424 3182 2544 3210
rect 2608 3194 2636 3606
rect 2320 3120 2372 3126
rect 2318 3088 2320 3097
rect 2372 3088 2374 3097
rect 2318 3023 2374 3032
rect 2228 2984 2280 2990
rect 2042 2952 2098 2961
rect 2228 2926 2280 2932
rect 2042 2887 2098 2896
rect 2516 2802 2544 3182
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2792 3058 2820 3946
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 1780 2638 1900 2666
rect 2332 2774 2544 2802
rect 1582 2272 1638 2281
rect 1582 2207 1638 2216
rect 1398 1592 1454 1601
rect 1398 1527 1454 1536
rect 1780 480 1808 2638
rect 2332 480 2360 2774
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 1737 2544 2246
rect 2502 1728 2558 1737
rect 2502 1663 2558 1672
rect 2608 649 2636 2926
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2792 2310 2820 2790
rect 2870 2680 2926 2689
rect 2870 2615 2926 2624
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2594 640 2650 649
rect 2594 575 2650 584
rect 2884 480 2912 2615
rect 3160 2281 3188 6734
rect 3252 5137 3280 6870
rect 3238 5128 3294 5137
rect 3344 5098 3372 7414
rect 3238 5063 3294 5072
rect 3332 5092 3384 5098
rect 3252 3738 3280 5063
rect 3332 5034 3384 5040
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3252 3194 3280 3674
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3330 2408 3386 2417
rect 3330 2343 3386 2352
rect 3146 2272 3202 2281
rect 3146 2207 3202 2216
rect 3344 1601 3372 2343
rect 3330 1592 3386 1601
rect 3330 1527 3386 1536
rect 3436 480 3464 7942
rect 3514 7440 3570 7449
rect 3514 7375 3570 7384
rect 3528 7177 3556 7375
rect 3712 7256 3740 8366
rect 3620 7228 3740 7256
rect 3514 7168 3570 7177
rect 3514 7103 3570 7112
rect 3528 5914 3556 7103
rect 3620 7002 3648 7228
rect 3698 7168 3754 7177
rect 3698 7103 3754 7112
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3606 6896 3662 6905
rect 3606 6831 3608 6840
rect 3660 6831 3662 6840
rect 3608 6802 3660 6808
rect 3712 6769 3740 7103
rect 3698 6760 3754 6769
rect 3608 6724 3660 6730
rect 3698 6695 3754 6704
rect 3608 6666 3660 6672
rect 3620 6390 3648 6666
rect 3804 6633 3832 10231
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3790 6624 3846 6633
rect 3790 6559 3846 6568
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3620 5914 3648 6122
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3528 3602 3556 4422
rect 3620 3670 3648 5102
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3514 3496 3570 3505
rect 3712 3466 3740 6394
rect 3792 5092 3844 5098
rect 3792 5034 3844 5040
rect 3514 3431 3570 3440
rect 3700 3460 3752 3466
rect 3528 2689 3556 3431
rect 3700 3402 3752 3408
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3514 2680 3570 2689
rect 3514 2615 3570 2624
rect 3712 2514 3740 2790
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3620 1601 3648 2382
rect 3804 2009 3832 5034
rect 3896 4729 3924 9862
rect 3988 9217 4016 10639
rect 4080 10112 4108 10764
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4080 10084 4292 10112
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 3974 9208 4030 9217
rect 3974 9143 4030 9152
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3988 8634 4016 9046
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4080 7993 4108 9959
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4172 9382 4200 9454
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4172 8090 4200 9046
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4066 7984 4122 7993
rect 4066 7919 4122 7928
rect 4068 7404 4120 7410
rect 4120 7364 4200 7392
rect 4068 7346 4120 7352
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3988 7002 4016 7278
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3988 6662 4016 6938
rect 4080 6662 4108 7142
rect 4172 6769 4200 7364
rect 4158 6760 4214 6769
rect 4158 6695 4214 6704
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 4068 6656 4120 6662
rect 4120 6616 4200 6644
rect 4068 6598 4120 6604
rect 3988 6118 4016 6598
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5778 4016 6054
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4080 5681 4108 5782
rect 4066 5672 4122 5681
rect 4172 5642 4200 6616
rect 4264 6458 4292 10084
rect 4540 10062 4568 10406
rect 4632 10266 4660 10950
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4540 9518 4568 9998
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4066 5607 4122 5616
rect 4160 5636 4212 5642
rect 4080 5370 4108 5607
rect 4160 5578 4212 5584
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4264 5250 4292 5646
rect 4080 5234 4292 5250
rect 4068 5228 4292 5234
rect 4120 5222 4292 5228
rect 4068 5170 4120 5176
rect 4356 5148 4384 9386
rect 4540 9178 4568 9454
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4540 8090 4568 8298
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4632 7546 4660 7890
rect 4724 7546 4752 17224
rect 4908 15337 4936 22086
rect 4988 21004 5040 21010
rect 4988 20946 5040 20952
rect 5000 20398 5028 20946
rect 4988 20392 5040 20398
rect 4988 20334 5040 20340
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 5000 16250 5028 16730
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4894 15328 4950 15337
rect 4894 15263 4950 15272
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4816 13394 4844 14554
rect 5092 13870 5120 27520
rect 5448 25492 5500 25498
rect 5448 25434 5500 25440
rect 5172 25424 5224 25430
rect 5172 25366 5224 25372
rect 5184 24954 5212 25366
rect 5172 24948 5224 24954
rect 5172 24890 5224 24896
rect 5460 23338 5488 25434
rect 5644 25226 5672 27520
rect 5632 25220 5684 25226
rect 5632 25162 5684 25168
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6092 24812 6144 24818
rect 6092 24754 6144 24760
rect 6104 24138 6132 24754
rect 6092 24132 6144 24138
rect 6092 24074 6144 24080
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5908 23792 5960 23798
rect 5906 23760 5908 23769
rect 5960 23760 5962 23769
rect 5906 23695 5962 23704
rect 6012 23662 6040 24006
rect 6092 23860 6144 23866
rect 6092 23802 6144 23808
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 5906 23352 5962 23361
rect 5460 23322 5580 23338
rect 5172 23316 5224 23322
rect 5460 23316 5592 23322
rect 5460 23310 5540 23316
rect 5172 23258 5224 23264
rect 5906 23287 5962 23296
rect 5540 23258 5592 23264
rect 5184 22574 5212 23258
rect 5552 22778 5580 23258
rect 5920 23254 5948 23287
rect 5908 23248 5960 23254
rect 5960 23208 6040 23236
rect 5908 23190 5960 23196
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 6012 22778 6040 23208
rect 5540 22772 5592 22778
rect 5460 22732 5540 22760
rect 5172 22568 5224 22574
rect 5172 22510 5224 22516
rect 5264 21344 5316 21350
rect 5264 21286 5316 21292
rect 5276 21078 5304 21286
rect 5460 21146 5488 22732
rect 5540 22714 5592 22720
rect 6000 22772 6052 22778
rect 6000 22714 6052 22720
rect 5540 22160 5592 22166
rect 5540 22102 5592 22108
rect 5552 21690 5580 22102
rect 5632 22024 5684 22030
rect 6104 21978 6132 23802
rect 6196 22556 6224 27520
rect 6460 25220 6512 25226
rect 6460 25162 6512 25168
rect 6274 24712 6330 24721
rect 6274 24647 6330 24656
rect 6288 24206 6316 24647
rect 6368 24336 6420 24342
rect 6368 24278 6420 24284
rect 6276 24200 6328 24206
rect 6276 24142 6328 24148
rect 6288 23866 6316 24142
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 6380 23798 6408 24278
rect 6368 23792 6420 23798
rect 6368 23734 6420 23740
rect 6276 23520 6328 23526
rect 6276 23462 6328 23468
rect 6288 23118 6316 23462
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 6288 22710 6316 23054
rect 6276 22704 6328 22710
rect 6276 22646 6328 22652
rect 6196 22528 6316 22556
rect 6288 21978 6316 22528
rect 5684 21972 6132 21978
rect 5632 21966 6132 21972
rect 5644 21950 6132 21966
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 6000 21344 6052 21350
rect 6104 21332 6132 21950
rect 6052 21304 6132 21332
rect 6196 21950 6316 21978
rect 6000 21286 6052 21292
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 5264 21072 5316 21078
rect 5264 21014 5316 21020
rect 5276 20058 5304 21014
rect 5460 20466 5488 21082
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5172 19984 5224 19990
rect 5172 19926 5224 19932
rect 5184 19514 5212 19926
rect 5448 19780 5500 19786
rect 5448 19722 5500 19728
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5460 19292 5488 19722
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5632 19304 5684 19310
rect 5460 19272 5632 19292
rect 5684 19272 5686 19281
rect 5460 19264 5630 19272
rect 6012 19242 6040 21286
rect 5630 19207 5686 19216
rect 6000 19236 6052 19242
rect 6000 19178 6052 19184
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5460 18970 5488 19110
rect 5448 18964 5500 18970
rect 5368 18924 5448 18952
rect 5368 17814 5396 18924
rect 5448 18906 5500 18912
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6196 18329 6224 21950
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6288 21146 6316 21830
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 6288 20602 6316 21082
rect 6276 20596 6328 20602
rect 6276 20538 6328 20544
rect 6288 20330 6316 20538
rect 6276 20324 6328 20330
rect 6276 20266 6328 20272
rect 6368 18352 6420 18358
rect 6182 18320 6238 18329
rect 6182 18255 6238 18264
rect 6366 18320 6368 18329
rect 6420 18320 6422 18329
rect 6366 18255 6422 18264
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5356 17808 5408 17814
rect 5356 17750 5408 17756
rect 5368 17270 5396 17750
rect 5460 17338 5488 18158
rect 6276 17808 6328 17814
rect 6276 17750 6328 17756
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6288 17338 6316 17750
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 5356 17264 5408 17270
rect 5356 17206 5408 17212
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5264 16176 5316 16182
rect 5262 16144 5264 16153
rect 5316 16144 5318 16153
rect 5262 16079 5318 16088
rect 5368 14278 5396 16390
rect 5460 15570 5488 17138
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5736 16794 5764 16934
rect 6274 16824 6330 16833
rect 5724 16788 5776 16794
rect 6274 16759 6330 16768
rect 5724 16730 5776 16736
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5460 15162 5488 15506
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5460 14482 5488 15098
rect 5552 14550 5580 16390
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5998 16280 6054 16289
rect 5998 16215 6054 16224
rect 6012 16114 6040 16215
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 5828 15638 5856 15914
rect 6012 15706 6040 16050
rect 6196 15910 6224 16662
rect 6184 15904 6236 15910
rect 6182 15872 6184 15881
rect 6236 15872 6238 15881
rect 6182 15807 6238 15816
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 5816 15632 5868 15638
rect 5816 15574 5868 15580
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6012 15162 6040 15506
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6012 14618 6040 15098
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6196 14618 6224 14962
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4816 12986 4844 13330
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 5092 12850 5120 13126
rect 5368 12918 5396 14214
rect 5460 13938 5488 14418
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4816 11830 4844 12174
rect 4804 11824 4856 11830
rect 4802 11792 4804 11801
rect 4856 11792 4858 11801
rect 4802 11727 4858 11736
rect 4802 11656 4858 11665
rect 4802 11591 4858 11600
rect 4816 11286 4844 11591
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4816 10266 4844 11222
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4908 9897 4936 12582
rect 5552 12481 5580 13942
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5538 12472 5594 12481
rect 5448 12436 5500 12442
rect 5538 12407 5594 12416
rect 5448 12378 5500 12384
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5184 11218 5212 11630
rect 5460 11558 5488 12378
rect 6012 12374 6040 13874
rect 6288 13394 6316 16759
rect 6368 16176 6420 16182
rect 6368 16118 6420 16124
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11898 6040 12310
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5552 11354 5580 11562
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5092 10470 5120 11018
rect 5368 10606 5396 11018
rect 5460 10810 5488 11154
rect 6104 11121 6132 13126
rect 6288 12986 6316 13330
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6380 12866 6408 16118
rect 6472 16046 6500 25162
rect 6748 24834 6776 27520
rect 7012 25356 7064 25362
rect 7012 25298 7064 25304
rect 6564 24806 6776 24834
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6458 13968 6514 13977
rect 6458 13903 6514 13912
rect 6288 12838 6408 12866
rect 6472 12850 6500 13903
rect 6460 12844 6512 12850
rect 6090 11112 6146 11121
rect 6090 11047 6146 11056
rect 6000 11008 6052 11014
rect 5998 10976 6000 10985
rect 6052 10976 6054 10985
rect 5622 10908 5918 10928
rect 5998 10911 6054 10920
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5630 10568 5686 10577
rect 5080 10464 5132 10470
rect 5552 10441 5580 10542
rect 5630 10503 5686 10512
rect 5080 10406 5132 10412
rect 5538 10432 5594 10441
rect 4894 9888 4950 9897
rect 4894 9823 4950 9832
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 8430 4936 9318
rect 4986 9208 5042 9217
rect 4986 9143 5042 9152
rect 5000 8673 5028 9143
rect 4986 8664 5042 8673
rect 4986 8599 5042 8608
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4908 7886 4936 8366
rect 4896 7880 4948 7886
rect 4802 7848 4858 7857
rect 4896 7822 4948 7828
rect 4802 7783 4858 7792
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4724 7206 4752 7482
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4816 6089 4844 7783
rect 4908 7342 4936 7822
rect 5092 7732 5120 10406
rect 5538 10367 5594 10376
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5276 9110 5304 9862
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5448 8968 5500 8974
rect 5552 8956 5580 10134
rect 5644 9994 5672 10503
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10305 5764 10406
rect 5722 10296 5778 10305
rect 5722 10231 5778 10240
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5500 8928 5580 8956
rect 5448 8910 5500 8916
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5184 7954 5212 8842
rect 5276 8090 5304 8910
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 8401 5396 8774
rect 5354 8392 5410 8401
rect 5354 8327 5410 8336
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5264 7744 5316 7750
rect 5092 7712 5264 7732
rect 5316 7712 5318 7721
rect 5092 7704 5262 7712
rect 5262 7647 5318 7656
rect 5460 7546 5488 8910
rect 6104 8838 6132 9998
rect 6288 9654 6316 12838
rect 6460 12786 6512 12792
rect 6564 12782 6592 24806
rect 7024 24614 7052 25298
rect 7012 24608 7064 24614
rect 7012 24550 7064 24556
rect 6920 24132 6972 24138
rect 6920 24074 6972 24080
rect 6932 24018 6960 24074
rect 6840 23990 6960 24018
rect 6736 22976 6788 22982
rect 6642 22944 6698 22953
rect 6736 22918 6788 22924
rect 6642 22879 6698 22888
rect 6656 22681 6684 22879
rect 6642 22672 6698 22681
rect 6642 22607 6698 22616
rect 6656 16182 6684 22607
rect 6748 22574 6776 22918
rect 6736 22568 6788 22574
rect 6736 22510 6788 22516
rect 6840 22234 6868 23990
rect 6920 23792 6972 23798
rect 6920 23734 6972 23740
rect 6932 23361 6960 23734
rect 6918 23352 6974 23361
rect 6918 23287 6974 23296
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6748 21010 6776 21830
rect 6826 21448 6882 21457
rect 6826 21383 6882 21392
rect 6840 21350 6868 21383
rect 6932 21350 6960 22714
rect 7024 22642 7052 24550
rect 7104 23724 7156 23730
rect 7104 23666 7156 23672
rect 7116 23186 7144 23666
rect 7196 23656 7248 23662
rect 7196 23598 7248 23604
rect 7104 23180 7156 23186
rect 7104 23122 7156 23128
rect 7116 22778 7144 23122
rect 7208 22778 7236 23598
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 7024 22098 7052 22578
rect 7012 22092 7064 22098
rect 7012 22034 7064 22040
rect 7024 21690 7052 22034
rect 7012 21684 7064 21690
rect 7012 21626 7064 21632
rect 6828 21344 6880 21350
rect 6828 21286 6880 21292
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 6748 20058 6776 20946
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6840 19938 6868 21286
rect 6932 21146 6960 21286
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 6932 20058 6960 21082
rect 7116 20602 7144 22714
rect 7300 22658 7328 27520
rect 7748 25152 7800 25158
rect 7748 25094 7800 25100
rect 7656 24744 7708 24750
rect 7656 24686 7708 24692
rect 7380 24608 7432 24614
rect 7380 24550 7432 24556
rect 7392 23594 7420 24550
rect 7668 24138 7696 24686
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 7380 23588 7432 23594
rect 7380 23530 7432 23536
rect 7472 23588 7524 23594
rect 7472 23530 7524 23536
rect 7484 23322 7512 23530
rect 7656 23520 7708 23526
rect 7656 23462 7708 23468
rect 7472 23316 7524 23322
rect 7472 23258 7524 23264
rect 7668 23225 7696 23462
rect 7654 23216 7710 23225
rect 7380 23180 7432 23186
rect 7654 23151 7710 23160
rect 7380 23122 7432 23128
rect 7392 22710 7420 23122
rect 7208 22630 7328 22658
rect 7380 22704 7432 22710
rect 7380 22646 7432 22652
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6748 19910 6868 19938
rect 6644 16176 6696 16182
rect 6644 16118 6696 16124
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6564 12617 6592 12718
rect 6550 12608 6606 12617
rect 6550 12543 6606 12552
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6380 11286 6408 12242
rect 6458 11384 6514 11393
rect 6458 11319 6460 11328
rect 6512 11319 6514 11328
rect 6460 11290 6512 11296
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 6472 10810 6500 11290
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6656 10248 6684 15982
rect 6748 14906 6776 19910
rect 6932 19310 6960 19994
rect 7116 19922 7144 20538
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 7116 19514 7144 19858
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 7116 18902 7144 19110
rect 7104 18896 7156 18902
rect 7104 18838 7156 18844
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6840 17746 6868 18566
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6840 16658 6868 17070
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6840 16182 6868 16594
rect 6932 16250 6960 18770
rect 7116 18426 7144 18838
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 7024 15162 7052 16934
rect 7116 16114 7144 17070
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7116 15706 7144 16050
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6748 14878 6868 14906
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6748 13841 6776 14758
rect 6734 13832 6790 13841
rect 6734 13767 6736 13776
rect 6788 13767 6790 13776
rect 6736 13738 6788 13744
rect 6748 13530 6776 13738
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6840 13410 6868 14878
rect 6932 13462 6960 15030
rect 6472 10220 6684 10248
rect 6748 13382 6868 13410
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4908 6458 4936 7278
rect 5170 6760 5226 6769
rect 5170 6695 5226 6704
rect 5078 6488 5134 6497
rect 4896 6452 4948 6458
rect 5184 6458 5212 6695
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5078 6423 5134 6432
rect 5172 6452 5224 6458
rect 4896 6394 4948 6400
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4802 6080 4858 6089
rect 4802 6015 4858 6024
rect 4620 5840 4672 5846
rect 4618 5808 4620 5817
rect 4712 5840 4764 5846
rect 4672 5808 4674 5817
rect 4436 5772 4488 5778
rect 4712 5782 4764 5788
rect 4618 5743 4674 5752
rect 4436 5714 4488 5720
rect 4158 5128 4214 5137
rect 4158 5063 4160 5072
rect 4212 5063 4214 5072
rect 4264 5120 4384 5148
rect 4160 5034 4212 5040
rect 3882 4720 3938 4729
rect 3882 4655 3938 4664
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3974 4584 4030 4593
rect 3896 3738 3924 4558
rect 3974 4519 4030 4528
rect 3988 4078 4016 4519
rect 4080 4146 4108 4626
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 4080 3670 4108 3878
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3884 3460 3936 3466
rect 3884 3402 3936 3408
rect 3790 2000 3846 2009
rect 3790 1935 3846 1944
rect 3606 1592 3662 1601
rect 3606 1527 3662 1536
rect 3896 480 3924 3402
rect 3988 2922 4016 3538
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 3988 2582 4016 2858
rect 3976 2576 4028 2582
rect 3976 2518 4028 2524
rect 4080 1714 4108 3606
rect 4172 3369 4200 3878
rect 4264 3466 4292 5120
rect 4448 5030 4476 5714
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4010 4384 4422
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 4158 3360 4214 3369
rect 4158 3295 4214 3304
rect 3988 1686 4108 1714
rect 3988 1193 4016 1686
rect 4066 1456 4122 1465
rect 4066 1391 4122 1400
rect 3974 1184 4030 1193
rect 3974 1119 4030 1128
rect 202 0 258 480
rect 662 0 718 480
rect 1214 0 1270 480
rect 1766 0 1822 480
rect 2318 0 2374 480
rect 2870 0 2926 480
rect 3422 0 3478 480
rect 3882 0 3938 480
rect 4080 377 4108 1391
rect 4172 785 4200 3295
rect 4356 2854 4384 3946
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4356 2582 4384 2790
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 4158 776 4214 785
rect 4158 711 4214 720
rect 4448 480 4476 4966
rect 4540 1873 4568 5306
rect 4632 5302 4660 5743
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4724 5166 4752 5782
rect 4712 5160 4764 5166
rect 4618 5128 4674 5137
rect 4712 5102 4764 5108
rect 4618 5063 4674 5072
rect 4632 4826 4660 5063
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4632 4282 4660 4762
rect 4724 4758 4752 5102
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4816 4554 4844 6015
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4632 3097 4660 3606
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4618 3088 4674 3097
rect 4618 3023 4674 3032
rect 4526 1864 4582 1873
rect 4526 1799 4582 1808
rect 4632 1057 4660 3023
rect 4724 2310 4752 3470
rect 4908 2650 4936 6190
rect 5092 6186 5120 6423
rect 5172 6394 5224 6400
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 5092 6089 5120 6122
rect 5078 6080 5134 6089
rect 5078 6015 5134 6024
rect 5092 5914 5120 6015
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5460 5778 5488 6598
rect 5552 6322 5580 8502
rect 6104 8498 6132 8774
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6288 7698 6316 9590
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6012 7670 6316 7698
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5552 5914 5580 6258
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 5092 2666 5120 5238
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5460 5030 5488 5170
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5460 4729 5488 4966
rect 5552 4826 5580 5510
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5446 4720 5502 4729
rect 5446 4655 5502 4664
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5446 4312 5502 4321
rect 5622 4304 5918 4324
rect 5502 4270 5580 4298
rect 5446 4247 5502 4256
rect 5552 4010 5580 4270
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5000 2638 5120 2666
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 4618 1048 4674 1057
rect 4618 983 4674 992
rect 5000 480 5028 2638
rect 5356 2372 5408 2378
rect 5356 2314 5408 2320
rect 5368 2281 5396 2314
rect 5354 2272 5410 2281
rect 5354 2207 5410 2216
rect 5552 480 5580 3674
rect 5644 3466 5672 3878
rect 5736 3641 5764 4082
rect 6012 3738 6040 7670
rect 6182 7576 6238 7585
rect 6182 7511 6238 7520
rect 6276 7540 6328 7546
rect 6196 7478 6224 7511
rect 6276 7482 6328 7488
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6104 7002 6132 7346
rect 6196 7342 6224 7373
rect 6184 7336 6236 7342
rect 6288 7290 6316 7482
rect 6380 7324 6408 9046
rect 6472 7478 6500 10220
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6656 9897 6684 10066
rect 6642 9888 6698 9897
rect 6642 9823 6698 9832
rect 6748 9110 6776 13382
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6932 12442 6960 12854
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6932 11694 6960 12038
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6932 10470 6960 11018
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6840 9654 6868 9930
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6460 7472 6512 7478
rect 6460 7414 6512 7420
rect 6656 7410 6684 8570
rect 6748 7818 6776 8774
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6840 7546 6868 8978
rect 6932 8838 6960 9386
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8242 6960 8774
rect 7024 8430 7052 13126
rect 7104 12368 7156 12374
rect 7104 12310 7156 12316
rect 7116 8616 7144 12310
rect 7208 9353 7236 22630
rect 7760 22506 7788 25094
rect 7748 22500 7800 22506
rect 7748 22442 7800 22448
rect 7760 22234 7788 22442
rect 7748 22228 7800 22234
rect 7748 22170 7800 22176
rect 7380 22024 7432 22030
rect 7852 22012 7880 27520
rect 7932 25220 7984 25226
rect 7932 25162 7984 25168
rect 7944 24750 7972 25162
rect 8404 24834 8432 27520
rect 8576 25424 8628 25430
rect 8576 25366 8628 25372
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8496 24886 8524 25230
rect 8036 24806 8432 24834
rect 8484 24880 8536 24886
rect 8484 24822 8536 24828
rect 7932 24744 7984 24750
rect 7932 24686 7984 24692
rect 7944 24410 7972 24686
rect 7932 24404 7984 24410
rect 7932 24346 7984 24352
rect 7380 21966 7432 21972
rect 7484 21984 7880 22012
rect 7392 21486 7420 21966
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7392 20806 7420 21422
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7392 19922 7420 20742
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7392 18290 7420 18702
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7392 17882 7420 18226
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7392 16998 7420 17818
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 16726 7420 16934
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 7484 16538 7512 21984
rect 7748 21616 7800 21622
rect 7748 21558 7800 21564
rect 7760 21078 7788 21558
rect 7748 21072 7800 21078
rect 7748 21014 7800 21020
rect 7562 20632 7618 20641
rect 7562 20567 7618 20576
rect 7576 19360 7604 20567
rect 7576 19332 7788 19360
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 7576 18970 7604 19178
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7576 17814 7604 18906
rect 7564 17808 7616 17814
rect 7564 17750 7616 17756
rect 7654 17640 7710 17649
rect 7654 17575 7656 17584
rect 7708 17575 7710 17584
rect 7656 17546 7708 17552
rect 7760 16572 7788 19332
rect 7932 18352 7984 18358
rect 7932 18294 7984 18300
rect 7944 17814 7972 18294
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 7930 17368 7986 17377
rect 7930 17303 7986 17312
rect 7760 16544 7880 16572
rect 7300 16510 7512 16538
rect 7300 11914 7328 16510
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7392 16017 7420 16390
rect 7378 16008 7434 16017
rect 7378 15943 7380 15952
rect 7432 15943 7434 15952
rect 7380 15914 7432 15920
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 7484 15094 7512 15574
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7392 14550 7420 14758
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 7668 14482 7696 15302
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7470 13560 7526 13569
rect 7470 13495 7472 13504
rect 7524 13495 7526 13504
rect 7472 13466 7524 13472
rect 7378 13016 7434 13025
rect 7378 12951 7434 12960
rect 7392 12850 7420 12951
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7484 12442 7512 13466
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7300 11886 7512 11914
rect 7378 11792 7434 11801
rect 7378 11727 7434 11736
rect 7392 11014 7420 11727
rect 7380 11008 7432 11014
rect 7300 10968 7380 10996
rect 7300 10606 7328 10968
rect 7380 10950 7432 10956
rect 7484 10849 7512 11886
rect 7470 10840 7526 10849
rect 7470 10775 7526 10784
rect 7576 10690 7604 13126
rect 7746 10840 7802 10849
rect 7746 10775 7802 10784
rect 7392 10662 7604 10690
rect 7656 10668 7708 10674
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7194 9344 7250 9353
rect 7194 9279 7250 9288
rect 7286 8664 7342 8673
rect 7116 8588 7236 8616
rect 7286 8599 7342 8608
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6932 8214 7052 8242
rect 7024 8129 7052 8214
rect 7010 8120 7066 8129
rect 7010 8055 7066 8064
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 7024 7342 7052 7686
rect 7116 7546 7144 8434
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7208 7426 7236 8588
rect 7300 8498 7328 8599
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7286 8120 7342 8129
rect 7286 8055 7342 8064
rect 7300 7721 7328 8055
rect 7286 7712 7342 7721
rect 7286 7647 7342 7656
rect 7116 7398 7236 7426
rect 7012 7336 7064 7342
rect 6380 7296 6500 7324
rect 6236 7284 6316 7290
rect 6184 7278 6316 7284
rect 6196 7262 6316 7278
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6196 5896 6224 7262
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6104 5868 6224 5896
rect 6104 5574 6132 5868
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6090 5400 6146 5409
rect 6090 5335 6146 5344
rect 6104 5166 6132 5335
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 6104 3670 6132 4966
rect 6196 4826 6224 5714
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6288 4706 6316 7142
rect 6366 6352 6422 6361
rect 6366 6287 6422 6296
rect 6196 4678 6316 4706
rect 6196 3777 6224 4678
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 6182 3768 6238 3777
rect 6182 3703 6238 3712
rect 6092 3664 6144 3670
rect 5722 3632 5778 3641
rect 6092 3606 6144 3612
rect 5722 3567 5778 3576
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6104 3194 6132 3606
rect 6184 3460 6236 3466
rect 6184 3402 6236 3408
rect 6196 3233 6224 3402
rect 6182 3224 6238 3233
rect 6092 3188 6144 3194
rect 6182 3159 6238 3168
rect 6092 3130 6144 3136
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 6012 2281 6040 2314
rect 5998 2272 6054 2281
rect 5622 2204 5918 2224
rect 5998 2207 6054 2216
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6090 1592 6146 1601
rect 6090 1527 6146 1536
rect 6104 480 6132 1527
rect 6288 1329 6316 3946
rect 6380 3398 6408 6287
rect 6472 6118 6500 7296
rect 7012 7278 7064 7284
rect 7116 7274 7144 7398
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7010 7032 7066 7041
rect 7010 6967 7066 6976
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6840 6186 6868 6802
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 6225 6960 6598
rect 6918 6216 6974 6225
rect 6828 6180 6880 6186
rect 6918 6151 6974 6160
rect 6828 6122 6880 6128
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6564 4214 6592 4626
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6472 4078 6500 4109
rect 6460 4072 6512 4078
rect 6458 4040 6460 4049
rect 6512 4040 6514 4049
rect 6458 3975 6514 3984
rect 6472 3738 6500 3975
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6564 2990 6592 3470
rect 6552 2984 6604 2990
rect 6550 2952 6552 2961
rect 6604 2952 6606 2961
rect 6550 2887 6606 2896
rect 6274 1320 6330 1329
rect 6274 1255 6330 1264
rect 6656 480 6684 6054
rect 6840 5817 6868 6122
rect 6826 5808 6882 5817
rect 6826 5743 6882 5752
rect 6734 5400 6790 5409
rect 6734 5335 6790 5344
rect 6748 5098 6776 5335
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6840 4758 6868 5743
rect 7024 5370 7052 6967
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7116 5250 7144 7210
rect 7300 6882 7328 7647
rect 7392 7177 7420 10662
rect 7656 10610 7708 10616
rect 7668 10266 7696 10610
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7484 7750 7512 10202
rect 7654 9752 7710 9761
rect 7760 9738 7788 10775
rect 7710 9710 7788 9738
rect 7654 9687 7710 9696
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7576 9042 7604 9386
rect 7654 9344 7710 9353
rect 7654 9279 7710 9288
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7576 8634 7604 8978
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7562 8256 7618 8265
rect 7562 8191 7618 8200
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 7410 7512 7686
rect 7576 7478 7604 8191
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7378 7168 7434 7177
rect 7378 7103 7434 7112
rect 7392 7002 7420 7103
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7300 6854 7512 6882
rect 7378 6352 7434 6361
rect 7378 6287 7434 6296
rect 7194 6216 7250 6225
rect 7392 6186 7420 6287
rect 7194 6151 7196 6160
rect 7248 6151 7250 6160
rect 7380 6180 7432 6186
rect 7196 6122 7248 6128
rect 7380 6122 7432 6128
rect 7024 5222 7144 5250
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6748 3602 6776 4422
rect 6840 4282 6868 4694
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 7024 3210 7052 5222
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7116 3913 7144 3946
rect 7102 3904 7158 3913
rect 7102 3839 7158 3848
rect 7208 3398 7236 6122
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7300 5953 7328 6054
rect 7286 5944 7342 5953
rect 7286 5879 7288 5888
rect 7340 5879 7342 5888
rect 7288 5850 7340 5856
rect 7300 5370 7328 5850
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7300 3670 7328 4150
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7024 3182 7236 3210
rect 7300 3194 7328 3606
rect 7392 3466 7420 4082
rect 7484 3534 7512 6854
rect 7668 5098 7696 9279
rect 7760 6254 7788 9710
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7852 5794 7880 16544
rect 7944 12374 7972 17303
rect 8036 16833 8064 24806
rect 8496 24342 8524 24822
rect 8588 24614 8616 25366
rect 8576 24608 8628 24614
rect 8576 24550 8628 24556
rect 8116 24336 8168 24342
rect 8116 24278 8168 24284
rect 8484 24336 8536 24342
rect 8484 24278 8536 24284
rect 8128 23526 8156 24278
rect 8300 24200 8352 24206
rect 8300 24142 8352 24148
rect 8312 23866 8340 24142
rect 8300 23860 8352 23866
rect 8300 23802 8352 23808
rect 8496 23610 8524 24278
rect 8404 23582 8524 23610
rect 8116 23520 8168 23526
rect 8116 23462 8168 23468
rect 8404 23202 8432 23582
rect 8116 23180 8168 23186
rect 8116 23122 8168 23128
rect 8312 23174 8432 23202
rect 8128 23066 8156 23122
rect 8312 23066 8340 23174
rect 8128 23038 8340 23066
rect 8128 22098 8156 23038
rect 8588 22817 8616 24550
rect 8668 24404 8720 24410
rect 8668 24346 8720 24352
rect 8680 23662 8708 24346
rect 8668 23656 8720 23662
rect 8668 23598 8720 23604
rect 8680 23322 8708 23598
rect 8668 23316 8720 23322
rect 8668 23258 8720 23264
rect 8574 22808 8630 22817
rect 8680 22778 8708 23258
rect 8574 22743 8630 22752
rect 8668 22772 8720 22778
rect 8668 22714 8720 22720
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 8220 21690 8248 22102
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8312 20602 8340 20878
rect 8956 20777 8984 27520
rect 9508 23905 9536 27520
rect 10060 24698 10088 27520
rect 10612 25786 10640 27520
rect 10612 25758 10732 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 9864 24676 9916 24682
rect 10060 24670 10180 24698
rect 9864 24618 9916 24624
rect 9876 24410 9904 24618
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9864 24404 9916 24410
rect 9864 24346 9916 24352
rect 9678 24304 9734 24313
rect 9678 24239 9734 24248
rect 9494 23896 9550 23905
rect 9494 23831 9550 23840
rect 9218 23080 9274 23089
rect 9218 23015 9274 23024
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 9126 21856 9182 21865
rect 9048 21350 9076 21830
rect 9126 21791 9182 21800
rect 9140 21690 9168 21791
rect 9128 21684 9180 21690
rect 9128 21626 9180 21632
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 9048 20874 9076 21286
rect 9036 20868 9088 20874
rect 9036 20810 9088 20816
rect 8942 20768 8998 20777
rect 8942 20703 8998 20712
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8220 19922 8248 20198
rect 8312 20058 8340 20538
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 8220 19378 8248 19858
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 8220 19242 8248 19314
rect 9036 19304 9088 19310
rect 9036 19246 9088 19252
rect 8208 19236 8260 19242
rect 8208 19178 8260 19184
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8022 16824 8078 16833
rect 8022 16759 8078 16768
rect 8128 15722 8156 18158
rect 8772 17921 8800 19110
rect 9048 18970 9076 19246
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 9232 18601 9260 23015
rect 9692 22658 9720 24239
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9784 22778 9812 23462
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9692 22630 9812 22658
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9416 21418 9444 21830
rect 9404 21412 9456 21418
rect 9404 21354 9456 21360
rect 9416 20602 9444 21354
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 9600 20312 9628 20742
rect 9680 20324 9732 20330
rect 9600 20284 9680 20312
rect 9680 20266 9732 20272
rect 9496 20256 9548 20262
rect 9496 20198 9548 20204
rect 9508 19718 9536 20198
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9692 19514 9720 20266
rect 9784 19938 9812 22630
rect 9876 22098 9904 24346
rect 9968 22574 9996 24550
rect 10046 23352 10102 23361
rect 10046 23287 10048 23296
rect 10100 23287 10102 23296
rect 10048 23258 10100 23264
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 10060 22778 10088 23122
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 9956 22568 10008 22574
rect 9956 22510 10008 22516
rect 9968 22234 9996 22510
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 10060 21146 10088 21422
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9968 20466 9996 20946
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9968 20058 9996 20402
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9784 19910 9996 19938
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9784 19378 9812 19790
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9218 18592 9274 18601
rect 9218 18527 9274 18536
rect 9232 18290 9260 18527
rect 9310 18456 9366 18465
rect 9310 18391 9366 18400
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 8758 17912 8814 17921
rect 9232 17882 9260 18226
rect 8758 17847 8814 17856
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8220 17338 8248 17614
rect 9140 17338 9168 17682
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 8220 16794 8248 17274
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8036 15694 8248 15722
rect 8036 15570 8064 15694
rect 8116 15632 8168 15638
rect 8116 15574 8168 15580
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 8036 15026 8064 15302
rect 8128 15162 8156 15574
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 8220 13818 8248 15694
rect 8680 15638 8708 16050
rect 8772 16046 8800 16730
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8772 15706 8800 15982
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8668 15632 8720 15638
rect 8298 15600 8354 15609
rect 8668 15574 8720 15580
rect 8298 15535 8300 15544
rect 8352 15535 8354 15544
rect 8300 15506 8352 15512
rect 8312 15162 8340 15506
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8772 15337 8800 15438
rect 8758 15328 8814 15337
rect 8758 15263 8814 15272
rect 9324 15178 9352 18391
rect 9588 18352 9640 18358
rect 9588 18294 9640 18300
rect 9402 17912 9458 17921
rect 9402 17847 9458 17856
rect 9416 16590 9444 17847
rect 9494 17096 9550 17105
rect 9494 17031 9550 17040
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 9232 15150 9352 15178
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 8404 14618 8432 14826
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8220 13790 8340 13818
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8220 13326 8248 13670
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8220 12986 8248 13262
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8116 12708 8168 12714
rect 8116 12650 8168 12656
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 8036 12186 8064 12582
rect 8128 12306 8156 12650
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 7944 12158 8064 12186
rect 7944 7206 7972 12158
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 10441 8064 12038
rect 8128 11898 8156 12242
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8220 11694 8248 12922
rect 8312 12170 8340 13790
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8220 11354 8248 11630
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8312 10742 8340 12106
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8312 10470 8340 10542
rect 8300 10464 8352 10470
rect 8022 10432 8078 10441
rect 8300 10406 8352 10412
rect 8022 10367 8078 10376
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 8036 6633 8064 10367
rect 8312 9178 8340 10406
rect 8390 9616 8446 9625
rect 8390 9551 8446 9560
rect 8404 9518 8432 9551
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8128 7886 8156 8774
rect 8312 8650 8340 9114
rect 8220 8634 8340 8650
rect 8208 8628 8340 8634
rect 8260 8622 8340 8628
rect 8208 8570 8260 8576
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8312 8106 8340 8502
rect 8220 8078 8340 8106
rect 8220 7954 8248 8078
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7546 8156 7822
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8220 7002 8248 7890
rect 8312 7546 8340 7958
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8404 7313 8432 9318
rect 8496 8498 8524 13126
rect 9048 12646 9076 14758
rect 9140 13308 9168 15030
rect 9232 14929 9260 15150
rect 9218 14920 9274 14929
rect 9218 14855 9274 14864
rect 9232 13444 9260 14855
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9416 14278 9444 14758
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9416 13841 9444 14214
rect 9402 13832 9458 13841
rect 9402 13767 9458 13776
rect 9508 13546 9536 17031
rect 9600 13705 9628 18294
rect 9784 18272 9812 19110
rect 9876 18698 9904 19654
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9784 18244 9904 18272
rect 9770 18184 9826 18193
rect 9680 18148 9732 18154
rect 9770 18119 9826 18128
rect 9680 18090 9732 18096
rect 9692 16969 9720 18090
rect 9784 18086 9812 18119
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9678 16960 9734 16969
rect 9678 16895 9734 16904
rect 9586 13696 9642 13705
rect 9586 13631 9642 13640
rect 9508 13518 9628 13546
rect 9232 13416 9536 13444
rect 9140 13280 9352 13308
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 8668 12232 8720 12238
rect 9048 12209 9076 12310
rect 9128 12232 9180 12238
rect 8668 12174 8720 12180
rect 9034 12200 9090 12209
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8588 11150 8616 12038
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8574 10840 8630 10849
rect 8574 10775 8630 10784
rect 8588 10062 8616 10775
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 9178 8616 9998
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8390 7304 8446 7313
rect 8390 7239 8446 7248
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8300 6792 8352 6798
rect 8298 6760 8300 6769
rect 8352 6760 8354 6769
rect 8298 6695 8354 6704
rect 8392 6656 8444 6662
rect 8022 6624 8078 6633
rect 8392 6598 8444 6604
rect 8022 6559 8078 6568
rect 8024 6384 8076 6390
rect 8024 6326 8076 6332
rect 7760 5766 7880 5794
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7760 4434 7788 5766
rect 8036 5681 8064 6326
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 7838 5672 7894 5681
rect 7838 5607 7840 5616
rect 7892 5607 7894 5616
rect 8022 5672 8078 5681
rect 8022 5607 8078 5616
rect 7840 5578 7892 5584
rect 7668 4406 7788 4434
rect 7668 3777 7696 4406
rect 8220 3942 8248 6258
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8208 3936 8260 3942
rect 8312 3913 8340 5510
rect 8208 3878 8260 3884
rect 8298 3904 8354 3913
rect 8298 3839 8354 3848
rect 7654 3768 7710 3777
rect 7654 3703 7710 3712
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7208 480 7236 3182
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7300 2650 7328 3130
rect 7392 2990 7420 3402
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7668 480 7696 3703
rect 8206 3632 8262 3641
rect 7840 3596 7892 3602
rect 8206 3567 8262 3576
rect 7840 3538 7892 3544
rect 7852 3505 7880 3538
rect 7838 3496 7894 3505
rect 7838 3431 7894 3440
rect 7852 2990 7880 3431
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 8220 480 8248 3567
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 8312 2650 8340 3402
rect 8404 2689 8432 6598
rect 8588 6458 8616 8570
rect 8680 8430 8708 12174
rect 9324 12209 9352 13280
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 9128 12174 9180 12180
rect 9310 12200 9366 12209
rect 9034 12135 9090 12144
rect 9048 11830 9076 12135
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8772 10062 8800 10950
rect 8944 10804 8996 10810
rect 9048 10792 9076 11222
rect 8996 10764 9076 10792
rect 8944 10746 8996 10752
rect 9048 10266 9076 10764
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9034 10160 9090 10169
rect 9034 10095 9090 10104
rect 9048 10062 9076 10095
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 8772 9926 8800 9998
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8772 9586 8800 9862
rect 9048 9722 9076 9998
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8852 8492 8904 8498
rect 8844 8440 8852 8480
rect 8844 8434 8904 8440
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8680 8090 8708 8366
rect 8844 8344 8872 8434
rect 8956 8362 8984 8978
rect 8944 8356 8996 8362
rect 8844 8316 8892 8344
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8864 6934 8892 8316
rect 8944 8298 8996 8304
rect 8956 8090 8984 8298
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8852 6928 8904 6934
rect 8758 6896 8814 6905
rect 8852 6870 8904 6876
rect 8758 6831 8814 6840
rect 9036 6860 9088 6866
rect 8576 6452 8628 6458
rect 8496 6412 8576 6440
rect 8496 5370 8524 6412
rect 8576 6394 8628 6400
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8496 3194 8524 3674
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8588 2825 8616 5510
rect 8772 5098 8800 6831
rect 9036 6802 9088 6808
rect 9048 5574 9076 6802
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8680 4026 8708 4966
rect 8772 4826 8800 5034
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8680 3998 8800 4026
rect 8956 4010 8984 4422
rect 8574 2816 8630 2825
rect 8574 2751 8630 2760
rect 8390 2680 8446 2689
rect 8300 2644 8352 2650
rect 8390 2615 8446 2624
rect 8300 2586 8352 2592
rect 8772 480 8800 3998
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 8956 3738 8984 3946
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9048 3505 9076 5510
rect 9140 5030 9168 12174
rect 9220 12164 9272 12170
rect 9310 12135 9366 12144
rect 9220 12106 9272 12112
rect 9232 11354 9260 12106
rect 9416 12102 9444 12650
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9508 11898 9536 13416
rect 9600 12238 9628 13518
rect 9784 12594 9812 17138
rect 9876 16946 9904 18244
rect 9968 17377 9996 19910
rect 10048 19236 10100 19242
rect 10048 19178 10100 19184
rect 10060 18834 10088 19178
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 10060 17882 10088 18770
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 9954 17368 10010 17377
rect 9954 17303 10010 17312
rect 10152 17202 10180 24670
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10612 23866 10640 24142
rect 10600 23860 10652 23866
rect 10600 23802 10652 23808
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10598 23216 10654 23225
rect 10598 23151 10654 23160
rect 10612 23050 10640 23151
rect 10600 23044 10652 23050
rect 10600 22986 10652 22992
rect 10704 22545 10732 25758
rect 11060 25356 11112 25362
rect 11060 25298 11112 25304
rect 10784 25152 10836 25158
rect 10784 25094 10836 25100
rect 10968 25152 11020 25158
rect 10968 25094 11020 25100
rect 10796 24614 10824 25094
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 10784 24608 10836 24614
rect 10784 24550 10836 24556
rect 10796 23610 10824 24550
rect 10888 23730 10916 24754
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 10796 23582 10916 23610
rect 10690 22536 10746 22545
rect 10690 22471 10746 22480
rect 10692 22432 10744 22438
rect 10692 22374 10744 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10508 22092 10560 22098
rect 10508 22034 10560 22040
rect 10520 21554 10548 22034
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10612 21332 10640 21966
rect 10704 21690 10732 22374
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10692 21344 10744 21350
rect 10612 21304 10692 21332
rect 10692 21286 10744 21292
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10704 21078 10732 21286
rect 10796 21146 10824 22034
rect 10888 22001 10916 23582
rect 10874 21992 10930 22001
rect 10874 21927 10930 21936
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10692 21072 10744 21078
rect 10692 21014 10744 21020
rect 10704 20262 10732 21014
rect 10782 20360 10838 20369
rect 10782 20295 10838 20304
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10796 20058 10824 20295
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10232 19984 10284 19990
rect 10232 19926 10284 19932
rect 10244 19242 10272 19926
rect 10598 19816 10654 19825
rect 10598 19751 10654 19760
rect 10612 19310 10640 19751
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10692 18896 10744 18902
rect 10692 18838 10744 18844
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10244 18154 10272 18702
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 10244 17082 10272 17750
rect 10704 17542 10732 18838
rect 10888 18442 10916 21830
rect 10980 21332 11008 25094
rect 11072 24614 11100 25298
rect 11164 24834 11192 27520
rect 11520 25424 11572 25430
rect 11520 25366 11572 25372
rect 11426 24848 11482 24857
rect 11164 24806 11376 24834
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 11072 24313 11100 24550
rect 11152 24336 11204 24342
rect 11058 24304 11114 24313
rect 11152 24278 11204 24284
rect 11058 24239 11114 24248
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 11072 23118 11100 23530
rect 11164 23526 11192 24278
rect 11152 23520 11204 23526
rect 11152 23462 11204 23468
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11072 22778 11100 23054
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 11348 21434 11376 24806
rect 11426 24783 11482 24792
rect 11440 21894 11468 24783
rect 11532 24614 11560 25366
rect 11520 24608 11572 24614
rect 11520 24550 11572 24556
rect 11532 23361 11560 24550
rect 11518 23352 11574 23361
rect 11518 23287 11574 23296
rect 11532 22137 11560 23287
rect 11518 22128 11574 22137
rect 11518 22063 11574 22072
rect 11428 21888 11480 21894
rect 11428 21830 11480 21836
rect 11244 21412 11296 21418
rect 11348 21406 11652 21434
rect 11244 21354 11296 21360
rect 11060 21344 11112 21350
rect 10980 21304 11060 21332
rect 10980 20602 11008 21304
rect 11060 21286 11112 21292
rect 11256 20602 11284 21354
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11348 20505 11376 21286
rect 11518 20768 11574 20777
rect 11518 20703 11574 20712
rect 11334 20496 11390 20505
rect 11334 20431 11390 20440
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11072 19174 11100 19994
rect 11256 19922 11284 20198
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11256 19310 11284 19858
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 11060 19168 11112 19174
rect 11164 19145 11192 19178
rect 11060 19110 11112 19116
rect 11150 19136 11206 19145
rect 11150 19071 11206 19080
rect 11244 18896 11296 18902
rect 11242 18864 11244 18873
rect 11296 18864 11298 18873
rect 11242 18799 11298 18808
rect 11348 18748 11376 20431
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 11440 19825 11468 19858
rect 11426 19816 11482 19825
rect 11426 19751 11482 19760
rect 11428 19236 11480 19242
rect 11428 19178 11480 19184
rect 11440 18970 11468 19178
rect 11428 18964 11480 18970
rect 11428 18906 11480 18912
rect 10796 18414 10916 18442
rect 11256 18720 11376 18748
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10152 17054 10272 17082
rect 10152 16998 10180 17054
rect 10140 16992 10192 16998
rect 10046 16960 10102 16969
rect 9876 16918 9996 16946
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9876 15366 9904 16730
rect 9968 15994 9996 16918
rect 10140 16934 10192 16940
rect 10046 16895 10102 16904
rect 10060 16726 10088 16895
rect 10048 16720 10100 16726
rect 10152 16697 10180 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10048 16662 10100 16668
rect 10138 16688 10194 16697
rect 10060 16250 10088 16662
rect 10138 16623 10194 16632
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10612 16182 10640 16526
rect 10600 16176 10652 16182
rect 10600 16118 10652 16124
rect 9968 15966 10180 15994
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9968 15570 9996 15846
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9876 14498 9904 15302
rect 9968 15162 9996 15506
rect 9956 15156 10008 15162
rect 10008 15116 10088 15144
rect 9956 15098 10008 15104
rect 9956 14884 10008 14890
rect 9956 14826 10008 14832
rect 9968 14618 9996 14826
rect 10060 14618 10088 15116
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 9876 14482 9996 14498
rect 9876 14476 10008 14482
rect 9876 14470 9956 14476
rect 9956 14418 10008 14424
rect 9968 14074 9996 14418
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9968 13530 9996 14010
rect 10152 13977 10180 15966
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10324 15632 10376 15638
rect 10324 15574 10376 15580
rect 10336 15162 10364 15574
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10612 14074 10640 14350
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10138 13968 10194 13977
rect 10138 13903 10194 13912
rect 10138 13696 10194 13705
rect 10138 13631 10194 13640
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9968 12850 9996 13466
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9956 12640 10008 12646
rect 9784 12566 9904 12594
rect 9956 12582 10008 12588
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9600 11218 9628 12038
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9692 11286 9720 11766
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9600 10266 9628 11154
rect 9692 10266 9720 11222
rect 9770 11112 9826 11121
rect 9770 11047 9772 11056
rect 9824 11047 9826 11056
rect 9772 11018 9824 11024
rect 9876 10985 9904 12566
rect 9968 11393 9996 12582
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10060 11898 10088 12242
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9954 11384 10010 11393
rect 9954 11319 10010 11328
rect 10060 11014 10088 11698
rect 10152 11626 10180 13631
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10336 12986 10364 13126
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12424 10732 17478
rect 10796 17218 10824 18414
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 10888 17921 10916 18294
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10874 17912 10930 17921
rect 10874 17847 10930 17856
rect 10980 17338 11008 18226
rect 11256 17678 11284 18720
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11348 18290 11376 18566
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11348 17882 11376 18022
rect 11336 17876 11388 17882
rect 11336 17818 11388 17824
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 11256 17270 11284 17614
rect 11244 17264 11296 17270
rect 10796 17190 11008 17218
rect 11244 17206 11296 17212
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10888 16794 10916 16934
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10782 14240 10838 14249
rect 10782 14175 10838 14184
rect 10796 12986 10824 14175
rect 10876 14000 10928 14006
rect 10874 13968 10876 13977
rect 10928 13968 10930 13977
rect 10874 13903 10930 13912
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10888 12918 10916 13466
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 10704 12396 10916 12424
rect 10690 12336 10746 12345
rect 10690 12271 10692 12280
rect 10744 12271 10746 12280
rect 10692 12242 10744 12248
rect 10704 11898 10732 12242
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10140 11620 10192 11626
rect 10140 11562 10192 11568
rect 10152 11354 10180 11562
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10796 11354 10824 12106
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10048 11008 10100 11014
rect 9862 10976 9918 10985
rect 10048 10950 10100 10956
rect 9862 10911 9918 10920
rect 10060 10810 10088 10950
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10796 10470 10824 11086
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 9862 10024 9918 10033
rect 9862 9959 9918 9968
rect 9218 9888 9274 9897
rect 9218 9823 9274 9832
rect 9232 7732 9260 9823
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9508 9178 9536 9522
rect 9678 9480 9734 9489
rect 9678 9415 9734 9424
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9692 9042 9720 9415
rect 9876 9178 9904 9959
rect 10520 9722 10548 10066
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9680 8560 9732 8566
rect 9310 8528 9366 8537
rect 9310 8463 9312 8472
rect 9364 8463 9366 8472
rect 9494 8528 9550 8537
rect 9680 8502 9732 8508
rect 9494 8463 9550 8472
rect 9312 8434 9364 8440
rect 9508 8430 9536 8463
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9692 8106 9720 8502
rect 9770 8392 9826 8401
rect 9770 8327 9826 8336
rect 9600 8078 9720 8106
rect 9600 8022 9628 8078
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9784 7954 9812 8327
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9312 7744 9364 7750
rect 9232 7704 9312 7732
rect 9312 7686 9364 7692
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9034 3496 9090 3505
rect 9034 3431 9090 3440
rect 9324 3369 9352 7686
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9494 7304 9550 7313
rect 9494 7239 9496 7248
rect 9548 7239 9550 7248
rect 9496 7210 9548 7216
rect 9508 7002 9536 7210
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9508 5914 9536 6666
rect 9600 6474 9628 7414
rect 9784 7002 9812 7890
rect 9876 7206 9904 8230
rect 10060 8090 10088 8978
rect 10152 8265 10180 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10704 9178 10732 10134
rect 10796 10062 10824 10406
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10796 9722 10824 9998
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10888 9450 10916 12396
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10520 8498 10548 8774
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10336 8401 10364 8434
rect 10322 8392 10378 8401
rect 10322 8327 10378 8336
rect 10138 8256 10194 8265
rect 10138 8191 10194 8200
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9600 6458 9720 6474
rect 9600 6452 9732 6458
rect 9600 6446 9680 6452
rect 9680 6394 9732 6400
rect 9680 6112 9732 6118
rect 9600 6060 9680 6066
rect 9600 6054 9732 6060
rect 9600 6038 9720 6054
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9600 5098 9628 6038
rect 9770 5808 9826 5817
rect 9680 5772 9732 5778
rect 9954 5808 10010 5817
rect 9826 5766 9904 5794
rect 9770 5743 9826 5752
rect 9680 5714 9732 5720
rect 9692 5681 9720 5714
rect 9678 5672 9734 5681
rect 9678 5607 9734 5616
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9588 5092 9640 5098
rect 9588 5034 9640 5040
rect 9784 4554 9812 5510
rect 9876 5370 9904 5766
rect 9954 5743 9956 5752
rect 10008 5743 10010 5752
rect 9956 5714 10008 5720
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9678 3904 9734 3913
rect 9310 3360 9366 3369
rect 9310 3295 9366 3304
rect 9310 3088 9366 3097
rect 9310 3023 9366 3032
rect 9324 480 9352 3023
rect 9508 2854 9536 3878
rect 9678 3839 9734 3848
rect 9692 3602 9720 3839
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9508 2650 9536 2790
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9692 921 9720 3334
rect 9784 2582 9812 4490
rect 9876 4078 9904 4558
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9876 3670 9904 4014
rect 9968 3738 9996 4626
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9968 1034 9996 2858
rect 10060 2553 10088 7822
rect 10784 7472 10836 7478
rect 10782 7440 10784 7449
rect 10836 7440 10838 7449
rect 10782 7375 10838 7384
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10704 7177 10732 7210
rect 10690 7168 10746 7177
rect 10289 7100 10585 7120
rect 10690 7103 10746 7112
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10888 6186 10916 8570
rect 10980 8294 11008 17190
rect 11440 17066 11468 17614
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 11428 17060 11480 17066
rect 11428 17002 11480 17008
rect 11164 16794 11192 17002
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 11072 15706 11100 16594
rect 11164 16114 11192 16730
rect 11440 16726 11468 17002
rect 11428 16720 11480 16726
rect 11428 16662 11480 16668
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11072 14822 11100 15642
rect 11152 15360 11204 15366
rect 11150 15328 11152 15337
rect 11204 15328 11206 15337
rect 11150 15263 11206 15272
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 11164 14278 11192 15030
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11164 13870 11192 14214
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11348 13258 11376 13670
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11440 13190 11468 16662
rect 11532 15745 11560 20703
rect 11624 16289 11652 21406
rect 11610 16280 11666 16289
rect 11610 16215 11666 16224
rect 11624 15881 11652 16215
rect 11610 15872 11666 15881
rect 11610 15807 11666 15816
rect 11518 15736 11574 15745
rect 11518 15671 11574 15680
rect 11716 13410 11744 27520
rect 12164 26308 12216 26314
rect 12164 26250 12216 26256
rect 11888 25288 11940 25294
rect 11888 25230 11940 25236
rect 11900 24886 11928 25230
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 11888 24880 11940 24886
rect 11888 24822 11940 24828
rect 11900 24614 11928 24822
rect 11888 24608 11940 24614
rect 11888 24550 11940 24556
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 11808 22817 11836 23122
rect 11794 22808 11850 22817
rect 11794 22743 11850 22752
rect 11808 22710 11836 22743
rect 11796 22704 11848 22710
rect 11796 22646 11848 22652
rect 11900 21962 11928 24550
rect 11888 21956 11940 21962
rect 11888 21898 11940 21904
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 11808 21418 11836 21830
rect 11900 21690 11928 21898
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11796 21412 11848 21418
rect 11796 21354 11848 21360
rect 11992 21146 12020 24890
rect 12072 24064 12124 24070
rect 12072 24006 12124 24012
rect 12084 23594 12112 24006
rect 12072 23588 12124 23594
rect 12072 23530 12124 23536
rect 12072 23248 12124 23254
rect 12072 23190 12124 23196
rect 12084 23089 12112 23190
rect 12070 23080 12126 23089
rect 12070 23015 12126 23024
rect 12084 22710 12112 23015
rect 12072 22704 12124 22710
rect 12072 22646 12124 22652
rect 11980 21140 12032 21146
rect 11980 21082 12032 21088
rect 11796 20256 11848 20262
rect 11796 20198 11848 20204
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11808 20058 11836 20198
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11808 19514 11836 19994
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11900 18834 11928 20198
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11900 18426 11928 18770
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11886 18320 11942 18329
rect 11886 18255 11942 18264
rect 11900 17882 11928 18255
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11992 16998 12020 21082
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11900 15978 11928 16526
rect 11978 16008 12034 16017
rect 11888 15972 11940 15978
rect 11978 15943 12034 15952
rect 11888 15914 11940 15920
rect 11900 15162 11928 15914
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11888 14340 11940 14346
rect 11888 14282 11940 14288
rect 11900 13530 11928 14282
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11624 13382 11744 13410
rect 11888 13388 11940 13394
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11072 12850 11100 13126
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 11072 12306 11100 12650
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11072 10266 11100 11154
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 9654 11100 9862
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11164 9586 11192 12038
rect 11256 11762 11284 12582
rect 11440 12374 11468 12786
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11532 11665 11560 13126
rect 11624 13025 11652 13382
rect 11888 13330 11940 13336
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11610 13016 11666 13025
rect 11610 12951 11666 12960
rect 11624 12617 11652 12951
rect 11610 12608 11666 12617
rect 11610 12543 11666 12552
rect 11716 12442 11744 13262
rect 11794 13152 11850 13161
rect 11794 13087 11850 13096
rect 11808 12889 11836 13087
rect 11900 12986 11928 13330
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11794 12880 11850 12889
rect 11794 12815 11850 12824
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11808 12374 11836 12815
rect 11886 12608 11942 12617
rect 11886 12543 11942 12552
rect 11796 12368 11848 12374
rect 11900 12345 11928 12543
rect 11796 12310 11848 12316
rect 11886 12336 11942 12345
rect 11808 11898 11836 12310
rect 11886 12271 11942 12280
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11518 11656 11574 11665
rect 11518 11591 11574 11600
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11256 10538 11284 11086
rect 11348 10810 11376 11154
rect 11518 10976 11574 10985
rect 11518 10911 11574 10920
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11244 10532 11296 10538
rect 11244 10474 11296 10480
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11164 9081 11192 9318
rect 11150 9072 11206 9081
rect 11150 9007 11206 9016
rect 11060 8968 11112 8974
rect 11256 8956 11284 9318
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11112 8928 11284 8956
rect 11060 8910 11112 8916
rect 11072 8634 11100 8910
rect 11348 8634 11376 8978
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11164 7274 11192 8026
rect 11440 8022 11468 10406
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11256 7410 11284 7686
rect 11440 7546 11468 7958
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 10966 6896 11022 6905
rect 10966 6831 10968 6840
rect 11020 6831 11022 6840
rect 11428 6860 11480 6866
rect 10968 6802 11020 6808
rect 11428 6802 11480 6808
rect 10980 6254 11008 6802
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10138 6080 10194 6089
rect 10138 6015 10194 6024
rect 10152 4826 10180 6015
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10888 5778 10916 6122
rect 11072 5896 11100 6734
rect 11242 6624 11298 6633
rect 11242 6559 11298 6568
rect 11256 6322 11284 6559
rect 11440 6458 11468 6802
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11072 5868 11192 5896
rect 10876 5772 10928 5778
rect 10928 5732 11008 5760
rect 10876 5714 10928 5720
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10152 4282 10180 4762
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10704 4214 10732 4966
rect 10888 4865 10916 5510
rect 10980 5370 11008 5732
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 10874 4856 10930 4865
rect 10874 4791 10930 4800
rect 10980 4570 11008 5306
rect 11164 5166 11192 5868
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 11440 5030 11468 5782
rect 11532 5545 11560 10911
rect 11888 9920 11940 9926
rect 11794 9888 11850 9897
rect 11888 9862 11940 9868
rect 11794 9823 11850 9832
rect 11808 9654 11836 9823
rect 11796 9648 11848 9654
rect 11900 9625 11928 9862
rect 11796 9590 11848 9596
rect 11886 9616 11942 9625
rect 11886 9551 11942 9560
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11610 8256 11666 8265
rect 11610 8191 11666 8200
rect 11624 8022 11652 8191
rect 11716 8022 11744 8570
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11624 7721 11652 7958
rect 11610 7712 11666 7721
rect 11610 7647 11666 7656
rect 11624 7478 11652 7647
rect 11716 7546 11744 7958
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11992 7018 12020 15943
rect 12084 8430 12112 18022
rect 12176 9466 12204 26250
rect 12268 18272 12296 27520
rect 12440 24608 12492 24614
rect 12360 24556 12440 24562
rect 12360 24550 12492 24556
rect 12360 24534 12480 24550
rect 12360 21729 12388 24534
rect 12440 23724 12492 23730
rect 12440 23666 12492 23672
rect 12452 22710 12480 23666
rect 12716 23248 12768 23254
rect 12716 23190 12768 23196
rect 12728 22778 12756 23190
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 12624 22568 12676 22574
rect 12624 22510 12676 22516
rect 12636 22098 12664 22510
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 12530 21992 12586 22001
rect 12530 21927 12586 21936
rect 12346 21720 12402 21729
rect 12544 21690 12572 21927
rect 12636 21865 12664 22034
rect 12622 21856 12678 21865
rect 12622 21791 12678 21800
rect 12346 21655 12402 21664
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12360 19174 12388 19246
rect 12348 19168 12400 19174
rect 12348 19110 12400 19116
rect 12268 18244 12388 18272
rect 12256 18148 12308 18154
rect 12256 18090 12308 18096
rect 12268 17882 12296 18090
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12360 15042 12388 18244
rect 12452 17814 12480 21558
rect 12532 21412 12584 21418
rect 12532 21354 12584 21360
rect 12544 21146 12572 21354
rect 12532 21140 12584 21146
rect 12532 21082 12584 21088
rect 12532 20528 12584 20534
rect 12530 20496 12532 20505
rect 12584 20496 12586 20505
rect 12530 20431 12586 20440
rect 12820 19990 12848 27520
rect 13372 24834 13400 27520
rect 13372 24806 13584 24834
rect 13452 22092 13504 22098
rect 13452 22034 13504 22040
rect 13084 21956 13136 21962
rect 13084 21898 13136 21904
rect 13096 21486 13124 21898
rect 13360 21684 13412 21690
rect 13360 21626 13412 21632
rect 13084 21480 13136 21486
rect 13084 21422 13136 21428
rect 13096 21146 13124 21422
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 12990 20904 13046 20913
rect 12990 20839 13046 20848
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12912 20466 12940 20742
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12900 20324 12952 20330
rect 12900 20266 12952 20272
rect 12912 20058 12940 20266
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12808 19984 12860 19990
rect 12808 19926 12860 19932
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12530 19272 12586 19281
rect 12912 19242 12940 19654
rect 12530 19207 12586 19216
rect 12900 19236 12952 19242
rect 12544 18426 12572 19207
rect 12900 19178 12952 19184
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12636 18748 12664 19110
rect 12716 18760 12768 18766
rect 12636 18720 12716 18748
rect 12716 18702 12768 18708
rect 12728 18426 12756 18702
rect 12912 18630 12940 19178
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12912 18154 12940 18566
rect 12900 18148 12952 18154
rect 12900 18090 12952 18096
rect 13004 18086 13032 20839
rect 13372 19514 13400 21626
rect 13464 21622 13492 22034
rect 13452 21616 13504 21622
rect 13452 21558 13504 21564
rect 13450 21040 13506 21049
rect 13450 20975 13506 20984
rect 13464 20602 13492 20975
rect 13452 20596 13504 20602
rect 13452 20538 13504 20544
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13464 19378 13492 20198
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13096 18329 13124 18566
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13082 18320 13138 18329
rect 13082 18255 13084 18264
rect 13136 18255 13138 18264
rect 13084 18226 13136 18232
rect 13096 18195 13124 18226
rect 13464 18086 13492 18362
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13004 17814 13032 18022
rect 13174 17912 13230 17921
rect 13174 17847 13230 17856
rect 13360 17876 13412 17882
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12992 17808 13044 17814
rect 12992 17750 13044 17756
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12452 15094 12480 16730
rect 12716 16720 12768 16726
rect 12820 16697 12848 17478
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12716 16662 12768 16668
rect 12806 16688 12862 16697
rect 12728 15910 12756 16662
rect 12806 16623 12862 16632
rect 12912 15978 12940 16934
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12728 15570 12756 15846
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12268 15014 12388 15042
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12268 12481 12296 15014
rect 12452 14822 12480 15030
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 12900 14884 12952 14890
rect 12900 14826 12952 14832
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12544 14278 12572 14826
rect 12912 14618 12940 14826
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 12532 14272 12584 14278
rect 12912 14249 12940 14554
rect 13004 14498 13032 17750
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 13096 17338 13124 17682
rect 13188 17678 13216 17847
rect 13360 17818 13412 17824
rect 13268 17808 13320 17814
rect 13268 17750 13320 17756
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13096 16726 13124 17274
rect 13084 16720 13136 16726
rect 13084 16662 13136 16668
rect 13188 16182 13216 17614
rect 13280 16250 13308 17750
rect 13372 17134 13400 17818
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13372 16794 13400 17070
rect 13464 17066 13492 18022
rect 13452 17060 13504 17066
rect 13452 17002 13504 17008
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13176 16176 13228 16182
rect 13176 16118 13228 16124
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 13096 14890 13124 15302
rect 13280 15162 13308 16186
rect 13358 16144 13414 16153
rect 13358 16079 13414 16088
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13084 14884 13136 14890
rect 13084 14826 13136 14832
rect 13004 14470 13124 14498
rect 12532 14214 12584 14220
rect 12898 14240 12954 14249
rect 12544 13802 12572 14214
rect 12898 14175 12954 14184
rect 12622 13832 12678 13841
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12532 13796 12584 13802
rect 12808 13796 12860 13802
rect 12622 13767 12678 13776
rect 12532 13738 12584 13744
rect 12360 13462 12388 13738
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 12544 13326 12572 13738
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12254 12472 12310 12481
rect 12254 12407 12310 12416
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12452 10282 12480 12378
rect 12636 12102 12664 13767
rect 12728 13756 12808 13784
rect 12728 13394 12756 13756
rect 12808 13738 12860 13744
rect 12806 13424 12862 13433
rect 12716 13388 12768 13394
rect 12806 13359 12862 13368
rect 12716 13330 12768 13336
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12728 12458 12756 12854
rect 12820 12594 12848 13359
rect 12898 13152 12954 13161
rect 12898 13087 12954 13096
rect 12912 12986 12940 13087
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12912 12782 12940 12922
rect 13096 12918 13124 14470
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 12900 12776 12952 12782
rect 13188 12764 13216 14350
rect 12900 12718 12952 12724
rect 13096 12736 13216 12764
rect 12820 12566 12940 12594
rect 12728 12442 12848 12458
rect 12728 12436 12860 12442
rect 12728 12430 12808 12436
rect 12808 12378 12860 12384
rect 12820 12347 12848 12378
rect 12714 12336 12770 12345
rect 12714 12271 12770 12280
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12532 11824 12584 11830
rect 12728 11801 12756 12271
rect 12912 12170 12940 12566
rect 12990 12336 13046 12345
rect 12990 12271 13046 12280
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 13004 12102 13032 12271
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 12532 11766 12584 11772
rect 12714 11792 12770 11801
rect 12544 10849 12572 11766
rect 12714 11727 12770 11736
rect 13004 11626 13032 12038
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 12714 11112 12770 11121
rect 12714 11047 12770 11056
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12530 10840 12586 10849
rect 12530 10775 12586 10784
rect 12636 10606 12664 10950
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12452 10254 12572 10282
rect 12440 10192 12492 10198
rect 12360 10140 12440 10146
rect 12360 10134 12492 10140
rect 12360 10118 12480 10134
rect 12360 9897 12388 10118
rect 12346 9888 12402 9897
rect 12346 9823 12402 9832
rect 12346 9616 12402 9625
rect 12544 9602 12572 10254
rect 12636 10062 12664 10542
rect 12728 10130 12756 11047
rect 12898 10704 12954 10713
rect 12898 10639 12954 10648
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12544 9574 12664 9602
rect 12346 9551 12402 9560
rect 12360 9500 12388 9551
rect 12360 9472 12572 9500
rect 12176 9438 12296 9466
rect 12268 9330 12296 9438
rect 12268 9302 12480 9330
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12268 7410 12296 9302
rect 12452 9178 12480 9302
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12360 8945 12388 8978
rect 12346 8936 12402 8945
rect 12346 8871 12402 8880
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12452 8106 12480 8502
rect 12360 8090 12480 8106
rect 12348 8084 12480 8090
rect 12400 8078 12480 8084
rect 12348 8026 12400 8032
rect 12544 7410 12572 9472
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 11992 6990 12112 7018
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11900 6118 11928 6734
rect 11992 6390 12020 6802
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 11888 6112 11940 6118
rect 11886 6080 11888 6089
rect 11940 6080 11942 6089
rect 11886 6015 11942 6024
rect 11992 5642 12020 6326
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 11518 5536 11574 5545
rect 11518 5471 11574 5480
rect 11518 5400 11574 5409
rect 11574 5358 11836 5386
rect 11518 5335 11574 5344
rect 11808 5273 11836 5358
rect 11518 5264 11574 5273
rect 11518 5199 11574 5208
rect 11794 5264 11850 5273
rect 11794 5199 11850 5208
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 10888 4542 11008 4570
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10046 2544 10102 2553
rect 10046 2479 10102 2488
rect 10046 1184 10102 1193
rect 10152 1170 10180 3878
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2650 10732 4150
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10796 2417 10824 3674
rect 10888 3602 10916 4542
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10980 3924 11008 4422
rect 11348 4321 11376 4966
rect 11532 4321 11560 5199
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11334 4312 11390 4321
rect 11334 4247 11390 4256
rect 11518 4312 11574 4321
rect 11518 4247 11574 4256
rect 11060 3936 11112 3942
rect 10980 3896 11060 3924
rect 11060 3878 11112 3884
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 11060 3596 11112 3602
rect 11112 3556 11192 3584
rect 11060 3538 11112 3544
rect 10888 3194 10916 3538
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10888 2990 10916 3130
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 11164 2854 11192 3556
rect 11426 2952 11482 2961
rect 11426 2887 11482 2896
rect 11152 2848 11204 2854
rect 10874 2816 10930 2825
rect 11152 2790 11204 2796
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 10874 2751 10930 2760
rect 10782 2408 10838 2417
rect 10782 2343 10838 2352
rect 10152 1142 10456 1170
rect 10046 1119 10102 1128
rect 9876 1006 9996 1034
rect 9678 912 9734 921
rect 9678 847 9734 856
rect 9876 480 9904 1006
rect 10060 785 10088 1119
rect 10046 776 10102 785
rect 10046 711 10102 720
rect 10428 480 10456 1142
rect 10888 480 10916 2751
rect 11164 2650 11192 2790
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11256 2582 11284 2790
rect 11244 2576 11296 2582
rect 11150 2544 11206 2553
rect 11244 2518 11296 2524
rect 11150 2479 11152 2488
rect 11204 2479 11206 2488
rect 11152 2450 11204 2456
rect 11440 480 11468 2887
rect 11716 2854 11744 4966
rect 12084 4622 12112 6990
rect 12360 6866 12388 7278
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12452 6254 12480 6598
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12360 5574 12388 6122
rect 12348 5568 12400 5574
rect 12162 5536 12218 5545
rect 12348 5510 12400 5516
rect 12162 5471 12218 5480
rect 12176 4826 12204 5471
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12084 4282 12112 4558
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11900 2378 11928 4014
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11532 1465 11560 2246
rect 11518 1456 11574 1465
rect 11518 1391 11574 1400
rect 11992 480 12020 4150
rect 12084 2922 12112 4218
rect 12176 4146 12204 4762
rect 12360 4690 12388 5510
rect 12452 5370 12480 6190
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12440 5160 12492 5166
rect 12636 5114 12664 9574
rect 12728 9178 12756 10066
rect 12912 9654 12940 10639
rect 12900 9648 12952 9654
rect 13096 9625 13124 12736
rect 13372 12374 13400 16079
rect 13450 15328 13506 15337
rect 13450 15263 13506 15272
rect 13360 12368 13412 12374
rect 13360 12310 13412 12316
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13188 12209 13216 12242
rect 13464 12238 13492 15263
rect 13268 12232 13320 12238
rect 13174 12200 13230 12209
rect 13268 12174 13320 12180
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13174 12135 13230 12144
rect 13188 11354 13216 12135
rect 13280 11626 13308 12174
rect 13360 12164 13412 12170
rect 13360 12106 13412 12112
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13280 11121 13308 11562
rect 13266 11112 13322 11121
rect 13266 11047 13268 11056
rect 13320 11047 13322 11056
rect 13268 11018 13320 11024
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13188 10198 13216 10746
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13188 9722 13216 10134
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13372 9654 13400 12106
rect 13464 11898 13492 12174
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13556 10538 13584 24806
rect 13634 23624 13690 23633
rect 13634 23559 13690 23568
rect 13648 22953 13676 23559
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13832 23322 13860 23462
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 13728 22976 13780 22982
rect 13634 22944 13690 22953
rect 13728 22918 13780 22924
rect 13634 22879 13690 22888
rect 13740 22273 13768 22918
rect 13818 22536 13874 22545
rect 13818 22471 13874 22480
rect 13726 22264 13782 22273
rect 13832 22234 13860 22471
rect 13726 22199 13782 22208
rect 13820 22228 13872 22234
rect 13820 22170 13872 22176
rect 13832 21690 13860 22170
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 13636 20800 13688 20806
rect 13636 20742 13688 20748
rect 13648 19281 13676 20742
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13740 20346 13768 20402
rect 13924 20346 13952 27520
rect 14004 25356 14056 25362
rect 14004 25298 14056 25304
rect 14016 24614 14044 25298
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 14016 20482 14044 24550
rect 14280 24200 14332 24206
rect 14280 24142 14332 24148
rect 14292 23526 14320 24142
rect 14188 23520 14240 23526
rect 14188 23462 14240 23468
rect 14280 23520 14332 23526
rect 14280 23462 14332 23468
rect 14200 22506 14228 23462
rect 14292 23225 14320 23462
rect 14278 23216 14334 23225
rect 14278 23151 14334 23160
rect 14188 22500 14240 22506
rect 14188 22442 14240 22448
rect 14200 22234 14228 22442
rect 14188 22228 14240 22234
rect 14188 22170 14240 22176
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14292 21078 14320 22170
rect 14188 21072 14240 21078
rect 14186 21040 14188 21049
rect 14280 21072 14332 21078
rect 14240 21040 14242 21049
rect 14096 21004 14148 21010
rect 14280 21014 14332 21020
rect 14186 20975 14242 20984
rect 14096 20946 14148 20952
rect 14108 20602 14136 20946
rect 14292 20602 14320 21014
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14016 20454 14136 20482
rect 13740 20318 13860 20346
rect 13924 20318 14044 20346
rect 13832 20210 13860 20318
rect 13832 20182 13952 20210
rect 13818 19952 13874 19961
rect 13818 19887 13820 19896
rect 13872 19887 13874 19896
rect 13820 19858 13872 19864
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13740 19417 13768 19654
rect 13832 19514 13860 19858
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13726 19408 13782 19417
rect 13726 19343 13782 19352
rect 13634 19272 13690 19281
rect 13634 19207 13690 19216
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 18834 13860 19110
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13924 18426 13952 20182
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 14016 16810 14044 20318
rect 14108 18222 14136 20454
rect 14292 20330 14320 20538
rect 14280 20324 14332 20330
rect 14280 20266 14332 20272
rect 14292 19990 14320 20266
rect 14188 19984 14240 19990
rect 14188 19926 14240 19932
rect 14280 19984 14332 19990
rect 14280 19926 14332 19932
rect 14200 19258 14228 19926
rect 14200 19230 14320 19258
rect 14292 19174 14320 19230
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14188 18148 14240 18154
rect 14188 18090 14240 18096
rect 14200 17882 14228 18090
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 13924 16782 14044 16810
rect 13818 15736 13874 15745
rect 13818 15671 13820 15680
rect 13872 15671 13874 15680
rect 13820 15642 13872 15648
rect 13924 15502 13952 16782
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 14016 16046 14044 16662
rect 14186 16552 14242 16561
rect 14186 16487 14242 16496
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 14094 16008 14150 16017
rect 14094 15943 14150 15952
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13924 15178 13952 15438
rect 13740 15162 13952 15178
rect 14016 15162 14044 15642
rect 13728 15156 13952 15162
rect 13780 15150 13952 15156
rect 14004 15156 14056 15162
rect 13728 15098 13780 15104
rect 14004 15098 14056 15104
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13740 13462 13768 13670
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13832 13274 13860 14214
rect 13740 13246 13860 13274
rect 13740 11778 13768 13246
rect 14016 12866 14044 15098
rect 14108 14278 14136 15943
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14200 13954 14228 16487
rect 14292 15745 14320 19110
rect 14278 15736 14334 15745
rect 14278 15671 14334 15680
rect 14384 15552 14412 27520
rect 14936 25242 14964 27520
rect 14844 25214 14964 25242
rect 14554 23896 14610 23905
rect 14554 23831 14610 23840
rect 14462 23352 14518 23361
rect 14462 23287 14518 23296
rect 14476 23118 14504 23287
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14476 22778 14504 23054
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14464 22092 14516 22098
rect 14464 22034 14516 22040
rect 14476 21690 14504 22034
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14464 19440 14516 19446
rect 14464 19382 14516 19388
rect 14292 15524 14412 15552
rect 14292 14414 14320 15524
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14292 14074 14320 14350
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14200 13926 14320 13954
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 14108 12986 14136 13398
rect 14186 13288 14242 13297
rect 14186 13223 14242 13232
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14016 12838 14136 12866
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13832 11898 13860 12310
rect 14016 12306 14044 12650
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13740 11750 13860 11778
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13360 9648 13412 9654
rect 12900 9590 12952 9596
rect 13082 9616 13138 9625
rect 13360 9590 13412 9596
rect 13450 9616 13506 9625
rect 13082 9551 13138 9560
rect 13450 9551 13506 9560
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 13082 8936 13138 8945
rect 13082 8871 13138 8880
rect 13096 8498 13124 8871
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12990 8392 13046 8401
rect 12714 7168 12770 7177
rect 12714 7103 12770 7112
rect 12728 6866 12756 7103
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12728 6458 12756 6802
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12728 5914 12756 6394
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12440 5102 12492 5108
rect 12452 4865 12480 5102
rect 12544 5086 12664 5114
rect 12716 5092 12768 5098
rect 12438 4856 12494 4865
rect 12438 4791 12494 4800
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12544 4570 12572 5086
rect 12716 5034 12768 5040
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12452 4542 12572 4570
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12360 4078 12388 4490
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12256 4004 12308 4010
rect 12256 3946 12308 3952
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 12268 2378 12296 3946
rect 12452 3369 12480 4542
rect 12636 4321 12664 4966
rect 12622 4312 12678 4321
rect 12622 4247 12678 4256
rect 12728 4162 12756 5034
rect 12636 4134 12756 4162
rect 12636 3924 12664 4134
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12544 3896 12664 3924
rect 12438 3360 12494 3369
rect 12438 3295 12494 3304
rect 12438 3088 12494 3097
rect 12438 3023 12494 3032
rect 12452 2582 12480 3023
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12256 2372 12308 2378
rect 12256 2314 12308 2320
rect 12544 480 12572 3896
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12636 2922 12664 3674
rect 12728 3641 12756 3946
rect 12714 3632 12770 3641
rect 12714 3567 12770 3576
rect 12714 3360 12770 3369
rect 12714 3295 12770 3304
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 12728 2582 12756 3295
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 12912 1902 12940 8366
rect 12990 8327 13046 8336
rect 13004 7954 13032 8327
rect 13464 8294 13492 9551
rect 13648 9518 13676 10406
rect 13740 10266 13768 11154
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13648 9382 13676 9454
rect 13636 9376 13688 9382
rect 13688 9336 13768 9364
rect 13636 9318 13688 9324
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13556 8362 13584 9046
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 13464 7818 13492 8230
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13280 7342 13308 7686
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13082 4992 13138 5001
rect 13082 4927 13138 4936
rect 12900 1896 12952 1902
rect 12900 1838 12952 1844
rect 13096 480 13124 4927
rect 13188 3942 13216 7142
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13280 3670 13308 4626
rect 13372 4146 13400 5170
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13268 3664 13320 3670
rect 13266 3632 13268 3641
rect 13320 3632 13322 3641
rect 13266 3567 13322 3576
rect 13358 3496 13414 3505
rect 13358 3431 13360 3440
rect 13412 3431 13414 3440
rect 13360 3402 13412 3408
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13188 1601 13216 2518
rect 13464 2514 13492 7754
rect 13556 5409 13584 8298
rect 13648 7886 13676 8774
rect 13740 8566 13768 9336
rect 13832 9110 13860 11750
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13924 9518 13952 9862
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13924 8634 13952 9454
rect 14016 9217 14044 11086
rect 14002 9208 14058 9217
rect 14002 9143 14058 9152
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13924 8022 13952 8570
rect 14108 8514 14136 12838
rect 14200 12442 14228 13223
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14200 11694 14228 12378
rect 14292 11778 14320 13926
rect 14384 11914 14412 15370
rect 14476 14498 14504 19382
rect 14568 18442 14596 23831
rect 14740 23520 14792 23526
rect 14740 23462 14792 23468
rect 14648 23180 14700 23186
rect 14648 23122 14700 23128
rect 14660 22778 14688 23122
rect 14648 22772 14700 22778
rect 14648 22714 14700 22720
rect 14646 22400 14702 22409
rect 14646 22335 14702 22344
rect 14660 20641 14688 22335
rect 14752 21690 14780 23462
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 14740 21480 14792 21486
rect 14740 21422 14792 21428
rect 14646 20632 14702 20641
rect 14646 20567 14702 20576
rect 14752 19514 14780 21422
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14740 18896 14792 18902
rect 14740 18838 14792 18844
rect 14752 18601 14780 18838
rect 14738 18592 14794 18601
rect 14738 18527 14794 18536
rect 14568 18414 14688 18442
rect 14752 18426 14780 18527
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14568 17882 14596 18226
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14568 15620 14596 15846
rect 14660 15722 14688 18414
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 14660 15694 14780 15722
rect 14568 15592 14688 15620
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 14822 14596 15438
rect 14660 14958 14688 15592
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14556 14816 14608 14822
rect 14554 14784 14556 14793
rect 14608 14784 14610 14793
rect 14554 14719 14610 14728
rect 14752 14498 14780 15694
rect 14476 14470 14596 14498
rect 14660 14482 14780 14498
rect 14384 11886 14504 11914
rect 14292 11750 14412 11778
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 14292 10130 14320 11562
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14200 9761 14228 9930
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14186 9752 14242 9761
rect 14186 9687 14242 9696
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14016 8486 14136 8514
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13912 8016 13964 8022
rect 13912 7958 13964 7964
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13648 6934 13676 7822
rect 13740 7546 13768 7958
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13924 7478 13952 7958
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 13636 6928 13688 6934
rect 13636 6870 13688 6876
rect 14016 6798 14044 8486
rect 14200 8090 14228 8910
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14186 7576 14242 7585
rect 14186 7511 14242 7520
rect 14200 6934 14228 7511
rect 14188 6928 14240 6934
rect 14188 6870 14240 6876
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 14016 6089 14044 6598
rect 14002 6080 14058 6089
rect 14058 6038 14136 6066
rect 14002 6015 14058 6024
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13832 5658 13860 5714
rect 13740 5630 13860 5658
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13542 5400 13598 5409
rect 13542 5335 13598 5344
rect 13634 5264 13690 5273
rect 13634 5199 13690 5208
rect 13648 4826 13676 5199
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13556 4010 13584 4694
rect 13648 4282 13676 4762
rect 13740 4486 13768 5630
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 13174 1592 13230 1601
rect 13174 1527 13230 1536
rect 13648 480 13676 3878
rect 13740 3670 13768 4422
rect 13832 3738 13860 5510
rect 13924 5030 13952 5646
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 14016 4554 14044 5782
rect 14108 5166 14136 6038
rect 14292 5642 14320 9862
rect 14384 9518 14412 11750
rect 14476 9659 14504 11886
rect 14462 9650 14518 9659
rect 14462 9585 14518 9594
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14476 7410 14504 9454
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14108 4826 14136 5102
rect 14280 5092 14332 5098
rect 14280 5034 14332 5040
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14292 4729 14320 5034
rect 14278 4720 14334 4729
rect 14278 4655 14334 4664
rect 14004 4548 14056 4554
rect 14004 4490 14056 4496
rect 14384 4128 14412 6734
rect 14568 6236 14596 14470
rect 14648 14476 14780 14482
rect 14700 14470 14780 14476
rect 14648 14418 14700 14424
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14660 13802 14688 14214
rect 14752 14074 14780 14470
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14660 12986 14688 13738
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14660 10810 14688 11154
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14660 9178 14688 10066
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14660 8362 14688 8910
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14660 8022 14688 8298
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 14660 7410 14688 7958
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14660 7002 14688 7346
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14476 6208 14596 6236
rect 14476 5370 14504 6208
rect 14554 5944 14610 5953
rect 14554 5879 14610 5888
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14476 4282 14504 5306
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14292 4100 14412 4128
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13832 2689 13860 3674
rect 14292 3233 14320 4100
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14384 3466 14412 3946
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14476 3534 14504 3878
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 14278 3224 14334 3233
rect 14476 3194 14504 3470
rect 14278 3159 14334 3168
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 13818 2680 13874 2689
rect 13818 2615 13874 2624
rect 14186 2544 14242 2553
rect 14186 2479 14242 2488
rect 14200 2009 14228 2479
rect 14476 2446 14504 3130
rect 14464 2440 14516 2446
rect 14370 2408 14426 2417
rect 14464 2382 14516 2388
rect 14370 2343 14372 2352
rect 14424 2343 14426 2352
rect 14372 2314 14424 2320
rect 14568 2281 14596 5879
rect 14646 5536 14702 5545
rect 14646 5471 14702 5480
rect 14660 4729 14688 5471
rect 14646 4720 14702 4729
rect 14646 4655 14702 4664
rect 14554 2272 14610 2281
rect 14554 2207 14610 2216
rect 14186 2000 14242 2009
rect 14186 1935 14242 1944
rect 14646 2000 14702 2009
rect 14646 1935 14702 1944
rect 14188 1896 14240 1902
rect 14188 1838 14240 1844
rect 14200 480 14228 1838
rect 14660 480 14688 1935
rect 14752 1601 14780 14010
rect 14844 12594 14872 25214
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15488 24698 15516 27520
rect 15120 24670 15516 24698
rect 15120 24614 15148 24670
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 15580 24313 15608 24550
rect 15566 24304 15622 24313
rect 15292 24268 15344 24274
rect 15566 24239 15622 24248
rect 15292 24210 15344 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15304 23866 15332 24210
rect 15292 23860 15344 23866
rect 15292 23802 15344 23808
rect 15936 23248 15988 23254
rect 15934 23216 15936 23225
rect 15988 23216 15990 23225
rect 15934 23151 15990 23160
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15016 22704 15068 22710
rect 15016 22646 15068 22652
rect 15028 22234 15056 22646
rect 15016 22228 15068 22234
rect 15016 22170 15068 22176
rect 15396 22098 15424 22918
rect 15856 22506 15884 23054
rect 15948 22658 15976 23151
rect 16040 22778 16068 27520
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 15948 22630 16068 22658
rect 15844 22500 15896 22506
rect 15844 22442 15896 22448
rect 16040 22438 16068 22630
rect 16028 22432 16080 22438
rect 16026 22400 16028 22409
rect 16080 22400 16082 22409
rect 16026 22335 16082 22344
rect 15842 22264 15898 22273
rect 15842 22199 15844 22208
rect 15896 22199 15898 22208
rect 15844 22170 15896 22176
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15396 21350 15424 21830
rect 15660 21412 15712 21418
rect 15660 21354 15712 21360
rect 15752 21412 15804 21418
rect 15752 21354 15804 21360
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15028 21146 15056 21286
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 15672 21078 15700 21354
rect 15660 21072 15712 21078
rect 15382 21040 15438 21049
rect 15660 21014 15712 21020
rect 15764 21010 15792 21354
rect 15856 21146 15884 22170
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 16040 21350 16068 21966
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 16040 21026 16068 21286
rect 15948 21010 16068 21026
rect 15382 20975 15438 20984
rect 15752 21004 15804 21010
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15292 19304 15344 19310
rect 15290 19272 15292 19281
rect 15344 19272 15346 19281
rect 15290 19207 15346 19216
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15290 19136 15346 19145
rect 15028 18970 15056 19110
rect 15290 19071 15346 19080
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15304 17610 15332 19071
rect 15396 18714 15424 20975
rect 15752 20946 15804 20952
rect 15936 21004 16068 21010
rect 15988 20998 16068 21004
rect 15936 20946 15988 20952
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15672 20398 15700 20878
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 15672 20058 15700 20334
rect 16040 20262 16068 20998
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 15934 19816 15990 19825
rect 15844 19780 15896 19786
rect 15934 19751 15990 19760
rect 15844 19722 15896 19728
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 15474 19408 15530 19417
rect 15474 19343 15530 19352
rect 15488 19242 15516 19343
rect 15580 19242 15608 19654
rect 15476 19236 15528 19242
rect 15476 19178 15528 19184
rect 15568 19236 15620 19242
rect 15568 19178 15620 19184
rect 15488 18970 15516 19178
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15658 18864 15714 18873
rect 15658 18799 15660 18808
rect 15712 18799 15714 18808
rect 15660 18770 15712 18776
rect 15396 18686 15516 18714
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15396 18290 15424 18566
rect 15384 18284 15436 18290
rect 15384 18226 15436 18232
rect 15382 18184 15438 18193
rect 15382 18119 15384 18128
rect 15436 18119 15438 18128
rect 15384 18090 15436 18096
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 15396 17490 15424 17682
rect 15304 17462 15424 17490
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15304 16998 15332 17462
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15304 16561 15332 16934
rect 15488 16794 15516 18686
rect 15672 18442 15700 18770
rect 15672 18426 15792 18442
rect 15672 18420 15804 18426
rect 15672 18414 15752 18420
rect 15752 18362 15804 18368
rect 15856 18306 15884 19722
rect 15948 18902 15976 19751
rect 16040 19718 16068 20198
rect 16132 19786 16160 24550
rect 16592 24426 16620 27520
rect 16500 24410 16620 24426
rect 16488 24404 16620 24410
rect 16540 24398 16620 24404
rect 16488 24346 16540 24352
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16408 23866 16436 24210
rect 17144 23866 17172 27520
rect 17696 25514 17724 27520
rect 17512 25486 17724 25514
rect 17406 24440 17462 24449
rect 17512 24410 17540 25486
rect 18248 24698 18276 27520
rect 17880 24670 18276 24698
rect 18326 24712 18382 24721
rect 17682 24440 17738 24449
rect 17406 24375 17462 24384
rect 17500 24404 17552 24410
rect 17420 24274 17448 24375
rect 17682 24375 17684 24384
rect 17500 24346 17552 24352
rect 17736 24375 17738 24384
rect 17684 24346 17736 24352
rect 17408 24268 17460 24274
rect 17408 24210 17460 24216
rect 17420 23866 17448 24210
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 17132 23860 17184 23866
rect 17132 23802 17184 23808
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 16856 23656 16908 23662
rect 16854 23624 16856 23633
rect 16908 23624 16910 23633
rect 16854 23559 16910 23568
rect 17880 23322 17908 24670
rect 18326 24647 18382 24656
rect 17868 23316 17920 23322
rect 17868 23258 17920 23264
rect 17958 23216 18014 23225
rect 16764 23180 16816 23186
rect 17958 23151 17960 23160
rect 16764 23122 16816 23128
rect 18012 23151 18014 23160
rect 17960 23122 18012 23128
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 16212 22432 16264 22438
rect 16212 22374 16264 22380
rect 16224 22098 16252 22374
rect 16316 22234 16344 22510
rect 16776 22438 16804 23122
rect 17972 22778 18000 23122
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16212 22092 16264 22098
rect 16212 22034 16264 22040
rect 16120 19780 16172 19786
rect 16120 19722 16172 19728
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 16224 19394 16252 22034
rect 16776 21457 16804 22374
rect 16948 22092 17000 22098
rect 16948 22034 17000 22040
rect 16960 21690 16988 22034
rect 17038 21992 17094 22001
rect 17038 21927 17040 21936
rect 17092 21927 17094 21936
rect 17040 21898 17092 21904
rect 18340 21690 18368 24647
rect 18800 24449 18828 27520
rect 18786 24440 18842 24449
rect 18786 24375 18842 24384
rect 18694 23896 18750 23905
rect 18694 23831 18696 23840
rect 18748 23831 18750 23840
rect 18696 23802 18748 23808
rect 18512 23656 18564 23662
rect 18512 23598 18564 23604
rect 16948 21684 17000 21690
rect 16948 21626 17000 21632
rect 18328 21684 18380 21690
rect 18328 21626 18380 21632
rect 18328 21480 18380 21486
rect 16762 21448 16818 21457
rect 18328 21422 18380 21428
rect 16762 21383 16818 21392
rect 16488 21072 16540 21078
rect 16488 21014 16540 21020
rect 16500 19990 16528 21014
rect 18050 20496 18106 20505
rect 18340 20466 18368 21422
rect 18050 20431 18106 20440
rect 18328 20460 18380 20466
rect 18064 20398 18092 20431
rect 18328 20402 18380 20408
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 16488 19984 16540 19990
rect 16488 19926 16540 19932
rect 17222 19952 17278 19961
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16316 19514 16344 19858
rect 16500 19514 16528 19926
rect 17222 19887 17278 19896
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16040 19366 16252 19394
rect 16302 19408 16358 19417
rect 15936 18896 15988 18902
rect 15936 18838 15988 18844
rect 15764 18278 15884 18306
rect 15948 18290 15976 18838
rect 15936 18284 15988 18290
rect 15764 17746 15792 18278
rect 15936 18226 15988 18232
rect 15842 17912 15898 17921
rect 15842 17847 15898 17856
rect 15856 17814 15884 17847
rect 15948 17814 15976 18226
rect 15844 17808 15896 17814
rect 15844 17750 15896 17756
rect 15936 17808 15988 17814
rect 15936 17750 15988 17756
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15856 17338 15884 17750
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 15856 17105 15884 17274
rect 15842 17096 15898 17105
rect 15842 17031 15898 17040
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15290 16552 15346 16561
rect 15290 16487 15346 16496
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 15570 15332 16390
rect 15488 16114 15516 16730
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 15144 15332 15506
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15120 15116 15332 15144
rect 15120 14618 15148 15116
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 14936 13433 14964 13942
rect 15396 13938 15424 15302
rect 15488 14550 15516 15846
rect 15580 15434 15608 16594
rect 15856 16590 15884 16934
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 16250 15884 16526
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15580 14890 15608 15370
rect 15568 14884 15620 14890
rect 15568 14826 15620 14832
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 15028 13462 15056 13738
rect 15120 13530 15148 13874
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15016 13456 15068 13462
rect 14922 13424 14978 13433
rect 15016 13398 15068 13404
rect 14922 13359 14978 13368
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15488 12646 15516 13126
rect 15476 12640 15528 12646
rect 14844 12566 15056 12594
rect 15476 12582 15528 12588
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 14844 12102 14872 12310
rect 15028 12170 15056 12566
rect 15382 12472 15438 12481
rect 15382 12407 15438 12416
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14844 10810 14872 12038
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15212 11150 15240 11630
rect 15304 11626 15332 12038
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15304 11354 15332 11562
rect 15396 11370 15424 12407
rect 15488 12170 15516 12582
rect 15580 12306 15608 14826
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15672 14414 15700 14758
rect 15948 14618 15976 15574
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 16040 14498 16068 19366
rect 16302 19343 16358 19352
rect 16118 18320 16174 18329
rect 16118 18255 16174 18264
rect 16132 18154 16160 18255
rect 16120 18148 16172 18154
rect 16120 18090 16172 18096
rect 16316 16153 16344 19343
rect 16396 17808 16448 17814
rect 16396 17750 16448 17756
rect 16408 17338 16436 17750
rect 16396 17332 16448 17338
rect 16396 17274 16448 17280
rect 16670 16688 16726 16697
rect 16670 16623 16726 16632
rect 16302 16144 16358 16153
rect 16302 16079 16358 16088
rect 16684 16046 16712 16623
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16302 15872 16358 15881
rect 16302 15807 16358 15816
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16132 15162 16160 15438
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16132 14550 16160 15098
rect 15948 14470 16068 14498
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15672 13734 15700 14350
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15672 13326 15700 13670
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15750 13288 15806 13297
rect 15672 12646 15700 13262
rect 15750 13223 15806 13232
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15292 11348 15344 11354
rect 15396 11342 15516 11370
rect 15292 11290 15344 11296
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 15304 10674 15332 11290
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15488 10198 15516 11342
rect 15580 11268 15608 12242
rect 15764 12050 15792 13223
rect 15842 12336 15898 12345
rect 15842 12271 15898 12280
rect 15856 12238 15884 12271
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15672 12022 15792 12050
rect 15672 11506 15700 12022
rect 15856 11914 15884 12174
rect 15764 11898 15884 11914
rect 15752 11892 15884 11898
rect 15804 11886 15884 11892
rect 15752 11834 15804 11840
rect 15672 11478 15792 11506
rect 15660 11280 15712 11286
rect 15580 11240 15660 11268
rect 15660 11222 15712 11228
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15476 10192 15528 10198
rect 15382 10160 15438 10169
rect 15476 10134 15528 10140
rect 15382 10095 15438 10104
rect 15396 9994 15424 10095
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15488 9722 15516 10134
rect 15580 9926 15608 10406
rect 15568 9920 15620 9926
rect 15566 9888 15568 9897
rect 15620 9888 15622 9897
rect 15566 9823 15622 9832
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 14830 9616 14886 9625
rect 14830 9551 14886 9560
rect 14844 7206 14872 9551
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15212 8945 15240 9318
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15198 8936 15254 8945
rect 15198 8871 15254 8880
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14924 7880 14976 7886
rect 14922 7848 14924 7857
rect 14976 7848 14978 7857
rect 14922 7783 14978 7792
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14844 3738 14872 4966
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14844 3505 14872 3674
rect 14830 3496 14886 3505
rect 14830 3431 14886 3440
rect 14844 2922 14872 3431
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 14936 2650 14964 2926
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14738 1592 14794 1601
rect 14738 1527 14794 1536
rect 15304 1034 15332 8774
rect 15396 8634 15424 8978
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15396 8537 15424 8570
rect 15382 8528 15438 8537
rect 15382 8463 15438 8472
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 15396 7018 15424 7890
rect 15488 7449 15516 9658
rect 15568 7472 15620 7478
rect 15474 7440 15530 7449
rect 15568 7414 15620 7420
rect 15474 7375 15530 7384
rect 15396 6990 15516 7018
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15396 6458 15424 6802
rect 15488 6746 15516 6990
rect 15580 6905 15608 7414
rect 15566 6896 15622 6905
rect 15566 6831 15622 6840
rect 15488 6718 15608 6746
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15382 5536 15438 5545
rect 15382 5471 15438 5480
rect 15396 5370 15424 5471
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15212 1006 15332 1034
rect 15212 480 15240 1006
rect 15488 610 15516 6598
rect 15580 4826 15608 6718
rect 15672 5778 15700 10474
rect 15764 8401 15792 11478
rect 15948 11234 15976 14470
rect 16132 13462 16160 14486
rect 16120 13456 16172 13462
rect 16120 13398 16172 13404
rect 16132 12986 16160 13398
rect 16316 13161 16344 15807
rect 17236 15638 17264 19887
rect 17590 19816 17646 19825
rect 17590 19751 17592 19760
rect 17644 19751 17646 19760
rect 17592 19722 17644 19728
rect 18524 17921 18552 23598
rect 19062 23488 19118 23497
rect 19062 23423 19118 23432
rect 19076 22114 19104 23423
rect 19352 23338 19380 27520
rect 19904 25786 19932 27520
rect 19536 25758 19932 25786
rect 19536 24721 19564 25758
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19522 24712 19578 24721
rect 19522 24647 19578 24656
rect 19982 24712 20038 24721
rect 19982 24647 20038 24656
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19996 24410 20024 24647
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 20168 24268 20220 24274
rect 20168 24210 20220 24216
rect 20180 23526 20208 24210
rect 20456 23905 20484 27520
rect 20442 23896 20498 23905
rect 21008 23866 21036 27520
rect 21560 24721 21588 27520
rect 21546 24712 21602 24721
rect 21546 24647 21602 24656
rect 22006 23896 22062 23905
rect 20442 23831 20498 23840
rect 20996 23860 21048 23866
rect 22006 23831 22008 23840
rect 20996 23802 21048 23808
rect 22060 23831 22062 23840
rect 22008 23802 22060 23808
rect 22112 23746 22140 27520
rect 22664 23798 22692 27520
rect 23216 23905 23244 27520
rect 23480 25220 23532 25226
rect 23480 25162 23532 25168
rect 23202 23896 23258 23905
rect 23202 23831 23258 23840
rect 21928 23718 22140 23746
rect 22652 23792 22704 23798
rect 22652 23734 22704 23740
rect 20720 23656 20772 23662
rect 20718 23624 20720 23633
rect 21824 23656 21876 23662
rect 20772 23624 20774 23633
rect 21824 23598 21876 23604
rect 20718 23559 20774 23568
rect 19524 23520 19576 23526
rect 19524 23462 19576 23468
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 19260 23322 19380 23338
rect 19248 23316 19380 23322
rect 19300 23310 19380 23316
rect 19248 23258 19300 23264
rect 19076 22086 19288 22114
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19168 19174 19196 19858
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 19168 18737 19196 19110
rect 19154 18728 19210 18737
rect 19154 18663 19210 18672
rect 18510 17912 18566 17921
rect 18510 17847 18566 17856
rect 18420 15972 18472 15978
rect 18420 15914 18472 15920
rect 17224 15632 17276 15638
rect 17224 15574 17276 15580
rect 17408 15632 17460 15638
rect 17408 15574 17460 15580
rect 17236 15162 17264 15574
rect 17420 15473 17448 15574
rect 18432 15570 18460 15914
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18236 15496 18288 15502
rect 17406 15464 17462 15473
rect 18236 15438 18288 15444
rect 17406 15399 17462 15408
rect 17420 15162 17448 15399
rect 18050 15192 18106 15201
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17408 15156 17460 15162
rect 18248 15162 18276 15438
rect 18432 15162 18460 15506
rect 18050 15127 18106 15136
rect 18236 15156 18288 15162
rect 17408 15098 17460 15104
rect 17498 14784 17554 14793
rect 17498 14719 17554 14728
rect 17512 14618 17540 14719
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16408 13870 16436 14418
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17052 13530 17080 13806
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16578 13424 16634 13433
rect 16578 13359 16634 13368
rect 16302 13152 16358 13161
rect 16302 13087 16358 13096
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16132 12782 16160 12922
rect 16120 12776 16172 12782
rect 16026 12744 16082 12753
rect 16120 12718 16172 12724
rect 16026 12679 16082 12688
rect 15856 11206 15976 11234
rect 15750 8392 15806 8401
rect 15750 8327 15806 8336
rect 15764 6458 15792 8327
rect 15856 7834 15884 11206
rect 15934 11112 15990 11121
rect 15934 11047 15990 11056
rect 15948 10062 15976 11047
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15948 9178 15976 9998
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15856 7806 15976 7834
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15856 7274 15884 7686
rect 15844 7268 15896 7274
rect 15844 7210 15896 7216
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15764 6118 15792 6394
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15856 5642 15884 7210
rect 15948 5846 15976 7806
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 15844 5636 15896 5642
rect 15844 5578 15896 5584
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15580 4282 15608 4762
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15580 4049 15608 4218
rect 15672 4214 15700 4422
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15566 4040 15622 4049
rect 15566 3975 15622 3984
rect 15476 604 15528 610
rect 15476 546 15528 552
rect 15764 480 15792 5578
rect 15948 5370 15976 5782
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 15948 5001 15976 5306
rect 15934 4992 15990 5001
rect 15934 4927 15990 4936
rect 16040 3670 16068 12679
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 16500 11014 16528 12582
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16500 10470 16528 10950
rect 16592 10606 16620 13359
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16776 11898 16804 12242
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 17130 11792 17186 11801
rect 17130 11727 17186 11736
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16856 10532 16908 10538
rect 16856 10474 16908 10480
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 16132 9489 16160 10134
rect 16118 9480 16174 9489
rect 16118 9415 16120 9424
rect 16172 9415 16174 9424
rect 16120 9386 16172 9392
rect 16394 9208 16450 9217
rect 16394 9143 16450 9152
rect 16408 9042 16436 9143
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16132 7954 16160 8366
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 16132 7410 16160 7686
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16132 6458 16160 7346
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16212 4548 16264 4554
rect 16212 4490 16264 4496
rect 16224 3942 16252 4490
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 16028 3664 16080 3670
rect 16028 3606 16080 3612
rect 16224 3233 16252 3878
rect 16210 3224 16266 3233
rect 16210 3159 16266 3168
rect 16316 480 16344 8774
rect 16408 8634 16436 8978
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16500 8480 16528 10406
rect 16868 9722 16896 10474
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16868 9518 16896 9658
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16408 8452 16528 8480
rect 16408 7954 16436 8452
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16408 7206 16436 7890
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16408 6798 16436 7142
rect 16500 6866 16528 8298
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16592 7274 16620 7890
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16408 6168 16436 6598
rect 16500 6322 16528 6802
rect 16684 6662 16712 6802
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16776 6458 16804 7142
rect 16960 7002 16988 7142
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16488 6180 16540 6186
rect 16408 6140 16488 6168
rect 16488 6122 16540 6128
rect 16500 6089 16528 6122
rect 16486 6080 16542 6089
rect 16486 6015 16542 6024
rect 16500 5846 16528 6015
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 16408 5409 16436 5782
rect 16394 5400 16450 5409
rect 16394 5335 16396 5344
rect 16448 5335 16450 5344
rect 16396 5306 16448 5312
rect 16488 5296 16540 5302
rect 16488 5238 16540 5244
rect 16500 3670 16528 5238
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16960 4826 16988 4966
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16592 4282 16620 4490
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 16592 3534 16620 4218
rect 16684 3602 16712 4626
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16868 3942 16896 4422
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16500 2854 16528 3402
rect 16592 2990 16620 3470
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16488 2848 16540 2854
rect 16488 2790 16540 2796
rect 16500 2530 16528 2790
rect 16684 2650 16712 3538
rect 16868 3194 16896 3878
rect 16960 3738 16988 3946
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17144 3126 17172 11727
rect 18064 9586 18092 15127
rect 18236 15098 18288 15104
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18510 13968 18566 13977
rect 18510 13903 18566 13912
rect 18524 13394 18552 13903
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18524 12986 18552 13330
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17236 5234 17264 7142
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17420 5166 17448 6054
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17236 4690 17264 4966
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17420 4010 17448 4626
rect 17408 4004 17460 4010
rect 17408 3946 17460 3952
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 17512 2666 17540 9318
rect 17590 7984 17646 7993
rect 17590 7919 17646 7928
rect 17604 7546 17632 7919
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 18064 7392 18092 9522
rect 18064 7364 18184 7392
rect 18050 7304 18106 7313
rect 18050 7239 18052 7248
rect 18104 7239 18106 7248
rect 18052 7210 18104 7216
rect 18050 6760 18106 6769
rect 18050 6695 18106 6704
rect 18064 6322 18092 6695
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17880 5658 17908 5714
rect 17604 5030 17632 5646
rect 17880 5630 18000 5658
rect 17972 5166 18000 5630
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17682 4312 17738 4321
rect 17682 4247 17738 4256
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 17420 2638 17540 2666
rect 16500 2514 16620 2530
rect 16500 2508 16632 2514
rect 16500 2502 16580 2508
rect 16580 2450 16632 2456
rect 16856 604 16908 610
rect 16856 546 16908 552
rect 16868 480 16896 546
rect 17420 480 17448 2638
rect 17696 2553 17724 4247
rect 17866 3088 17922 3097
rect 18156 3058 18184 7364
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18340 6497 18368 6598
rect 18326 6488 18382 6497
rect 18326 6423 18382 6432
rect 18524 6361 18552 7142
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18510 6352 18566 6361
rect 18510 6287 18566 6296
rect 18708 5953 18736 6598
rect 18694 5944 18750 5953
rect 18694 5879 18750 5888
rect 18892 5370 18920 6734
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 18984 5914 19012 6122
rect 18972 5908 19024 5914
rect 18972 5850 19024 5856
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18602 5128 18658 5137
rect 18326 4856 18382 4865
rect 18326 4791 18382 4800
rect 18340 4010 18368 4791
rect 18524 4554 18552 5102
rect 18602 5063 18604 5072
rect 18656 5063 18658 5072
rect 18604 5034 18656 5040
rect 18512 4548 18564 4554
rect 18512 4490 18564 4496
rect 18510 4448 18566 4457
rect 18510 4383 18566 4392
rect 18328 4004 18380 4010
rect 18328 3946 18380 3952
rect 17866 3023 17922 3032
rect 18144 3052 18196 3058
rect 17880 2553 17908 3023
rect 18144 2994 18196 3000
rect 18156 2961 18184 2994
rect 18142 2952 18198 2961
rect 18142 2887 18198 2896
rect 18326 2680 18382 2689
rect 18326 2615 18382 2624
rect 17682 2544 17738 2553
rect 17682 2479 17738 2488
rect 17866 2544 17922 2553
rect 17866 2479 17922 2488
rect 18340 2378 18368 2615
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18064 2009 18092 2246
rect 18050 2000 18106 2009
rect 18050 1935 18106 1944
rect 17866 1456 17922 1465
rect 17866 1391 17922 1400
rect 17880 480 17908 1391
rect 18524 626 18552 4383
rect 19076 3602 19104 7278
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 18708 3058 18736 3538
rect 19076 3194 19104 3538
rect 19260 3482 19288 22086
rect 19536 20913 19564 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19522 20904 19578 20913
rect 19522 20839 19578 20848
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 20180 19417 20208 23462
rect 21732 23180 21784 23186
rect 21732 23122 21784 23128
rect 21744 22778 21772 23122
rect 21732 22772 21784 22778
rect 21732 22714 21784 22720
rect 21744 22545 21772 22714
rect 21730 22536 21786 22545
rect 21730 22471 21786 22480
rect 20904 21004 20956 21010
rect 20904 20946 20956 20952
rect 20916 20262 20944 20946
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20916 19990 20944 20198
rect 20904 19984 20956 19990
rect 20904 19926 20956 19932
rect 20166 19408 20222 19417
rect 20166 19343 20222 19352
rect 21548 19304 21600 19310
rect 21548 19246 21600 19252
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 21560 18290 21588 19246
rect 21548 18284 21600 18290
rect 21548 18226 21600 18232
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 21284 17649 21312 18158
rect 21270 17640 21326 17649
rect 21270 17575 21326 17584
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19444 12306 19472 13262
rect 20166 13152 20222 13161
rect 20166 13087 20222 13096
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19444 11898 19472 12242
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19522 7440 19578 7449
rect 19522 7375 19578 7384
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19352 6225 19380 6598
rect 19338 6216 19394 6225
rect 19338 6151 19394 6160
rect 19432 6112 19484 6118
rect 19430 6080 19432 6089
rect 19484 6080 19486 6089
rect 19430 6015 19486 6024
rect 19536 5914 19564 7375
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19430 5536 19486 5545
rect 19430 5471 19486 5480
rect 19444 5370 19472 5471
rect 19536 5386 19564 5850
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 19432 5364 19484 5370
rect 19536 5358 19656 5386
rect 19432 5306 19484 5312
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19536 4826 19564 5238
rect 19628 5098 19656 5358
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19996 5098 20024 5306
rect 20088 5234 20116 5510
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 19616 5092 19668 5098
rect 19616 5034 19668 5040
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 19614 4720 19670 4729
rect 19614 4655 19616 4664
rect 19668 4655 19670 4664
rect 19616 4626 19668 4632
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19444 4321 19472 4422
rect 19430 4312 19486 4321
rect 19430 4247 19486 4256
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 19260 3454 19380 3482
rect 19248 3392 19300 3398
rect 19246 3360 19248 3369
rect 19300 3360 19302 3369
rect 19246 3295 19302 3304
rect 19352 3194 19380 3454
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19352 3074 19380 3130
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 19260 3046 19380 3074
rect 18970 2952 19026 2961
rect 18970 2887 19026 2896
rect 18432 598 18552 626
rect 18432 480 18460 598
rect 18984 480 19012 2887
rect 19260 2825 19288 3046
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19246 2816 19302 2825
rect 19246 2751 19302 2760
rect 19352 2650 19380 2926
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19444 1329 19472 3946
rect 19430 1320 19486 1329
rect 19430 1255 19486 1264
rect 19536 480 19564 4218
rect 19628 4214 19656 4626
rect 19890 4584 19946 4593
rect 19890 4519 19946 4528
rect 19904 4486 19932 4519
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19616 4208 19668 4214
rect 19616 4150 19668 4156
rect 20180 4078 20208 13087
rect 20272 4282 20300 15302
rect 21836 15201 21864 23598
rect 21928 21146 21956 23718
rect 22006 23624 22062 23633
rect 22006 23559 22062 23568
rect 22020 23322 22048 23559
rect 23492 23474 23520 25162
rect 23768 23633 23796 27520
rect 24320 25226 24348 27520
rect 24308 25220 24360 25226
rect 24308 25162 24360 25168
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 23754 23624 23810 23633
rect 23754 23559 23810 23568
rect 23400 23446 23520 23474
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 21916 21140 21968 21146
rect 21916 21082 21968 21088
rect 23400 19174 23428 23446
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24872 22001 24900 27520
rect 25424 24313 25452 27520
rect 25976 25158 26004 27520
rect 25964 25152 26016 25158
rect 25964 25094 26016 25100
rect 25410 24304 25466 24313
rect 25410 24239 25466 24248
rect 26528 23225 26556 27520
rect 27080 24857 27108 27520
rect 27066 24848 27122 24857
rect 27066 24783 27122 24792
rect 26514 23216 26570 23225
rect 26514 23151 26570 23160
rect 24858 21992 24914 22001
rect 24858 21927 24914 21936
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 27632 21418 27660 27520
rect 26240 21412 26292 21418
rect 26240 21354 26292 21360
rect 27620 21412 27672 21418
rect 27620 21354 27672 21360
rect 24122 21040 24178 21049
rect 24122 20975 24178 20984
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 24136 16017 24164 20975
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24122 16008 24178 16017
rect 24122 15943 24178 15952
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 21822 15192 21878 15201
rect 24289 15184 24585 15204
rect 21822 15127 21878 15136
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 26252 13297 26280 21354
rect 26238 13288 26294 13297
rect 26238 13223 26294 13232
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 25962 12336 26018 12345
rect 25962 12271 26018 12280
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20352 5704 20404 5710
rect 20350 5672 20352 5681
rect 20404 5672 20406 5681
rect 20350 5607 20406 5616
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20260 4276 20312 4282
rect 20260 4218 20312 4224
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20076 4004 20128 4010
rect 20076 3946 20128 3952
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19616 3528 19668 3534
rect 19614 3496 19616 3505
rect 19668 3496 19670 3505
rect 19614 3431 19670 3440
rect 19628 3194 19656 3431
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19616 3188 19668 3194
rect 19616 3130 19668 3136
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19904 1601 19932 2450
rect 19996 1737 20024 3334
rect 19982 1728 20038 1737
rect 19982 1663 20038 1672
rect 19890 1592 19946 1601
rect 19890 1527 19946 1536
rect 20088 480 20116 3946
rect 20180 2922 20208 4014
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20168 2916 20220 2922
rect 20168 2858 20220 2864
rect 20180 2650 20208 2858
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 20272 649 20300 3334
rect 20364 2825 20392 3878
rect 20350 2816 20406 2825
rect 20350 2751 20406 2760
rect 20456 2514 20484 4966
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20444 2508 20496 2514
rect 20444 2450 20496 2456
rect 20548 921 20576 4558
rect 20640 4049 20668 12038
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 21362 10840 21418 10849
rect 24289 10832 24585 10852
rect 21362 10775 21418 10784
rect 20902 9480 20958 9489
rect 20902 9415 20958 9424
rect 20720 5160 20772 5166
rect 20718 5128 20720 5137
rect 20772 5128 20774 5137
rect 20718 5063 20774 5072
rect 20916 4690 20944 9415
rect 20994 5808 21050 5817
rect 20994 5743 21050 5752
rect 21008 5370 21036 5743
rect 20996 5364 21048 5370
rect 20996 5306 21048 5312
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20720 4548 20772 4554
rect 20720 4490 20772 4496
rect 20626 4040 20682 4049
rect 20626 3975 20682 3984
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20640 2650 20668 2926
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 20534 912 20590 921
rect 20534 847 20590 856
rect 20258 640 20314 649
rect 20258 575 20314 584
rect 20640 480 20668 2314
rect 20732 610 20760 4490
rect 20916 4282 20944 4626
rect 21088 4480 21140 4486
rect 21086 4448 21088 4457
rect 21140 4448 21142 4457
rect 21086 4383 21142 4392
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 21272 4072 21324 4078
rect 21272 4014 21324 4020
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20916 2854 20944 3538
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 21284 2553 21312 4014
rect 21376 3738 21404 10775
rect 22006 9888 22062 9897
rect 22006 9823 22062 9832
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 21468 4185 21496 4422
rect 21454 4176 21510 4185
rect 21454 4111 21510 4120
rect 21638 4040 21694 4049
rect 21638 3975 21694 3984
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 21376 2990 21404 3674
rect 21364 2984 21416 2990
rect 21364 2926 21416 2932
rect 21270 2544 21326 2553
rect 21270 2479 21326 2488
rect 20720 604 20772 610
rect 20720 546 20772 552
rect 21180 604 21232 610
rect 21180 546 21232 552
rect 21192 480 21220 546
rect 21652 480 21680 3975
rect 22020 3602 22048 9823
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 22466 5400 22522 5409
rect 24289 5392 24585 5412
rect 22466 5335 22522 5344
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 22008 3596 22060 3602
rect 22008 3538 22060 3544
rect 21824 3392 21876 3398
rect 21824 3334 21876 3340
rect 21836 1057 21864 3334
rect 22020 3194 22048 3538
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22204 2961 22232 3334
rect 22388 3233 22416 3878
rect 22374 3224 22430 3233
rect 22374 3159 22430 3168
rect 22190 2952 22246 2961
rect 22190 2887 22246 2896
rect 22098 2816 22154 2825
rect 22098 2751 22154 2760
rect 21822 1048 21878 1057
rect 21822 983 21878 992
rect 22112 626 22140 2751
rect 22480 2514 22508 5335
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 23662 3496 23718 3505
rect 22744 3460 22796 3466
rect 23662 3431 23718 3440
rect 22744 3402 22796 3408
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22204 785 22232 2246
rect 22190 776 22246 785
rect 22190 711 22246 720
rect 22112 598 22232 626
rect 22204 480 22232 598
rect 22756 480 22784 3402
rect 23676 3058 23704 3431
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 24858 3088 24914 3097
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 23296 2644 23348 2650
rect 23296 2586 23348 2592
rect 23308 480 23336 2586
rect 23860 480 23888 3062
rect 24858 3023 24914 3032
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 24044 1737 24072 2450
rect 24124 2372 24176 2378
rect 24124 2314 24176 2320
rect 24030 1728 24086 1737
rect 24030 1663 24086 1672
rect 24136 1170 24164 2314
rect 24216 2304 24268 2310
rect 24216 2246 24268 2252
rect 24228 1465 24256 2246
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24214 1456 24270 1465
rect 24214 1391 24270 1400
rect 24136 1142 24440 1170
rect 24412 480 24440 1142
rect 24872 480 24900 3023
rect 25410 2408 25466 2417
rect 25410 2343 25466 2352
rect 25424 480 25452 2343
rect 25976 480 26004 12271
rect 27618 6760 27674 6769
rect 27618 6695 27674 6704
rect 27066 4992 27122 5001
rect 27066 4927 27122 4936
rect 26514 3632 26570 3641
rect 26514 3567 26570 3576
rect 26528 480 26556 3567
rect 27080 480 27108 4927
rect 27632 480 27660 6695
rect 4066 368 4122 377
rect 4066 303 4122 312
rect 4434 0 4490 480
rect 4986 0 5042 480
rect 5538 0 5594 480
rect 6090 0 6146 480
rect 6642 0 6698 480
rect 7194 0 7250 480
rect 7654 0 7710 480
rect 8206 0 8262 480
rect 8758 0 8814 480
rect 9310 0 9366 480
rect 9862 0 9918 480
rect 10414 0 10470 480
rect 10874 0 10930 480
rect 11426 0 11482 480
rect 11978 0 12034 480
rect 12530 0 12586 480
rect 13082 0 13138 480
rect 13634 0 13690 480
rect 14186 0 14242 480
rect 14646 0 14702 480
rect 15198 0 15254 480
rect 15750 0 15806 480
rect 16302 0 16358 480
rect 16854 0 16910 480
rect 17406 0 17462 480
rect 17866 0 17922 480
rect 18418 0 18474 480
rect 18970 0 19026 480
rect 19522 0 19578 480
rect 20074 0 20130 480
rect 20626 0 20682 480
rect 21178 0 21234 480
rect 21638 0 21694 480
rect 22190 0 22246 480
rect 22742 0 22798 480
rect 23294 0 23350 480
rect 23846 0 23902 480
rect 24398 0 24454 480
rect 24858 0 24914 480
rect 25410 0 25466 480
rect 25962 0 26018 480
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 3238 27648 3294 27704
rect 1674 25744 1730 25800
rect 662 24248 718 24304
rect 1490 24520 1546 24576
rect 2226 26968 2282 27024
rect 1766 24656 1822 24712
rect 1398 23704 1454 23760
rect 202 23568 258 23624
rect 1950 23568 2006 23624
rect 1950 23024 2006 23080
rect 3146 24248 3202 24304
rect 2778 23160 2834 23216
rect 2318 21936 2374 21992
rect 2502 21956 2558 21992
rect 2502 21936 2504 21956
rect 2504 21936 2556 21956
rect 2556 21936 2558 21956
rect 2502 21392 2558 21448
rect 570 11192 626 11248
rect 1674 13504 1730 13560
rect 2870 22108 2872 22128
rect 2872 22108 2924 22128
rect 2924 22108 2926 22128
rect 2870 22072 2926 22108
rect 1858 17448 1914 17504
rect 1766 12960 1822 13016
rect 1582 10376 1638 10432
rect 1490 8472 1546 8528
rect 1214 7656 1270 7712
rect 662 3712 718 3768
rect 1582 7112 1638 7168
rect 1398 6160 1454 6216
rect 1398 3596 1454 3632
rect 1398 3576 1400 3596
rect 1400 3576 1452 3596
rect 1452 3576 1454 3596
rect 1766 12724 1768 12744
rect 1768 12724 1820 12744
rect 1820 12724 1822 12744
rect 1766 12688 1822 12724
rect 2686 19352 2742 19408
rect 2594 18264 2650 18320
rect 2042 15272 2098 15328
rect 2042 14320 2098 14376
rect 2226 13796 2282 13832
rect 2226 13776 2228 13796
rect 2228 13776 2280 13796
rect 2280 13776 2282 13796
rect 2134 13676 2136 13696
rect 2136 13676 2188 13696
rect 2188 13676 2190 13696
rect 2134 13640 2190 13676
rect 1950 12960 2006 13016
rect 1858 9444 1914 9480
rect 1858 9424 1860 9444
rect 1860 9424 1912 9444
rect 1912 9424 1914 9444
rect 1858 8608 1914 8664
rect 2870 18672 2926 18728
rect 3330 24384 3386 24440
rect 3698 23840 3754 23896
rect 4066 26308 4122 26344
rect 4066 26288 4068 26308
rect 4068 26288 4120 26308
rect 4120 26288 4122 26308
rect 4066 25064 4122 25120
rect 4434 24556 4436 24576
rect 4436 24556 4488 24576
rect 4488 24556 4490 24576
rect 3974 23296 4030 23352
rect 3698 23024 3754 23080
rect 4434 24520 4490 24556
rect 3974 22616 4030 22672
rect 3330 20984 3386 21040
rect 3882 22480 3938 22536
rect 3698 19760 3754 19816
rect 4250 21392 4306 21448
rect 3974 21256 4030 21312
rect 4434 20304 4490 20360
rect 4066 18672 4122 18728
rect 4066 18128 4122 18184
rect 3974 17856 4030 17912
rect 2870 12860 2872 12880
rect 2872 12860 2924 12880
rect 2924 12860 2926 12880
rect 2870 12824 2926 12860
rect 2686 11736 2742 11792
rect 1766 6024 1822 6080
rect 1950 5072 2006 5128
rect 2134 6432 2190 6488
rect 2318 5888 2374 5944
rect 2686 11464 2742 11520
rect 3146 11600 3202 11656
rect 2502 6976 2558 7032
rect 2962 8880 3018 8936
rect 2870 7792 2926 7848
rect 2962 6024 3018 6080
rect 3514 9036 3570 9072
rect 3514 9016 3516 9036
rect 3516 9016 3568 9036
rect 3568 9016 3570 9036
rect 3422 8336 3478 8392
rect 3974 15816 4030 15872
rect 4710 23704 4766 23760
rect 4986 23604 4988 23624
rect 4988 23604 5040 23624
rect 5040 23604 5042 23624
rect 4986 23568 5042 23604
rect 4986 22480 5042 22536
rect 4434 15564 4490 15600
rect 4434 15544 4436 15564
rect 4436 15544 4488 15564
rect 4488 15544 4490 15564
rect 3974 13368 4030 13424
rect 4158 13252 4214 13288
rect 4158 13232 4160 13252
rect 4160 13232 4212 13252
rect 4212 13232 4214 13252
rect 3974 12144 4030 12200
rect 4434 12316 4436 12336
rect 4436 12316 4488 12336
rect 4488 12316 4490 12336
rect 4434 12280 4490 12316
rect 4342 11500 4344 11520
rect 4344 11500 4396 11520
rect 4396 11500 4398 11520
rect 4342 11464 4398 11500
rect 3974 10648 4030 10704
rect 3790 10240 3846 10296
rect 3698 8472 3754 8528
rect 3238 6976 3294 7032
rect 2778 5480 2834 5536
rect 2502 4548 2558 4584
rect 2502 4528 2504 4548
rect 2504 4528 2556 4548
rect 2556 4528 2558 4548
rect 2686 5072 2742 5128
rect 2594 4256 2650 4312
rect 2594 3884 2596 3904
rect 2596 3884 2648 3904
rect 2648 3884 2650 3904
rect 2594 3848 2650 3884
rect 2502 3340 2504 3360
rect 2504 3340 2556 3360
rect 2556 3340 2558 3360
rect 2502 3304 2558 3340
rect 2318 3068 2320 3088
rect 2320 3068 2372 3088
rect 2372 3068 2374 3088
rect 2318 3032 2374 3068
rect 2042 2896 2098 2952
rect 1582 2216 1638 2272
rect 1398 1536 1454 1592
rect 2502 1672 2558 1728
rect 2870 2624 2926 2680
rect 2594 584 2650 640
rect 3238 5072 3294 5128
rect 3330 2352 3386 2408
rect 3146 2216 3202 2272
rect 3330 1536 3386 1592
rect 3514 7384 3570 7440
rect 3514 7112 3570 7168
rect 3698 7112 3754 7168
rect 3606 6860 3662 6896
rect 3606 6840 3608 6860
rect 3608 6840 3660 6860
rect 3660 6840 3662 6860
rect 3698 6704 3754 6760
rect 3790 6568 3846 6624
rect 3514 3440 3570 3496
rect 3514 2624 3570 2680
rect 4066 9968 4122 10024
rect 3974 9152 4030 9208
rect 4066 7928 4122 7984
rect 4158 6704 4214 6760
rect 4066 5616 4122 5672
rect 4894 15272 4950 15328
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5906 23740 5908 23760
rect 5908 23740 5960 23760
rect 5960 23740 5962 23760
rect 5906 23704 5962 23740
rect 5906 23296 5962 23352
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 6274 24656 6330 24712
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5630 19252 5632 19272
rect 5632 19252 5684 19272
rect 5684 19252 5686 19272
rect 5630 19216 5686 19252
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 6182 18264 6238 18320
rect 6366 18300 6368 18320
rect 6368 18300 6420 18320
rect 6420 18300 6422 18320
rect 6366 18264 6422 18300
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5262 16124 5264 16144
rect 5264 16124 5316 16144
rect 5316 16124 5318 16144
rect 5262 16088 5318 16124
rect 6274 16768 6330 16824
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5998 16224 6054 16280
rect 6182 15852 6184 15872
rect 6184 15852 6236 15872
rect 6236 15852 6238 15872
rect 6182 15816 6238 15852
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 4802 11772 4804 11792
rect 4804 11772 4856 11792
rect 4856 11772 4858 11792
rect 4802 11736 4858 11772
rect 4802 11600 4858 11656
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5538 12416 5594 12472
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6458 13912 6514 13968
rect 6090 11056 6146 11112
rect 5998 10956 6000 10976
rect 6000 10956 6052 10976
rect 6052 10956 6054 10976
rect 5998 10920 6054 10956
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5630 10512 5686 10568
rect 4894 9832 4950 9888
rect 4986 9152 5042 9208
rect 4986 8608 5042 8664
rect 4802 7792 4858 7848
rect 5538 10376 5594 10432
rect 5722 10240 5778 10296
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5354 8336 5410 8392
rect 5262 7692 5264 7712
rect 5264 7692 5316 7712
rect 5316 7692 5318 7712
rect 5262 7656 5318 7692
rect 6642 22888 6698 22944
rect 6642 22616 6698 22672
rect 6918 23296 6974 23352
rect 6826 21392 6882 21448
rect 7654 23160 7710 23216
rect 6550 12552 6606 12608
rect 6458 11348 6514 11384
rect 6458 11328 6460 11348
rect 6460 11328 6512 11348
rect 6512 11328 6514 11348
rect 6734 13796 6790 13832
rect 6734 13776 6736 13796
rect 6736 13776 6788 13796
rect 6788 13776 6790 13796
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5170 6704 5226 6760
rect 5078 6432 5134 6488
rect 4802 6024 4858 6080
rect 4618 5788 4620 5808
rect 4620 5788 4672 5808
rect 4672 5788 4674 5808
rect 4618 5752 4674 5788
rect 4158 5092 4214 5128
rect 4158 5072 4160 5092
rect 4160 5072 4212 5092
rect 4212 5072 4214 5092
rect 3882 4664 3938 4720
rect 3974 4528 4030 4584
rect 3790 1944 3846 2000
rect 3606 1536 3662 1592
rect 4158 3304 4214 3360
rect 4066 1400 4122 1456
rect 3974 1128 4030 1184
rect 4158 720 4214 776
rect 4618 5072 4674 5128
rect 4618 3032 4674 3088
rect 4526 1808 4582 1864
rect 5078 6024 5134 6080
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5446 4664 5502 4720
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5446 4256 5502 4312
rect 4618 992 4674 1048
rect 5354 2216 5410 2272
rect 6182 7520 6238 7576
rect 6642 9832 6698 9888
rect 7562 20576 7618 20632
rect 7654 17604 7710 17640
rect 7654 17584 7656 17604
rect 7656 17584 7708 17604
rect 7708 17584 7710 17604
rect 7930 17312 7986 17368
rect 7378 15972 7434 16008
rect 7378 15952 7380 15972
rect 7380 15952 7432 15972
rect 7432 15952 7434 15972
rect 7470 13524 7526 13560
rect 7470 13504 7472 13524
rect 7472 13504 7524 13524
rect 7524 13504 7526 13524
rect 7378 12960 7434 13016
rect 7378 11736 7434 11792
rect 7470 10784 7526 10840
rect 7746 10784 7802 10840
rect 7194 9288 7250 9344
rect 7286 8608 7342 8664
rect 7010 8064 7066 8120
rect 7286 8064 7342 8120
rect 7286 7656 7342 7712
rect 6090 5344 6146 5400
rect 6366 6296 6422 6352
rect 6182 3712 6238 3768
rect 5722 3576 5778 3632
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6182 3168 6238 3224
rect 5998 2216 6054 2272
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6090 1536 6146 1592
rect 7010 6976 7066 7032
rect 6918 6160 6974 6216
rect 6458 4020 6460 4040
rect 6460 4020 6512 4040
rect 6512 4020 6514 4040
rect 6458 3984 6514 4020
rect 6550 2932 6552 2952
rect 6552 2932 6604 2952
rect 6604 2932 6606 2952
rect 6550 2896 6606 2932
rect 6274 1264 6330 1320
rect 6826 5752 6882 5808
rect 6734 5344 6790 5400
rect 7654 9696 7710 9752
rect 7654 9288 7710 9344
rect 7562 8200 7618 8256
rect 7378 7112 7434 7168
rect 7378 6296 7434 6352
rect 7194 6180 7250 6216
rect 7194 6160 7196 6180
rect 7196 6160 7248 6180
rect 7248 6160 7250 6180
rect 7102 3848 7158 3904
rect 7286 5908 7342 5944
rect 7286 5888 7288 5908
rect 7288 5888 7340 5908
rect 7340 5888 7342 5908
rect 8574 22752 8630 22808
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 9678 24248 9734 24304
rect 9494 23840 9550 23896
rect 9218 23024 9274 23080
rect 9126 21800 9182 21856
rect 8942 20712 8998 20768
rect 8022 16768 8078 16824
rect 10046 23316 10102 23352
rect 10046 23296 10048 23316
rect 10048 23296 10100 23316
rect 10100 23296 10102 23316
rect 9218 18536 9274 18592
rect 9310 18400 9366 18456
rect 8758 17856 8814 17912
rect 8298 15564 8354 15600
rect 8298 15544 8300 15564
rect 8300 15544 8352 15564
rect 8352 15544 8354 15564
rect 8758 15272 8814 15328
rect 9402 17856 9458 17912
rect 9494 17040 9550 17096
rect 8022 10376 8078 10432
rect 8390 9560 8446 9616
rect 9218 14864 9274 14920
rect 9402 13776 9458 13832
rect 9770 18128 9826 18184
rect 9678 16904 9734 16960
rect 9586 13640 9642 13696
rect 8574 10784 8630 10840
rect 8390 7248 8446 7304
rect 8298 6740 8300 6760
rect 8300 6740 8352 6760
rect 8352 6740 8354 6760
rect 8298 6704 8354 6740
rect 8022 6568 8078 6624
rect 7838 5636 7894 5672
rect 7838 5616 7840 5636
rect 7840 5616 7892 5636
rect 7892 5616 7894 5636
rect 8022 5616 8078 5672
rect 8298 3848 8354 3904
rect 7654 3712 7710 3768
rect 8206 3576 8262 3632
rect 7838 3440 7894 3496
rect 9034 12144 9090 12200
rect 9034 10104 9090 10160
rect 8758 6840 8814 6896
rect 8574 2760 8630 2816
rect 8390 2624 8446 2680
rect 9310 12144 9366 12200
rect 9954 17312 10010 17368
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10598 23160 10654 23216
rect 10690 22480 10746 22536
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10874 21936 10930 21992
rect 10782 20304 10838 20360
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10598 19760 10654 19816
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 11058 24248 11114 24304
rect 11426 24792 11482 24848
rect 11518 23296 11574 23352
rect 11518 22072 11574 22128
rect 11518 20712 11574 20768
rect 11334 20440 11390 20496
rect 11150 19080 11206 19136
rect 11242 18844 11244 18864
rect 11244 18844 11296 18864
rect 11296 18844 11298 18864
rect 11242 18808 11298 18844
rect 11426 19760 11482 19816
rect 10046 16904 10102 16960
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10138 16632 10194 16688
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10138 13912 10194 13968
rect 10138 13640 10194 13696
rect 9770 11076 9826 11112
rect 9770 11056 9772 11076
rect 9772 11056 9824 11076
rect 9824 11056 9826 11076
rect 9954 11328 10010 11384
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10874 17856 10930 17912
rect 10782 14184 10838 14240
rect 10874 13948 10876 13968
rect 10876 13948 10928 13968
rect 10928 13948 10930 13968
rect 10874 13912 10930 13948
rect 10690 12300 10746 12336
rect 10690 12280 10692 12300
rect 10692 12280 10744 12300
rect 10744 12280 10746 12300
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 9862 10920 9918 10976
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 9862 9968 9918 10024
rect 9218 9832 9274 9888
rect 9678 9424 9734 9480
rect 9310 8492 9366 8528
rect 9310 8472 9312 8492
rect 9312 8472 9364 8492
rect 9364 8472 9366 8492
rect 9494 8472 9550 8528
rect 9770 8336 9826 8392
rect 9034 3440 9090 3496
rect 9494 7268 9550 7304
rect 9494 7248 9496 7268
rect 9496 7248 9548 7268
rect 9548 7248 9550 7268
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10322 8336 10378 8392
rect 10138 8200 10194 8256
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 9770 5752 9826 5808
rect 9678 5616 9734 5672
rect 9954 5772 10010 5808
rect 9954 5752 9956 5772
rect 9956 5752 10008 5772
rect 10008 5752 10010 5772
rect 9310 3304 9366 3360
rect 9310 3032 9366 3088
rect 9678 3848 9734 3904
rect 10782 7420 10784 7440
rect 10784 7420 10836 7440
rect 10836 7420 10838 7440
rect 10782 7384 10838 7420
rect 10690 7112 10746 7168
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 11150 15308 11152 15328
rect 11152 15308 11204 15328
rect 11204 15308 11206 15328
rect 11150 15272 11206 15308
rect 11610 16224 11666 16280
rect 11610 15816 11666 15872
rect 11518 15680 11574 15736
rect 11794 22752 11850 22808
rect 12070 23024 12126 23080
rect 11886 18264 11942 18320
rect 11978 15952 12034 16008
rect 11610 12960 11666 13016
rect 11610 12552 11666 12608
rect 11794 13096 11850 13152
rect 11794 12824 11850 12880
rect 11886 12552 11942 12608
rect 11886 12280 11942 12336
rect 11518 11600 11574 11656
rect 11518 10920 11574 10976
rect 11150 9016 11206 9072
rect 10966 6860 11022 6896
rect 10966 6840 10968 6860
rect 10968 6840 11020 6860
rect 11020 6840 11022 6860
rect 10138 6024 10194 6080
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 11242 6568 11298 6624
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10874 4800 10930 4856
rect 11794 9832 11850 9888
rect 11886 9560 11942 9616
rect 11610 8200 11666 8256
rect 11610 7656 11666 7712
rect 12530 21936 12586 21992
rect 12346 21664 12402 21720
rect 12622 21800 12678 21856
rect 12530 20476 12532 20496
rect 12532 20476 12584 20496
rect 12584 20476 12586 20496
rect 12530 20440 12586 20476
rect 12990 20848 13046 20904
rect 12530 19216 12586 19272
rect 13450 20984 13506 21040
rect 13082 18284 13138 18320
rect 13082 18264 13084 18284
rect 13084 18264 13136 18284
rect 13136 18264 13138 18284
rect 13174 17856 13230 17912
rect 12806 16632 12862 16688
rect 13358 16088 13414 16144
rect 12898 14184 12954 14240
rect 12622 13776 12678 13832
rect 12254 12416 12310 12472
rect 12806 13368 12862 13424
rect 12898 13096 12954 13152
rect 12714 12280 12770 12336
rect 12990 12280 13046 12336
rect 12714 11736 12770 11792
rect 12714 11056 12770 11112
rect 12530 10784 12586 10840
rect 12346 9832 12402 9888
rect 12346 9560 12402 9616
rect 12898 10648 12954 10704
rect 12346 8880 12402 8936
rect 11886 6060 11888 6080
rect 11888 6060 11940 6080
rect 11940 6060 11942 6080
rect 11886 6024 11942 6060
rect 11518 5480 11574 5536
rect 11518 5344 11574 5400
rect 11518 5208 11574 5264
rect 11794 5208 11850 5264
rect 10046 2488 10102 2544
rect 10046 1128 10102 1184
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11334 4256 11390 4312
rect 11518 4256 11574 4312
rect 11426 2896 11482 2952
rect 10874 2760 10930 2816
rect 10782 2352 10838 2408
rect 9678 856 9734 912
rect 10046 720 10102 776
rect 11150 2508 11206 2544
rect 11150 2488 11152 2508
rect 11152 2488 11204 2508
rect 11204 2488 11206 2508
rect 12162 5480 12218 5536
rect 11518 1400 11574 1456
rect 13450 15272 13506 15328
rect 13174 12144 13230 12200
rect 13266 11076 13322 11112
rect 13266 11056 13268 11076
rect 13268 11056 13320 11076
rect 13320 11056 13322 11076
rect 13634 23568 13690 23624
rect 13634 22888 13690 22944
rect 13818 22480 13874 22536
rect 13726 22208 13782 22264
rect 14278 23160 14334 23216
rect 14186 21020 14188 21040
rect 14188 21020 14240 21040
rect 14240 21020 14242 21040
rect 14186 20984 14242 21020
rect 13818 19916 13874 19952
rect 13818 19896 13820 19916
rect 13820 19896 13872 19916
rect 13872 19896 13874 19916
rect 13726 19352 13782 19408
rect 13634 19216 13690 19272
rect 13818 15700 13874 15736
rect 13818 15680 13820 15700
rect 13820 15680 13872 15700
rect 13872 15680 13874 15700
rect 14186 16496 14242 16552
rect 14094 15952 14150 16008
rect 14278 15680 14334 15736
rect 14554 23840 14610 23896
rect 14462 23296 14518 23352
rect 14186 13232 14242 13288
rect 13082 9560 13138 9616
rect 13450 9560 13506 9616
rect 13082 8880 13138 8936
rect 12714 7112 12770 7168
rect 12438 4800 12494 4856
rect 12622 4256 12678 4312
rect 12438 3304 12494 3360
rect 12438 3032 12494 3088
rect 12714 3576 12770 3632
rect 12714 3304 12770 3360
rect 12990 8336 13046 8392
rect 13082 4936 13138 4992
rect 13266 3612 13268 3632
rect 13268 3612 13320 3632
rect 13320 3612 13322 3632
rect 13266 3576 13322 3612
rect 13358 3460 13414 3496
rect 13358 3440 13360 3460
rect 13360 3440 13412 3460
rect 13412 3440 13414 3460
rect 14002 9152 14058 9208
rect 14646 22344 14702 22400
rect 14646 20576 14702 20632
rect 14738 18536 14794 18592
rect 14554 14764 14556 14784
rect 14556 14764 14608 14784
rect 14608 14764 14610 14784
rect 14554 14728 14610 14764
rect 14186 9696 14242 9752
rect 14186 7520 14242 7576
rect 14002 6024 14058 6080
rect 13542 5344 13598 5400
rect 13634 5208 13690 5264
rect 13174 1536 13230 1592
rect 14462 9594 14518 9650
rect 14278 4664 14334 4720
rect 14554 5888 14610 5944
rect 14278 3168 14334 3224
rect 13818 2624 13874 2680
rect 14186 2488 14242 2544
rect 14370 2372 14426 2408
rect 14370 2352 14372 2372
rect 14372 2352 14424 2372
rect 14424 2352 14426 2372
rect 14646 5480 14702 5536
rect 14646 4664 14702 4720
rect 14554 2216 14610 2272
rect 14186 1944 14242 2000
rect 14646 1944 14702 2000
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15566 24248 15622 24304
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15934 23196 15936 23216
rect 15936 23196 15988 23216
rect 15988 23196 15990 23216
rect 15934 23160 15990 23196
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 16026 22380 16028 22400
rect 16028 22380 16080 22400
rect 16080 22380 16082 22400
rect 16026 22344 16082 22380
rect 15842 22228 15898 22264
rect 15842 22208 15844 22228
rect 15844 22208 15896 22228
rect 15896 22208 15898 22228
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15382 20984 15438 21040
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15290 19252 15292 19272
rect 15292 19252 15344 19272
rect 15344 19252 15346 19272
rect 15290 19216 15346 19252
rect 15290 19080 15346 19136
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15934 19760 15990 19816
rect 15474 19352 15530 19408
rect 15658 18828 15714 18864
rect 15658 18808 15660 18828
rect 15660 18808 15712 18828
rect 15712 18808 15714 18828
rect 15382 18148 15438 18184
rect 15382 18128 15384 18148
rect 15384 18128 15436 18148
rect 15436 18128 15438 18148
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 17406 24384 17462 24440
rect 17682 24404 17738 24440
rect 17682 24384 17684 24404
rect 17684 24384 17736 24404
rect 17736 24384 17738 24404
rect 16854 23604 16856 23624
rect 16856 23604 16908 23624
rect 16908 23604 16910 23624
rect 16854 23568 16910 23604
rect 18326 24656 18382 24712
rect 17958 23180 18014 23216
rect 17958 23160 17960 23180
rect 17960 23160 18012 23180
rect 18012 23160 18014 23180
rect 17038 21956 17094 21992
rect 17038 21936 17040 21956
rect 17040 21936 17092 21956
rect 17092 21936 17094 21956
rect 18786 24384 18842 24440
rect 18694 23860 18750 23896
rect 18694 23840 18696 23860
rect 18696 23840 18748 23860
rect 18748 23840 18750 23860
rect 16762 21392 16818 21448
rect 18050 20440 18106 20496
rect 17222 19896 17278 19952
rect 15842 17856 15898 17912
rect 15842 17040 15898 17096
rect 15290 16496 15346 16552
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14922 13368 14978 13424
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15382 12416 15438 12472
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 16302 19352 16358 19408
rect 16118 18264 16174 18320
rect 16670 16632 16726 16688
rect 16302 16088 16358 16144
rect 16302 15816 16358 15872
rect 15750 13232 15806 13288
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15842 12280 15898 12336
rect 15382 10104 15438 10160
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15566 9868 15568 9888
rect 15568 9868 15620 9888
rect 15620 9868 15622 9888
rect 15566 9832 15622 9868
rect 14830 9560 14886 9616
rect 15198 8880 15254 8936
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14922 7828 14924 7848
rect 14924 7828 14976 7848
rect 14976 7828 14978 7848
rect 14922 7792 14978 7828
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14830 3440 14886 3496
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 14738 1536 14794 1592
rect 15382 8472 15438 8528
rect 15474 7384 15530 7440
rect 15566 6840 15622 6896
rect 15382 5480 15438 5536
rect 17590 19780 17646 19816
rect 17590 19760 17592 19780
rect 17592 19760 17644 19780
rect 17644 19760 17646 19780
rect 19062 23432 19118 23488
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19522 24656 19578 24712
rect 19982 24656 20038 24712
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20442 23840 20498 23896
rect 21546 24656 21602 24712
rect 22006 23860 22062 23896
rect 22006 23840 22008 23860
rect 22008 23840 22060 23860
rect 22060 23840 22062 23860
rect 23202 23840 23258 23896
rect 20718 23604 20720 23624
rect 20720 23604 20772 23624
rect 20772 23604 20774 23624
rect 20718 23568 20774 23604
rect 19154 18672 19210 18728
rect 18510 17856 18566 17912
rect 17406 15408 17462 15464
rect 18050 15136 18106 15192
rect 17498 14728 17554 14784
rect 16578 13368 16634 13424
rect 16302 13096 16358 13152
rect 16026 12688 16082 12744
rect 15750 8336 15806 8392
rect 15934 11056 15990 11112
rect 15566 3984 15622 4040
rect 15934 4936 15990 4992
rect 17130 11736 17186 11792
rect 16118 9444 16174 9480
rect 16118 9424 16120 9444
rect 16120 9424 16172 9444
rect 16172 9424 16174 9444
rect 16394 9152 16450 9208
rect 16210 3168 16266 3224
rect 16486 6024 16542 6080
rect 16394 5364 16450 5400
rect 16394 5344 16396 5364
rect 16396 5344 16448 5364
rect 16448 5344 16450 5364
rect 18510 13912 18566 13968
rect 17590 7928 17646 7984
rect 18050 7268 18106 7304
rect 18050 7248 18052 7268
rect 18052 7248 18104 7268
rect 18104 7248 18106 7268
rect 18050 6704 18106 6760
rect 17682 4256 17738 4312
rect 17866 3032 17922 3088
rect 18326 6432 18382 6488
rect 18510 6296 18566 6352
rect 18694 5888 18750 5944
rect 18326 4800 18382 4856
rect 18602 5092 18658 5128
rect 18602 5072 18604 5092
rect 18604 5072 18656 5092
rect 18656 5072 18658 5092
rect 18510 4392 18566 4448
rect 18142 2896 18198 2952
rect 18326 2624 18382 2680
rect 17682 2488 17738 2544
rect 17866 2488 17922 2544
rect 18050 1944 18106 2000
rect 17866 1400 17922 1456
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19522 20848 19578 20904
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 21730 22480 21786 22536
rect 20166 19352 20222 19408
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 21270 17584 21326 17640
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 20166 13096 20222 13152
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19522 7384 19578 7440
rect 19338 6160 19394 6216
rect 19430 6060 19432 6080
rect 19432 6060 19484 6080
rect 19484 6060 19486 6080
rect 19430 6024 19486 6060
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19430 5480 19486 5536
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19614 4684 19670 4720
rect 19614 4664 19616 4684
rect 19616 4664 19668 4684
rect 19668 4664 19670 4684
rect 19430 4256 19486 4312
rect 19246 3340 19248 3360
rect 19248 3340 19300 3360
rect 19300 3340 19302 3360
rect 19246 3304 19302 3340
rect 18970 2896 19026 2952
rect 19246 2760 19302 2816
rect 19430 1264 19486 1320
rect 19890 4528 19946 4584
rect 22006 23568 22062 23624
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 23754 23568 23810 23624
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 25410 24248 25466 24304
rect 27066 24792 27122 24848
rect 26514 23160 26570 23216
rect 24858 21936 24914 21992
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24122 20984 24178 21040
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24122 15952 24178 16008
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 21822 15136 21878 15192
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 26238 13232 26294 13288
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 25962 12280 26018 12336
rect 20350 5652 20352 5672
rect 20352 5652 20404 5672
rect 20404 5652 20406 5672
rect 20350 5616 20406 5652
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19614 3476 19616 3496
rect 19616 3476 19668 3496
rect 19668 3476 19670 3496
rect 19614 3440 19670 3476
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 19982 1672 20038 1728
rect 19890 1536 19946 1592
rect 20350 2760 20406 2816
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 21362 10784 21418 10840
rect 20902 9424 20958 9480
rect 20718 5108 20720 5128
rect 20720 5108 20772 5128
rect 20772 5108 20774 5128
rect 20718 5072 20774 5108
rect 20994 5752 21050 5808
rect 20626 3984 20682 4040
rect 20534 856 20590 912
rect 20258 584 20314 640
rect 21086 4428 21088 4448
rect 21088 4428 21140 4448
rect 21140 4428 21142 4448
rect 21086 4392 21142 4428
rect 22006 9832 22062 9888
rect 21454 4120 21510 4176
rect 21638 3984 21694 4040
rect 21270 2488 21326 2544
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 22466 5344 22522 5400
rect 22374 3168 22430 3224
rect 22190 2896 22246 2952
rect 22098 2760 22154 2816
rect 21822 992 21878 1048
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 23662 3440 23718 3496
rect 22190 720 22246 776
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24858 3032 24914 3088
rect 24030 1672 24086 1728
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24214 1400 24270 1456
rect 25410 2352 25466 2408
rect 27618 6704 27674 6760
rect 27066 4936 27122 4992
rect 26514 3576 26570 3632
rect 4066 312 4122 368
<< metal3 >>
rect 0 27706 480 27736
rect 3233 27706 3299 27709
rect 0 27704 3299 27706
rect 0 27648 3238 27704
rect 3294 27648 3299 27704
rect 0 27646 3299 27648
rect 0 27616 480 27646
rect 3233 27643 3299 27646
rect 0 27026 480 27056
rect 2221 27026 2287 27029
rect 0 27024 2287 27026
rect 0 26968 2226 27024
rect 2282 26968 2287 27024
rect 0 26966 2287 26968
rect 0 26936 480 26966
rect 2221 26963 2287 26966
rect 0 26346 480 26376
rect 4061 26346 4127 26349
rect 0 26344 4127 26346
rect 0 26288 4066 26344
rect 4122 26288 4127 26344
rect 0 26286 4127 26288
rect 0 26256 480 26286
rect 4061 26283 4127 26286
rect 0 25802 480 25832
rect 1669 25802 1735 25805
rect 0 25800 1735 25802
rect 0 25744 1674 25800
rect 1730 25744 1735 25800
rect 0 25742 1735 25744
rect 0 25712 480 25742
rect 1669 25739 1735 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25122 480 25152
rect 4061 25122 4127 25125
rect 0 25120 4127 25122
rect 0 25064 4066 25120
rect 4122 25064 4127 25120
rect 0 25062 4127 25064
rect 0 25032 480 25062
rect 4061 25059 4127 25062
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 11421 24850 11487 24853
rect 27061 24850 27127 24853
rect 11421 24848 27127 24850
rect 11421 24792 11426 24848
rect 11482 24792 27066 24848
rect 27122 24792 27127 24848
rect 11421 24790 27127 24792
rect 11421 24787 11487 24790
rect 27061 24787 27127 24790
rect 1761 24714 1827 24717
rect 6269 24714 6335 24717
rect 1761 24712 6335 24714
rect 1761 24656 1766 24712
rect 1822 24656 6274 24712
rect 6330 24656 6335 24712
rect 1761 24654 6335 24656
rect 1761 24651 1827 24654
rect 6269 24651 6335 24654
rect 18321 24714 18387 24717
rect 19517 24714 19583 24717
rect 18321 24712 19583 24714
rect 18321 24656 18326 24712
rect 18382 24656 19522 24712
rect 19578 24656 19583 24712
rect 18321 24654 19583 24656
rect 18321 24651 18387 24654
rect 19517 24651 19583 24654
rect 19977 24714 20043 24717
rect 21541 24714 21607 24717
rect 19977 24712 21607 24714
rect 19977 24656 19982 24712
rect 20038 24656 21546 24712
rect 21602 24656 21607 24712
rect 19977 24654 21607 24656
rect 19977 24651 20043 24654
rect 21541 24651 21607 24654
rect 1485 24578 1551 24581
rect 4429 24578 4495 24581
rect 1485 24576 4495 24578
rect 1485 24520 1490 24576
rect 1546 24520 4434 24576
rect 4490 24520 4495 24576
rect 1485 24518 4495 24520
rect 1485 24515 1551 24518
rect 4429 24515 4495 24518
rect 10277 24512 10597 24513
rect 0 24442 480 24472
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 3325 24442 3391 24445
rect 17401 24442 17467 24445
rect 0 24440 3391 24442
rect 0 24384 3330 24440
rect 3386 24384 3391 24440
rect 0 24382 3391 24384
rect 0 24352 480 24382
rect 3325 24379 3391 24382
rect 11102 24440 17467 24442
rect 11102 24384 17406 24440
rect 17462 24384 17467 24440
rect 11102 24382 17467 24384
rect 11102 24309 11162 24382
rect 17401 24379 17467 24382
rect 17677 24442 17743 24445
rect 18781 24442 18847 24445
rect 17677 24440 18847 24442
rect 17677 24384 17682 24440
rect 17738 24384 18786 24440
rect 18842 24384 18847 24440
rect 17677 24382 18847 24384
rect 17677 24379 17743 24382
rect 18781 24379 18847 24382
rect 657 24306 723 24309
rect 3141 24306 3207 24309
rect 657 24304 3207 24306
rect 657 24248 662 24304
rect 718 24248 3146 24304
rect 3202 24248 3207 24304
rect 657 24246 3207 24248
rect 657 24243 723 24246
rect 3141 24243 3207 24246
rect 9673 24306 9739 24309
rect 11053 24306 11162 24309
rect 9673 24304 11162 24306
rect 9673 24248 9678 24304
rect 9734 24248 11058 24304
rect 11114 24248 11162 24304
rect 9673 24246 11162 24248
rect 15561 24306 15627 24309
rect 25405 24306 25471 24309
rect 15561 24304 25471 24306
rect 15561 24248 15566 24304
rect 15622 24248 25410 24304
rect 25466 24248 25471 24304
rect 15561 24246 25471 24248
rect 9673 24243 9739 24246
rect 11053 24243 11119 24246
rect 15561 24243 15627 24246
rect 25405 24243 25471 24246
rect 5610 23968 5930 23969
rect 0 23898 480 23928
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 3693 23898 3759 23901
rect 0 23896 3759 23898
rect 0 23840 3698 23896
rect 3754 23840 3759 23896
rect 0 23838 3759 23840
rect 0 23808 480 23838
rect 3693 23835 3759 23838
rect 9489 23898 9555 23901
rect 14549 23898 14615 23901
rect 9489 23896 14615 23898
rect 9489 23840 9494 23896
rect 9550 23840 14554 23896
rect 14610 23840 14615 23896
rect 9489 23838 14615 23840
rect 9489 23835 9555 23838
rect 14549 23835 14615 23838
rect 18689 23898 18755 23901
rect 20437 23898 20503 23901
rect 18689 23896 20503 23898
rect 18689 23840 18694 23896
rect 18750 23840 20442 23896
rect 20498 23840 20503 23896
rect 18689 23838 20503 23840
rect 18689 23835 18755 23838
rect 20437 23835 20503 23838
rect 22001 23898 22067 23901
rect 23197 23898 23263 23901
rect 22001 23896 23263 23898
rect 22001 23840 22006 23896
rect 22062 23840 23202 23896
rect 23258 23840 23263 23896
rect 22001 23838 23263 23840
rect 22001 23835 22067 23838
rect 23197 23835 23263 23838
rect 1393 23762 1459 23765
rect 4705 23762 4771 23765
rect 5901 23762 5967 23765
rect 1393 23760 5967 23762
rect 1393 23704 1398 23760
rect 1454 23704 4710 23760
rect 4766 23704 5906 23760
rect 5962 23704 5967 23760
rect 1393 23702 5967 23704
rect 1393 23699 1459 23702
rect 4705 23699 4771 23702
rect 5901 23699 5967 23702
rect 197 23626 263 23629
rect 1945 23626 2011 23629
rect 197 23624 2011 23626
rect 197 23568 202 23624
rect 258 23568 1950 23624
rect 2006 23568 2011 23624
rect 197 23566 2011 23568
rect 197 23563 263 23566
rect 1945 23563 2011 23566
rect 4981 23626 5047 23629
rect 13629 23626 13695 23629
rect 16849 23626 16915 23629
rect 20713 23626 20779 23629
rect 4981 23624 13554 23626
rect 4981 23568 4986 23624
rect 5042 23568 13554 23624
rect 4981 23566 13554 23568
rect 4981 23563 5047 23566
rect 13494 23490 13554 23566
rect 13629 23624 16915 23626
rect 13629 23568 13634 23624
rect 13690 23568 16854 23624
rect 16910 23568 16915 23624
rect 13629 23566 16915 23568
rect 13629 23563 13695 23566
rect 16849 23563 16915 23566
rect 19382 23624 20779 23626
rect 19382 23568 20718 23624
rect 20774 23568 20779 23624
rect 19382 23566 20779 23568
rect 19057 23490 19123 23493
rect 19382 23490 19442 23566
rect 20713 23563 20779 23566
rect 22001 23626 22067 23629
rect 23749 23626 23815 23629
rect 22001 23624 23815 23626
rect 22001 23568 22006 23624
rect 22062 23568 23754 23624
rect 23810 23568 23815 23624
rect 22001 23566 23815 23568
rect 22001 23563 22067 23566
rect 23749 23563 23815 23566
rect 13494 23488 19442 23490
rect 13494 23432 19062 23488
rect 19118 23432 19442 23488
rect 13494 23430 19442 23432
rect 19057 23427 19123 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 3969 23354 4035 23357
rect 5901 23354 5967 23357
rect 3969 23352 5967 23354
rect 3969 23296 3974 23352
rect 4030 23296 5906 23352
rect 5962 23296 5967 23352
rect 3969 23294 5967 23296
rect 3969 23291 4035 23294
rect 5901 23291 5967 23294
rect 6913 23354 6979 23357
rect 10041 23354 10107 23357
rect 6913 23352 10107 23354
rect 6913 23296 6918 23352
rect 6974 23296 10046 23352
rect 10102 23296 10107 23352
rect 6913 23294 10107 23296
rect 6913 23291 6979 23294
rect 10041 23291 10107 23294
rect 11513 23354 11579 23357
rect 14457 23354 14523 23357
rect 11513 23352 18154 23354
rect 11513 23296 11518 23352
rect 11574 23296 14462 23352
rect 14518 23296 18154 23352
rect 11513 23294 18154 23296
rect 11513 23291 11579 23294
rect 14457 23291 14523 23294
rect 0 23218 480 23248
rect 2773 23218 2839 23221
rect 7649 23218 7715 23221
rect 10593 23218 10659 23221
rect 14273 23218 14339 23221
rect 0 23216 2839 23218
rect 0 23160 2778 23216
rect 2834 23160 2839 23216
rect 0 23158 2839 23160
rect 0 23128 480 23158
rect 2773 23155 2839 23158
rect 3558 23216 10426 23218
rect 3558 23160 7654 23216
rect 7710 23160 10426 23216
rect 3558 23158 10426 23160
rect 1945 23082 2011 23085
rect 3558 23082 3618 23158
rect 7649 23155 7715 23158
rect 1945 23080 3618 23082
rect 1945 23024 1950 23080
rect 2006 23024 3618 23080
rect 1945 23022 3618 23024
rect 3693 23082 3759 23085
rect 9213 23082 9279 23085
rect 3693 23080 9279 23082
rect 3693 23024 3698 23080
rect 3754 23024 9218 23080
rect 9274 23024 9279 23080
rect 3693 23022 9279 23024
rect 10366 23082 10426 23158
rect 10593 23216 14339 23218
rect 10593 23160 10598 23216
rect 10654 23160 14278 23216
rect 14334 23160 14339 23216
rect 10593 23158 14339 23160
rect 10593 23155 10659 23158
rect 14273 23155 14339 23158
rect 15929 23218 15995 23221
rect 17953 23218 18019 23221
rect 15929 23216 18019 23218
rect 15929 23160 15934 23216
rect 15990 23160 17958 23216
rect 18014 23160 18019 23216
rect 15929 23158 18019 23160
rect 18094 23218 18154 23294
rect 26509 23218 26575 23221
rect 18094 23216 26575 23218
rect 18094 23160 26514 23216
rect 26570 23160 26575 23216
rect 18094 23158 26575 23160
rect 15929 23155 15995 23158
rect 17953 23155 18019 23158
rect 26509 23155 26575 23158
rect 12065 23082 12131 23085
rect 10366 23080 12131 23082
rect 10366 23024 12070 23080
rect 12126 23024 12131 23080
rect 10366 23022 12131 23024
rect 1945 23019 2011 23022
rect 3693 23019 3759 23022
rect 9213 23019 9279 23022
rect 12065 23019 12131 23022
rect 6637 22946 6703 22949
rect 13629 22946 13695 22949
rect 6637 22944 13695 22946
rect 6637 22888 6642 22944
rect 6698 22888 13634 22944
rect 13690 22888 13695 22944
rect 6637 22886 13695 22888
rect 6637 22883 6703 22886
rect 13629 22883 13695 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 8569 22810 8635 22813
rect 11789 22810 11855 22813
rect 8569 22808 11855 22810
rect 8569 22752 8574 22808
rect 8630 22752 11794 22808
rect 11850 22752 11855 22808
rect 8569 22750 11855 22752
rect 8569 22747 8635 22750
rect 11789 22747 11855 22750
rect 3969 22674 4035 22677
rect 6637 22674 6703 22677
rect 3969 22672 6703 22674
rect 3969 22616 3974 22672
rect 4030 22616 6642 22672
rect 6698 22616 6703 22672
rect 3969 22614 6703 22616
rect 3969 22611 4035 22614
rect 6637 22611 6703 22614
rect 0 22538 480 22568
rect 3877 22538 3943 22541
rect 0 22536 3943 22538
rect 0 22480 3882 22536
rect 3938 22480 3943 22536
rect 0 22478 3943 22480
rect 0 22448 480 22478
rect 3877 22475 3943 22478
rect 4981 22538 5047 22541
rect 10685 22538 10751 22541
rect 4981 22536 10751 22538
rect 4981 22480 4986 22536
rect 5042 22480 10690 22536
rect 10746 22480 10751 22536
rect 4981 22478 10751 22480
rect 4981 22475 5047 22478
rect 10685 22475 10751 22478
rect 13813 22538 13879 22541
rect 21725 22538 21791 22541
rect 13813 22536 21791 22538
rect 13813 22480 13818 22536
rect 13874 22480 21730 22536
rect 21786 22480 21791 22536
rect 13813 22478 21791 22480
rect 13813 22475 13879 22478
rect 21725 22475 21791 22478
rect 14641 22402 14707 22405
rect 16021 22402 16087 22405
rect 14641 22400 16087 22402
rect 14641 22344 14646 22400
rect 14702 22344 16026 22400
rect 16082 22344 16087 22400
rect 14641 22342 16087 22344
rect 14641 22339 14707 22342
rect 16021 22339 16087 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 13721 22266 13787 22269
rect 15837 22266 15903 22269
rect 13721 22264 15903 22266
rect 13721 22208 13726 22264
rect 13782 22208 15842 22264
rect 15898 22208 15903 22264
rect 13721 22206 15903 22208
rect 13721 22203 13787 22206
rect 15837 22203 15903 22206
rect 2865 22130 2931 22133
rect 11513 22130 11579 22133
rect 2865 22128 11579 22130
rect 2865 22072 2870 22128
rect 2926 22072 11518 22128
rect 11574 22072 11579 22128
rect 2865 22070 11579 22072
rect 2865 22067 2931 22070
rect 11513 22067 11579 22070
rect 0 21994 480 22024
rect 2313 21994 2379 21997
rect 0 21992 2379 21994
rect 0 21936 2318 21992
rect 2374 21936 2379 21992
rect 0 21934 2379 21936
rect 0 21904 480 21934
rect 2313 21931 2379 21934
rect 2497 21994 2563 21997
rect 10869 21994 10935 21997
rect 12525 21994 12591 21997
rect 2497 21992 7666 21994
rect 2497 21936 2502 21992
rect 2558 21936 7666 21992
rect 2497 21934 7666 21936
rect 2497 21931 2563 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 7606 21722 7666 21934
rect 10869 21992 12591 21994
rect 10869 21936 10874 21992
rect 10930 21936 12530 21992
rect 12586 21936 12591 21992
rect 10869 21934 12591 21936
rect 10869 21931 10935 21934
rect 12525 21931 12591 21934
rect 17033 21994 17099 21997
rect 24853 21994 24919 21997
rect 17033 21992 24919 21994
rect 17033 21936 17038 21992
rect 17094 21936 24858 21992
rect 24914 21936 24919 21992
rect 17033 21934 24919 21936
rect 17033 21931 17099 21934
rect 24853 21931 24919 21934
rect 9121 21858 9187 21861
rect 12617 21858 12683 21861
rect 9121 21856 12683 21858
rect 9121 21800 9126 21856
rect 9182 21800 12622 21856
rect 12678 21800 12683 21856
rect 9121 21798 12683 21800
rect 9121 21795 9187 21798
rect 12617 21795 12683 21798
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 12341 21722 12407 21725
rect 7606 21720 12407 21722
rect 7606 21664 12346 21720
rect 12402 21664 12407 21720
rect 7606 21662 12407 21664
rect 12341 21659 12407 21662
rect 2497 21450 2563 21453
rect 4245 21450 4311 21453
rect 2497 21448 4311 21450
rect 2497 21392 2502 21448
rect 2558 21392 4250 21448
rect 4306 21392 4311 21448
rect 2497 21390 4311 21392
rect 2497 21387 2563 21390
rect 4245 21387 4311 21390
rect 6821 21450 6887 21453
rect 16757 21450 16823 21453
rect 6821 21448 16823 21450
rect 6821 21392 6826 21448
rect 6882 21392 16762 21448
rect 16818 21392 16823 21448
rect 6821 21390 16823 21392
rect 6821 21387 6887 21390
rect 16757 21387 16823 21390
rect 0 21314 480 21344
rect 3969 21314 4035 21317
rect 0 21312 4035 21314
rect 0 21256 3974 21312
rect 4030 21256 4035 21312
rect 0 21254 4035 21256
rect 0 21224 480 21254
rect 3969 21251 4035 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 3325 21042 3391 21045
rect 13445 21042 13511 21045
rect 14181 21042 14247 21045
rect 15377 21042 15443 21045
rect 3325 21040 15443 21042
rect 3325 20984 3330 21040
rect 3386 20984 13450 21040
rect 13506 20984 14186 21040
rect 14242 20984 15382 21040
rect 15438 20984 15443 21040
rect 3325 20982 15443 20984
rect 3325 20979 3391 20982
rect 13445 20979 13511 20982
rect 14181 20979 14247 20982
rect 15377 20979 15443 20982
rect 24117 21042 24183 21045
rect 27520 21042 28000 21072
rect 24117 21040 28000 21042
rect 24117 20984 24122 21040
rect 24178 20984 28000 21040
rect 24117 20982 28000 20984
rect 24117 20979 24183 20982
rect 27520 20952 28000 20982
rect 12985 20906 13051 20909
rect 19517 20906 19583 20909
rect 12985 20904 19583 20906
rect 12985 20848 12990 20904
rect 13046 20848 19522 20904
rect 19578 20848 19583 20904
rect 12985 20846 19583 20848
rect 12985 20843 13051 20846
rect 19517 20843 19583 20846
rect 8937 20770 9003 20773
rect 11513 20770 11579 20773
rect 8937 20768 11579 20770
rect 8937 20712 8942 20768
rect 8998 20712 11518 20768
rect 11574 20712 11579 20768
rect 8937 20710 11579 20712
rect 8937 20707 9003 20710
rect 11513 20707 11579 20710
rect 5610 20704 5930 20705
rect 0 20634 480 20664
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 7557 20634 7623 20637
rect 14641 20634 14707 20637
rect 0 20574 4906 20634
rect 0 20544 480 20574
rect 4846 20498 4906 20574
rect 7557 20632 14707 20634
rect 7557 20576 7562 20632
rect 7618 20576 14646 20632
rect 14702 20576 14707 20632
rect 7557 20574 14707 20576
rect 7557 20571 7623 20574
rect 14641 20571 14707 20574
rect 11329 20498 11395 20501
rect 4846 20496 11395 20498
rect 4846 20440 11334 20496
rect 11390 20440 11395 20496
rect 4846 20438 11395 20440
rect 11329 20435 11395 20438
rect 12525 20498 12591 20501
rect 18045 20498 18111 20501
rect 12525 20496 18111 20498
rect 12525 20440 12530 20496
rect 12586 20440 18050 20496
rect 18106 20440 18111 20496
rect 12525 20438 18111 20440
rect 12525 20435 12591 20438
rect 18045 20435 18111 20438
rect 4429 20362 4495 20365
rect 10777 20362 10843 20365
rect 4429 20360 10843 20362
rect 4429 20304 4434 20360
rect 4490 20304 10782 20360
rect 10838 20304 10843 20360
rect 4429 20302 10843 20304
rect 4429 20299 4495 20302
rect 10777 20299 10843 20302
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 20030 4906 20090
rect 0 20000 480 20030
rect 4846 19954 4906 20030
rect 13813 19954 13879 19957
rect 17217 19954 17283 19957
rect 4846 19952 17283 19954
rect 4846 19896 13818 19952
rect 13874 19896 17222 19952
rect 17278 19896 17283 19952
rect 4846 19894 17283 19896
rect 13813 19891 13879 19894
rect 17217 19891 17283 19894
rect 3693 19818 3759 19821
rect 10593 19818 10659 19821
rect 11421 19818 11487 19821
rect 15929 19818 15995 19821
rect 17585 19818 17651 19821
rect 3693 19816 17651 19818
rect 3693 19760 3698 19816
rect 3754 19760 10598 19816
rect 10654 19760 11426 19816
rect 11482 19760 15934 19816
rect 15990 19760 17590 19816
rect 17646 19760 17651 19816
rect 3693 19758 17651 19760
rect 3693 19755 3759 19758
rect 10593 19755 10659 19758
rect 11421 19755 11487 19758
rect 15929 19755 15995 19758
rect 17585 19755 17651 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 0 19410 480 19440
rect 2681 19410 2747 19413
rect 0 19408 2747 19410
rect 0 19352 2686 19408
rect 2742 19352 2747 19408
rect 0 19350 2747 19352
rect 0 19320 480 19350
rect 2681 19347 2747 19350
rect 13721 19410 13787 19413
rect 15469 19410 15535 19413
rect 13721 19408 15535 19410
rect 13721 19352 13726 19408
rect 13782 19352 15474 19408
rect 15530 19352 15535 19408
rect 13721 19350 15535 19352
rect 13721 19347 13787 19350
rect 15469 19347 15535 19350
rect 16297 19410 16363 19413
rect 20161 19410 20227 19413
rect 16297 19408 20227 19410
rect 16297 19352 16302 19408
rect 16358 19352 20166 19408
rect 20222 19352 20227 19408
rect 16297 19350 20227 19352
rect 16297 19347 16363 19350
rect 20161 19347 20227 19350
rect 5625 19274 5691 19277
rect 12525 19274 12591 19277
rect 5625 19272 12591 19274
rect 5625 19216 5630 19272
rect 5686 19216 12530 19272
rect 12586 19216 12591 19272
rect 5625 19214 12591 19216
rect 5625 19211 5691 19214
rect 12525 19211 12591 19214
rect 13629 19274 13695 19277
rect 15285 19274 15351 19277
rect 13629 19272 15351 19274
rect 13629 19216 13634 19272
rect 13690 19216 15290 19272
rect 15346 19216 15351 19272
rect 13629 19214 15351 19216
rect 13629 19211 13695 19214
rect 15285 19211 15351 19214
rect 11145 19138 11211 19141
rect 15285 19138 15351 19141
rect 11145 19136 15351 19138
rect 11145 19080 11150 19136
rect 11206 19080 15290 19136
rect 15346 19080 15351 19136
rect 11145 19078 15351 19080
rect 11145 19075 11211 19078
rect 15285 19075 15351 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 11237 18866 11303 18869
rect 15653 18866 15719 18869
rect 11237 18864 15719 18866
rect 11237 18808 11242 18864
rect 11298 18808 15658 18864
rect 15714 18808 15719 18864
rect 11237 18806 15719 18808
rect 11237 18803 11303 18806
rect 15653 18803 15719 18806
rect 0 18730 480 18760
rect 2865 18730 2931 18733
rect 0 18728 2931 18730
rect 0 18672 2870 18728
rect 2926 18672 2931 18728
rect 0 18670 2931 18672
rect 0 18640 480 18670
rect 2865 18667 2931 18670
rect 4061 18730 4127 18733
rect 19149 18730 19215 18733
rect 4061 18728 19215 18730
rect 4061 18672 4066 18728
rect 4122 18672 19154 18728
rect 19210 18672 19215 18728
rect 4061 18670 19215 18672
rect 4061 18667 4127 18670
rect 19149 18667 19215 18670
rect 9213 18594 9279 18597
rect 14733 18594 14799 18597
rect 9213 18592 14799 18594
rect 9213 18536 9218 18592
rect 9274 18536 14738 18592
rect 14794 18536 14799 18592
rect 9213 18534 14799 18536
rect 9213 18531 9279 18534
rect 14733 18531 14799 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 9305 18458 9371 18461
rect 9305 18456 14842 18458
rect 9305 18400 9310 18456
rect 9366 18400 14842 18456
rect 9305 18398 14842 18400
rect 9305 18395 9371 18398
rect 2589 18322 2655 18325
rect 6177 18322 6243 18325
rect 2589 18320 6243 18322
rect 2589 18264 2594 18320
rect 2650 18264 6182 18320
rect 6238 18264 6243 18320
rect 2589 18262 6243 18264
rect 2589 18259 2655 18262
rect 6177 18259 6243 18262
rect 6361 18322 6427 18325
rect 11881 18322 11947 18325
rect 13077 18322 13143 18325
rect 6361 18320 13143 18322
rect 6361 18264 6366 18320
rect 6422 18264 11886 18320
rect 11942 18264 13082 18320
rect 13138 18264 13143 18320
rect 6361 18262 13143 18264
rect 14782 18322 14842 18398
rect 16113 18322 16179 18325
rect 14782 18320 16179 18322
rect 14782 18264 16118 18320
rect 16174 18264 16179 18320
rect 14782 18262 16179 18264
rect 6361 18259 6427 18262
rect 11881 18259 11947 18262
rect 13077 18259 13143 18262
rect 16113 18259 16179 18262
rect 0 18186 480 18216
rect 4061 18186 4127 18189
rect 0 18184 4127 18186
rect 0 18128 4066 18184
rect 4122 18128 4127 18184
rect 0 18126 4127 18128
rect 0 18096 480 18126
rect 4061 18123 4127 18126
rect 9765 18186 9831 18189
rect 15377 18186 15443 18189
rect 9765 18184 15443 18186
rect 9765 18128 9770 18184
rect 9826 18128 15382 18184
rect 15438 18128 15443 18184
rect 9765 18126 15443 18128
rect 9765 18123 9831 18126
rect 15377 18123 15443 18126
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 3969 17914 4035 17917
rect 8753 17914 8819 17917
rect 9397 17914 9463 17917
rect 3969 17912 9463 17914
rect 3969 17856 3974 17912
rect 4030 17856 8758 17912
rect 8814 17856 9402 17912
rect 9458 17856 9463 17912
rect 3969 17854 9463 17856
rect 3969 17851 4035 17854
rect 8753 17851 8819 17854
rect 9397 17851 9463 17854
rect 10869 17914 10935 17917
rect 13169 17914 13235 17917
rect 10869 17912 13235 17914
rect 10869 17856 10874 17912
rect 10930 17856 13174 17912
rect 13230 17856 13235 17912
rect 10869 17854 13235 17856
rect 10869 17851 10935 17854
rect 13169 17851 13235 17854
rect 15837 17914 15903 17917
rect 18505 17914 18571 17917
rect 15837 17912 18571 17914
rect 15837 17856 15842 17912
rect 15898 17856 18510 17912
rect 18566 17856 18571 17912
rect 15837 17854 18571 17856
rect 15837 17851 15903 17854
rect 18505 17851 18571 17854
rect 7649 17642 7715 17645
rect 21265 17642 21331 17645
rect 7649 17640 21331 17642
rect 7649 17584 7654 17640
rect 7710 17584 21270 17640
rect 21326 17584 21331 17640
rect 7649 17582 21331 17584
rect 7649 17579 7715 17582
rect 21265 17579 21331 17582
rect 0 17506 480 17536
rect 1853 17506 1919 17509
rect 0 17504 1919 17506
rect 0 17448 1858 17504
rect 1914 17448 1919 17504
rect 0 17446 1919 17448
rect 0 17416 480 17446
rect 1853 17443 1919 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 7925 17370 7991 17373
rect 9949 17370 10015 17373
rect 7925 17368 10015 17370
rect 7925 17312 7930 17368
rect 7986 17312 9954 17368
rect 10010 17312 10015 17368
rect 7925 17310 10015 17312
rect 7925 17307 7991 17310
rect 9949 17307 10015 17310
rect 9489 17098 9555 17101
rect 15837 17098 15903 17101
rect 9489 17096 15903 17098
rect 9489 17040 9494 17096
rect 9550 17040 15842 17096
rect 15898 17040 15903 17096
rect 9489 17038 15903 17040
rect 9489 17035 9555 17038
rect 15837 17035 15903 17038
rect 9673 16962 9739 16965
rect 10041 16962 10107 16965
rect 1350 16960 10107 16962
rect 1350 16904 9678 16960
rect 9734 16904 10046 16960
rect 10102 16904 10107 16960
rect 1350 16902 10107 16904
rect 0 16826 480 16856
rect 1350 16826 1410 16902
rect 9673 16899 9739 16902
rect 10041 16899 10107 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 0 16766 1410 16826
rect 6269 16826 6335 16829
rect 8017 16826 8083 16829
rect 6269 16824 8083 16826
rect 6269 16768 6274 16824
rect 6330 16768 8022 16824
rect 8078 16768 8083 16824
rect 6269 16766 8083 16768
rect 0 16736 480 16766
rect 6269 16763 6335 16766
rect 8017 16763 8083 16766
rect 10133 16690 10199 16693
rect 4800 16688 10199 16690
rect 4800 16632 10138 16688
rect 10194 16632 10199 16688
rect 4800 16630 10199 16632
rect 0 16282 480 16312
rect 4800 16282 4860 16630
rect 10133 16627 10199 16630
rect 12801 16690 12867 16693
rect 16665 16690 16731 16693
rect 12801 16688 16731 16690
rect 12801 16632 12806 16688
rect 12862 16632 16670 16688
rect 16726 16632 16731 16688
rect 12801 16630 16731 16632
rect 12801 16627 12867 16630
rect 16665 16627 16731 16630
rect 14181 16554 14247 16557
rect 15285 16554 15351 16557
rect 14181 16552 15351 16554
rect 14181 16496 14186 16552
rect 14242 16496 15290 16552
rect 15346 16496 15351 16552
rect 14181 16494 15351 16496
rect 14181 16491 14247 16494
rect 15285 16491 15351 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 16222 4860 16282
rect 5993 16282 6059 16285
rect 11605 16282 11671 16285
rect 5993 16280 11671 16282
rect 5993 16224 5998 16280
rect 6054 16224 11610 16280
rect 11666 16224 11671 16280
rect 5993 16222 11671 16224
rect 0 16192 480 16222
rect 5993 16219 6059 16222
rect 11605 16219 11671 16222
rect 5257 16146 5323 16149
rect 13353 16146 13419 16149
rect 16297 16146 16363 16149
rect 5257 16144 13419 16146
rect 5257 16088 5262 16144
rect 5318 16088 13358 16144
rect 13414 16088 13419 16144
rect 5257 16086 13419 16088
rect 5257 16083 5323 16086
rect 13353 16083 13419 16086
rect 13862 16144 16363 16146
rect 13862 16088 16302 16144
rect 16358 16088 16363 16144
rect 13862 16086 16363 16088
rect 7373 16010 7439 16013
rect 11973 16010 12039 16013
rect 13862 16010 13922 16086
rect 16297 16083 16363 16086
rect 7373 16008 13922 16010
rect 7373 15952 7378 16008
rect 7434 15952 11978 16008
rect 12034 15952 13922 16008
rect 7373 15950 13922 15952
rect 14089 16010 14155 16013
rect 24117 16010 24183 16013
rect 14089 16008 24183 16010
rect 14089 15952 14094 16008
rect 14150 15952 24122 16008
rect 24178 15952 24183 16008
rect 14089 15950 24183 15952
rect 7373 15947 7439 15950
rect 11973 15947 12039 15950
rect 14089 15947 14155 15950
rect 24117 15947 24183 15950
rect 3969 15874 4035 15877
rect 6177 15874 6243 15877
rect 3969 15872 6243 15874
rect 3969 15816 3974 15872
rect 4030 15816 6182 15872
rect 6238 15816 6243 15872
rect 3969 15814 6243 15816
rect 3969 15811 4035 15814
rect 6177 15811 6243 15814
rect 11605 15874 11671 15877
rect 16297 15874 16363 15877
rect 11605 15872 16363 15874
rect 11605 15816 11610 15872
rect 11666 15816 16302 15872
rect 16358 15816 16363 15872
rect 11605 15814 16363 15816
rect 11605 15811 11671 15814
rect 16297 15811 16363 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 11513 15738 11579 15741
rect 13813 15738 13879 15741
rect 14273 15738 14339 15741
rect 11513 15736 13879 15738
rect 11513 15680 11518 15736
rect 11574 15680 13818 15736
rect 13874 15680 13879 15736
rect 11513 15678 13879 15680
rect 11513 15675 11579 15678
rect 13813 15675 13879 15678
rect 14230 15736 14339 15738
rect 14230 15680 14278 15736
rect 14334 15680 14339 15736
rect 14230 15675 14339 15680
rect 0 15602 480 15632
rect 4429 15602 4495 15605
rect 8293 15602 8359 15605
rect 0 15542 1410 15602
rect 0 15512 480 15542
rect 1350 15466 1410 15542
rect 4429 15600 8359 15602
rect 4429 15544 4434 15600
rect 4490 15544 8298 15600
rect 8354 15544 8359 15600
rect 4429 15542 8359 15544
rect 4429 15539 4495 15542
rect 8293 15539 8359 15542
rect 14230 15466 14290 15675
rect 17401 15466 17467 15469
rect 1350 15464 17467 15466
rect 1350 15408 17406 15464
rect 17462 15408 17467 15464
rect 1350 15406 17467 15408
rect 17401 15403 17467 15406
rect 2037 15330 2103 15333
rect 4889 15330 4955 15333
rect 2037 15328 4955 15330
rect 2037 15272 2042 15328
rect 2098 15272 4894 15328
rect 4950 15272 4955 15328
rect 2037 15270 4955 15272
rect 2037 15267 2103 15270
rect 4889 15267 4955 15270
rect 8753 15330 8819 15333
rect 11145 15330 11211 15333
rect 13445 15330 13511 15333
rect 8753 15328 13511 15330
rect 8753 15272 8758 15328
rect 8814 15272 11150 15328
rect 11206 15272 13450 15328
rect 13506 15272 13511 15328
rect 8753 15270 13511 15272
rect 8753 15267 8819 15270
rect 11145 15267 11211 15270
rect 13445 15267 13511 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 18045 15194 18111 15197
rect 21817 15194 21883 15197
rect 18045 15192 21883 15194
rect 18045 15136 18050 15192
rect 18106 15136 21822 15192
rect 21878 15136 21883 15192
rect 18045 15134 21883 15136
rect 18045 15131 18111 15134
rect 21817 15131 21883 15134
rect 0 14922 480 14952
rect 9213 14922 9279 14925
rect 0 14920 9279 14922
rect 0 14864 9218 14920
rect 9274 14864 9279 14920
rect 0 14862 9279 14864
rect 0 14832 480 14862
rect 9213 14859 9279 14862
rect 14549 14786 14615 14789
rect 17493 14786 17559 14789
rect 14549 14784 17559 14786
rect 14549 14728 14554 14784
rect 14610 14728 17498 14784
rect 17554 14728 17559 14784
rect 14549 14726 17559 14728
rect 14549 14723 14615 14726
rect 17493 14723 17559 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 0 14378 480 14408
rect 2037 14378 2103 14381
rect 0 14376 2103 14378
rect 0 14320 2042 14376
rect 2098 14320 2103 14376
rect 0 14318 2103 14320
rect 0 14288 480 14318
rect 2037 14315 2103 14318
rect 10777 14242 10843 14245
rect 12893 14242 12959 14245
rect 10777 14240 12959 14242
rect 10777 14184 10782 14240
rect 10838 14184 12898 14240
rect 12954 14184 12959 14240
rect 10777 14182 12959 14184
rect 10777 14179 10843 14182
rect 12893 14179 12959 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 6453 13970 6519 13973
rect 10133 13970 10199 13973
rect 6453 13968 10199 13970
rect 6453 13912 6458 13968
rect 6514 13912 10138 13968
rect 10194 13912 10199 13968
rect 6453 13910 10199 13912
rect 6453 13907 6519 13910
rect 10133 13907 10199 13910
rect 10869 13970 10935 13973
rect 18505 13970 18571 13973
rect 10869 13968 18571 13970
rect 10869 13912 10874 13968
rect 10930 13912 18510 13968
rect 18566 13912 18571 13968
rect 10869 13910 18571 13912
rect 10869 13907 10935 13910
rect 18505 13907 18571 13910
rect 2221 13834 2287 13837
rect 6729 13834 6795 13837
rect 2221 13832 6795 13834
rect 2221 13776 2226 13832
rect 2282 13776 6734 13832
rect 6790 13776 6795 13832
rect 2221 13774 6795 13776
rect 2221 13771 2287 13774
rect 6729 13771 6795 13774
rect 9397 13834 9463 13837
rect 12617 13834 12683 13837
rect 9397 13832 12683 13834
rect 9397 13776 9402 13832
rect 9458 13776 12622 13832
rect 12678 13776 12683 13832
rect 9397 13774 12683 13776
rect 9397 13771 9463 13774
rect 12617 13771 12683 13774
rect 0 13698 480 13728
rect 2129 13698 2195 13701
rect 9581 13698 9647 13701
rect 10133 13698 10199 13701
rect 0 13638 1410 13698
rect 0 13608 480 13638
rect 1350 13426 1410 13638
rect 2129 13696 7666 13698
rect 2129 13640 2134 13696
rect 2190 13640 7666 13696
rect 2129 13638 7666 13640
rect 2129 13635 2195 13638
rect 1669 13562 1735 13565
rect 7465 13562 7531 13565
rect 1669 13560 7531 13562
rect 1669 13504 1674 13560
rect 1730 13504 7470 13560
rect 7526 13504 7531 13560
rect 1669 13502 7531 13504
rect 1669 13499 1735 13502
rect 7465 13499 7531 13502
rect 3969 13426 4035 13429
rect 1350 13424 4035 13426
rect 1350 13368 3974 13424
rect 4030 13368 4035 13424
rect 1350 13366 4035 13368
rect 7606 13426 7666 13638
rect 9581 13696 10199 13698
rect 9581 13640 9586 13696
rect 9642 13640 10138 13696
rect 10194 13640 10199 13696
rect 9581 13638 10199 13640
rect 9581 13635 9647 13638
rect 10133 13635 10199 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 12801 13426 12867 13429
rect 7606 13424 12867 13426
rect 7606 13368 12806 13424
rect 12862 13368 12867 13424
rect 7606 13366 12867 13368
rect 3969 13363 4035 13366
rect 12801 13363 12867 13366
rect 14917 13426 14983 13429
rect 16573 13426 16639 13429
rect 14917 13424 16639 13426
rect 14917 13368 14922 13424
rect 14978 13368 16578 13424
rect 16634 13368 16639 13424
rect 14917 13366 16639 13368
rect 14917 13363 14983 13366
rect 16573 13363 16639 13366
rect 4153 13290 4219 13293
rect 14181 13290 14247 13293
rect 4153 13288 14247 13290
rect 4153 13232 4158 13288
rect 4214 13232 14186 13288
rect 14242 13232 14247 13288
rect 4153 13230 14247 13232
rect 4153 13227 4219 13230
rect 14181 13227 14247 13230
rect 15745 13290 15811 13293
rect 26233 13290 26299 13293
rect 15745 13288 26299 13290
rect 15745 13232 15750 13288
rect 15806 13232 26238 13288
rect 26294 13232 26299 13288
rect 15745 13230 26299 13232
rect 15745 13227 15811 13230
rect 26233 13227 26299 13230
rect 11789 13154 11855 13157
rect 12893 13154 12959 13157
rect 11789 13152 12959 13154
rect 11789 13096 11794 13152
rect 11850 13096 12898 13152
rect 12954 13096 12959 13152
rect 11789 13094 12959 13096
rect 11789 13091 11855 13094
rect 12893 13091 12959 13094
rect 16297 13154 16363 13157
rect 20161 13154 20227 13157
rect 16297 13152 20227 13154
rect 16297 13096 16302 13152
rect 16358 13096 20166 13152
rect 20222 13096 20227 13152
rect 16297 13094 20227 13096
rect 16297 13091 16363 13094
rect 20161 13091 20227 13094
rect 5610 13088 5930 13089
rect 0 13018 480 13048
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 1761 13018 1827 13021
rect 1945 13018 2011 13021
rect 0 13016 2011 13018
rect 0 12960 1766 13016
rect 1822 12960 1950 13016
rect 2006 12960 2011 13016
rect 0 12958 2011 12960
rect 0 12928 480 12958
rect 1761 12955 1827 12958
rect 1945 12955 2011 12958
rect 7373 13018 7439 13021
rect 11605 13018 11671 13021
rect 7373 13016 11671 13018
rect 7373 12960 7378 13016
rect 7434 12960 11610 13016
rect 11666 12960 11671 13016
rect 7373 12958 11671 12960
rect 7373 12955 7439 12958
rect 11605 12955 11671 12958
rect 2865 12882 2931 12885
rect 11789 12882 11855 12885
rect 2865 12880 11855 12882
rect 2865 12824 2870 12880
rect 2926 12824 11794 12880
rect 11850 12824 11855 12880
rect 2865 12822 11855 12824
rect 2865 12819 2931 12822
rect 11789 12819 11855 12822
rect 1761 12746 1827 12749
rect 16021 12746 16087 12749
rect 1761 12744 16087 12746
rect 1761 12688 1766 12744
rect 1822 12688 16026 12744
rect 16082 12688 16087 12744
rect 1761 12686 16087 12688
rect 1761 12683 1827 12686
rect 16021 12683 16087 12686
rect 6545 12612 6611 12613
rect 6494 12610 6500 12612
rect 6454 12550 6500 12610
rect 6564 12608 6611 12612
rect 6606 12552 6611 12608
rect 6494 12548 6500 12550
rect 6564 12548 6611 12552
rect 6545 12547 6611 12548
rect 11605 12610 11671 12613
rect 11881 12610 11947 12613
rect 11605 12608 11947 12610
rect 11605 12552 11610 12608
rect 11666 12552 11886 12608
rect 11942 12552 11947 12608
rect 11605 12550 11947 12552
rect 11605 12547 11671 12550
rect 11881 12547 11947 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 5533 12474 5599 12477
rect 3006 12472 5599 12474
rect 3006 12416 5538 12472
rect 5594 12416 5599 12472
rect 3006 12414 5599 12416
rect 0 12338 480 12368
rect 3006 12338 3066 12414
rect 5533 12411 5599 12414
rect 12249 12474 12315 12477
rect 15377 12474 15443 12477
rect 12249 12472 15443 12474
rect 12249 12416 12254 12472
rect 12310 12416 15382 12472
rect 15438 12416 15443 12472
rect 12249 12414 15443 12416
rect 12249 12411 12315 12414
rect 15377 12411 15443 12414
rect 0 12278 3066 12338
rect 4429 12338 4495 12341
rect 10685 12338 10751 12341
rect 4429 12336 10751 12338
rect 4429 12280 4434 12336
rect 4490 12280 10690 12336
rect 10746 12280 10751 12336
rect 4429 12278 10751 12280
rect 0 12248 480 12278
rect 4429 12275 4495 12278
rect 10685 12275 10751 12278
rect 11881 12338 11947 12341
rect 12709 12338 12775 12341
rect 11881 12336 12775 12338
rect 11881 12280 11886 12336
rect 11942 12280 12714 12336
rect 12770 12280 12775 12336
rect 11881 12278 12775 12280
rect 11881 12275 11947 12278
rect 12709 12275 12775 12278
rect 12985 12338 13051 12341
rect 15837 12338 15903 12341
rect 25957 12338 26023 12341
rect 12985 12336 26023 12338
rect 12985 12280 12990 12336
rect 13046 12280 15842 12336
rect 15898 12280 25962 12336
rect 26018 12280 26023 12336
rect 12985 12278 26023 12280
rect 12985 12275 13051 12278
rect 15837 12275 15903 12278
rect 25957 12275 26023 12278
rect 3969 12202 4035 12205
rect 9029 12202 9095 12205
rect 3969 12200 9095 12202
rect 3969 12144 3974 12200
rect 4030 12144 9034 12200
rect 9090 12144 9095 12200
rect 3969 12142 9095 12144
rect 3969 12139 4035 12142
rect 9029 12139 9095 12142
rect 9305 12202 9371 12205
rect 13169 12202 13235 12205
rect 9305 12200 13235 12202
rect 9305 12144 9310 12200
rect 9366 12144 13174 12200
rect 13230 12144 13235 12200
rect 9305 12142 13235 12144
rect 9305 12139 9371 12142
rect 13169 12139 13235 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 0 11794 480 11824
rect 2681 11794 2747 11797
rect 0 11792 2747 11794
rect 0 11736 2686 11792
rect 2742 11736 2747 11792
rect 0 11734 2747 11736
rect 0 11704 480 11734
rect 2681 11731 2747 11734
rect 4797 11794 4863 11797
rect 7373 11794 7439 11797
rect 4797 11792 7439 11794
rect 4797 11736 4802 11792
rect 4858 11736 7378 11792
rect 7434 11736 7439 11792
rect 4797 11734 7439 11736
rect 4797 11731 4863 11734
rect 7373 11731 7439 11734
rect 12709 11794 12775 11797
rect 17125 11794 17191 11797
rect 12709 11792 17191 11794
rect 12709 11736 12714 11792
rect 12770 11736 17130 11792
rect 17186 11736 17191 11792
rect 12709 11734 17191 11736
rect 12709 11731 12775 11734
rect 17125 11731 17191 11734
rect 3141 11658 3207 11661
rect 4797 11658 4863 11661
rect 11513 11658 11579 11661
rect 3141 11656 11579 11658
rect 3141 11600 3146 11656
rect 3202 11600 4802 11656
rect 4858 11600 11518 11656
rect 11574 11600 11579 11656
rect 3141 11598 11579 11600
rect 3141 11595 3207 11598
rect 4797 11595 4863 11598
rect 11513 11595 11579 11598
rect 2681 11522 2747 11525
rect 4337 11522 4403 11525
rect 2681 11520 4403 11522
rect 2681 11464 2686 11520
rect 2742 11464 4342 11520
rect 4398 11464 4403 11520
rect 2681 11462 4403 11464
rect 2681 11459 2747 11462
rect 4337 11459 4403 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 6453 11386 6519 11389
rect 9949 11386 10015 11389
rect 3742 11384 10015 11386
rect 3742 11328 6458 11384
rect 6514 11328 9954 11384
rect 10010 11328 10015 11384
rect 3742 11326 10015 11328
rect 565 11250 631 11253
rect 3742 11250 3802 11326
rect 6453 11323 6519 11326
rect 9949 11323 10015 11326
rect 565 11248 3802 11250
rect 565 11192 570 11248
rect 626 11192 3802 11248
rect 565 11190 3802 11192
rect 565 11187 631 11190
rect 0 11114 480 11144
rect 6085 11114 6151 11117
rect 0 11112 6151 11114
rect 0 11056 6090 11112
rect 6146 11056 6151 11112
rect 0 11054 6151 11056
rect 0 11024 480 11054
rect 6085 11051 6151 11054
rect 9765 11114 9831 11117
rect 12709 11114 12775 11117
rect 9765 11112 12775 11114
rect 9765 11056 9770 11112
rect 9826 11056 12714 11112
rect 12770 11056 12775 11112
rect 9765 11054 12775 11056
rect 9765 11051 9831 11054
rect 12709 11051 12775 11054
rect 13261 11114 13327 11117
rect 15929 11114 15995 11117
rect 13261 11112 15995 11114
rect 13261 11056 13266 11112
rect 13322 11056 15934 11112
rect 15990 11056 15995 11112
rect 13261 11054 15995 11056
rect 13261 11051 13327 11054
rect 15929 11051 15995 11054
rect 5993 10978 6059 10981
rect 9857 10978 9923 10981
rect 11513 10978 11579 10981
rect 5993 10976 11579 10978
rect 5993 10920 5998 10976
rect 6054 10920 9862 10976
rect 9918 10920 11518 10976
rect 11574 10920 11579 10976
rect 5993 10918 11579 10920
rect 5993 10915 6059 10918
rect 9857 10915 9923 10918
rect 11513 10915 11579 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 7465 10842 7531 10845
rect 7741 10842 7807 10845
rect 7465 10840 7807 10842
rect 7465 10784 7470 10840
rect 7526 10784 7746 10840
rect 7802 10784 7807 10840
rect 7465 10782 7807 10784
rect 7465 10779 7531 10782
rect 7741 10779 7807 10782
rect 8569 10842 8635 10845
rect 12525 10842 12591 10845
rect 21357 10842 21423 10845
rect 8569 10840 12591 10842
rect 8569 10784 8574 10840
rect 8630 10784 12530 10840
rect 12586 10784 12591 10840
rect 8569 10782 12591 10784
rect 8569 10779 8635 10782
rect 12525 10779 12591 10782
rect 19382 10840 21423 10842
rect 19382 10784 21362 10840
rect 21418 10784 21423 10840
rect 19382 10782 21423 10784
rect 3969 10706 4035 10709
rect 12893 10706 12959 10709
rect 3969 10704 12959 10706
rect 3969 10648 3974 10704
rect 4030 10648 12898 10704
rect 12954 10648 12959 10704
rect 3969 10646 12959 10648
rect 3969 10643 4035 10646
rect 12893 10643 12959 10646
rect 5625 10570 5691 10573
rect 19382 10570 19442 10782
rect 21357 10779 21423 10782
rect 5625 10568 19442 10570
rect 5625 10512 5630 10568
rect 5686 10512 19442 10568
rect 5625 10510 19442 10512
rect 5625 10507 5691 10510
rect 0 10434 480 10464
rect 1577 10434 1643 10437
rect 0 10432 1643 10434
rect 0 10376 1582 10432
rect 1638 10376 1643 10432
rect 0 10374 1643 10376
rect 0 10344 480 10374
rect 1577 10371 1643 10374
rect 5533 10434 5599 10437
rect 8017 10434 8083 10437
rect 5533 10432 8083 10434
rect 5533 10376 5538 10432
rect 5594 10376 8022 10432
rect 8078 10376 8083 10432
rect 5533 10374 8083 10376
rect 5533 10371 5599 10374
rect 8017 10371 8083 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 3785 10298 3851 10301
rect 5717 10298 5783 10301
rect 3785 10296 5783 10298
rect 3785 10240 3790 10296
rect 3846 10240 5722 10296
rect 5778 10240 5783 10296
rect 3785 10238 5783 10240
rect 3785 10235 3851 10238
rect 5717 10235 5783 10238
rect 9029 10162 9095 10165
rect 15377 10162 15443 10165
rect 9029 10160 15443 10162
rect 9029 10104 9034 10160
rect 9090 10104 15382 10160
rect 15438 10104 15443 10160
rect 9029 10102 15443 10104
rect 9029 10099 9095 10102
rect 15377 10099 15443 10102
rect 4061 10026 4127 10029
rect 9857 10026 9923 10029
rect 4061 10024 9923 10026
rect 4061 9968 4066 10024
rect 4122 9968 9862 10024
rect 9918 9968 9923 10024
rect 4061 9966 9923 9968
rect 4061 9963 4127 9966
rect 9857 9963 9923 9966
rect 0 9890 480 9920
rect 4889 9890 4955 9893
rect 0 9888 4955 9890
rect 0 9832 4894 9888
rect 4950 9832 4955 9888
rect 0 9830 4955 9832
rect 0 9800 480 9830
rect 4889 9827 4955 9830
rect 6637 9890 6703 9893
rect 9213 9890 9279 9893
rect 6637 9888 9279 9890
rect 6637 9832 6642 9888
rect 6698 9832 9218 9888
rect 9274 9832 9279 9888
rect 6637 9830 9279 9832
rect 6637 9827 6703 9830
rect 9213 9827 9279 9830
rect 11789 9890 11855 9893
rect 12341 9890 12407 9893
rect 11789 9888 12407 9890
rect 11789 9832 11794 9888
rect 11850 9832 12346 9888
rect 12402 9832 12407 9888
rect 11789 9830 12407 9832
rect 11789 9827 11855 9830
rect 12341 9827 12407 9830
rect 15561 9890 15627 9893
rect 22001 9890 22067 9893
rect 15561 9888 22067 9890
rect 15561 9832 15566 9888
rect 15622 9832 22006 9888
rect 22062 9832 22067 9888
rect 15561 9830 22067 9832
rect 15561 9827 15627 9830
rect 22001 9827 22067 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 7649 9754 7715 9757
rect 14181 9754 14247 9757
rect 7649 9752 14247 9754
rect 7649 9696 7654 9752
rect 7710 9696 14186 9752
rect 14242 9696 14247 9752
rect 7649 9694 14247 9696
rect 7649 9691 7715 9694
rect 14181 9691 14247 9694
rect 14457 9652 14523 9655
rect 14457 9650 14658 9652
rect 8385 9618 8451 9621
rect 11881 9618 11947 9621
rect 12341 9618 12407 9621
rect 8385 9616 12407 9618
rect 8385 9560 8390 9616
rect 8446 9560 11886 9616
rect 11942 9560 12346 9616
rect 12402 9560 12407 9616
rect 8385 9558 12407 9560
rect 8385 9555 8451 9558
rect 11881 9555 11947 9558
rect 12341 9555 12407 9558
rect 13077 9618 13143 9621
rect 13445 9618 13511 9621
rect 13077 9616 13511 9618
rect 13077 9560 13082 9616
rect 13138 9560 13450 9616
rect 13506 9560 13511 9616
rect 14457 9594 14462 9650
rect 14518 9618 14658 9650
rect 14825 9618 14891 9621
rect 14518 9616 14891 9618
rect 14518 9594 14830 9616
rect 14457 9592 14830 9594
rect 14457 9589 14523 9592
rect 13077 9558 13511 9560
rect 14598 9560 14830 9592
rect 14886 9560 14891 9616
rect 14598 9558 14891 9560
rect 13077 9555 13143 9558
rect 13445 9555 13511 9558
rect 14825 9555 14891 9558
rect 1853 9482 1919 9485
rect 9673 9482 9739 9485
rect 16113 9482 16179 9485
rect 20897 9482 20963 9485
rect 1853 9480 9739 9482
rect 1853 9424 1858 9480
rect 1914 9424 9678 9480
rect 9734 9424 9739 9480
rect 1853 9422 9739 9424
rect 1853 9419 1919 9422
rect 9673 9419 9739 9422
rect 9814 9480 20963 9482
rect 9814 9424 16118 9480
rect 16174 9424 20902 9480
rect 20958 9424 20963 9480
rect 9814 9422 20963 9424
rect 7189 9346 7255 9349
rect 7649 9346 7715 9349
rect 9814 9346 9874 9422
rect 16113 9419 16179 9422
rect 20897 9419 20963 9422
rect 7189 9344 9874 9346
rect 7189 9288 7194 9344
rect 7250 9288 7654 9344
rect 7710 9288 9874 9344
rect 7189 9286 9874 9288
rect 7189 9283 7255 9286
rect 7649 9283 7715 9286
rect 10277 9280 10597 9281
rect 0 9210 480 9240
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 3969 9210 4035 9213
rect 0 9208 4035 9210
rect 0 9152 3974 9208
rect 4030 9152 4035 9208
rect 0 9150 4035 9152
rect 0 9120 480 9150
rect 3969 9147 4035 9150
rect 4981 9210 5047 9213
rect 6126 9210 6132 9212
rect 4981 9208 6132 9210
rect 4981 9152 4986 9208
rect 5042 9152 6132 9208
rect 4981 9150 6132 9152
rect 4981 9147 5047 9150
rect 6126 9148 6132 9150
rect 6196 9148 6202 9212
rect 13997 9210 14063 9213
rect 16389 9210 16455 9213
rect 13997 9208 16455 9210
rect 13997 9152 14002 9208
rect 14058 9152 16394 9208
rect 16450 9152 16455 9208
rect 13997 9150 16455 9152
rect 13997 9147 14063 9150
rect 16389 9147 16455 9150
rect 3509 9074 3575 9077
rect 11145 9074 11211 9077
rect 3509 9072 11211 9074
rect 3509 9016 3514 9072
rect 3570 9016 11150 9072
rect 11206 9016 11211 9072
rect 3509 9014 11211 9016
rect 3509 9011 3575 9014
rect 11145 9011 11211 9014
rect 2957 8938 3023 8941
rect 12341 8938 12407 8941
rect 2957 8936 12407 8938
rect 2957 8880 2962 8936
rect 3018 8880 12346 8936
rect 12402 8880 12407 8936
rect 2957 8878 12407 8880
rect 2957 8875 3023 8878
rect 12341 8875 12407 8878
rect 13077 8938 13143 8941
rect 15193 8938 15259 8941
rect 13077 8936 15259 8938
rect 13077 8880 13082 8936
rect 13138 8880 15198 8936
rect 15254 8880 15259 8936
rect 13077 8878 15259 8880
rect 13077 8875 13143 8878
rect 15193 8875 15259 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 1853 8666 1919 8669
rect 4981 8666 5047 8669
rect 1853 8664 5047 8666
rect 1853 8608 1858 8664
rect 1914 8608 4986 8664
rect 5042 8608 5047 8664
rect 1853 8606 5047 8608
rect 1853 8603 1919 8606
rect 4981 8603 5047 8606
rect 7281 8666 7347 8669
rect 7281 8664 14842 8666
rect 7281 8608 7286 8664
rect 7342 8608 14842 8664
rect 7281 8606 14842 8608
rect 7281 8603 7347 8606
rect 0 8530 480 8560
rect 1485 8530 1551 8533
rect 0 8528 1551 8530
rect 0 8472 1490 8528
rect 1546 8472 1551 8528
rect 0 8470 1551 8472
rect 0 8440 480 8470
rect 1485 8467 1551 8470
rect 3693 8530 3759 8533
rect 9305 8530 9371 8533
rect 3693 8528 9371 8530
rect 3693 8472 3698 8528
rect 3754 8472 9310 8528
rect 9366 8472 9371 8528
rect 3693 8470 9371 8472
rect 3693 8467 3759 8470
rect 9305 8467 9371 8470
rect 9489 8530 9555 8533
rect 14782 8530 14842 8606
rect 15377 8530 15443 8533
rect 9489 8528 13186 8530
rect 9489 8472 9494 8528
rect 9550 8472 13186 8528
rect 9489 8470 13186 8472
rect 14782 8528 15443 8530
rect 14782 8472 15382 8528
rect 15438 8472 15443 8528
rect 14782 8470 15443 8472
rect 9489 8467 9555 8470
rect 3182 8332 3188 8396
rect 3252 8394 3258 8396
rect 3417 8394 3483 8397
rect 3252 8392 3483 8394
rect 3252 8336 3422 8392
rect 3478 8336 3483 8392
rect 3252 8334 3483 8336
rect 3252 8332 3258 8334
rect 3417 8331 3483 8334
rect 5349 8394 5415 8397
rect 9765 8394 9831 8397
rect 5349 8392 9831 8394
rect 5349 8336 5354 8392
rect 5410 8336 9770 8392
rect 9826 8336 9831 8392
rect 5349 8334 9831 8336
rect 5349 8331 5415 8334
rect 9765 8331 9831 8334
rect 10317 8394 10383 8397
rect 12985 8394 13051 8397
rect 10317 8392 13051 8394
rect 10317 8336 10322 8392
rect 10378 8336 12990 8392
rect 13046 8336 13051 8392
rect 10317 8334 13051 8336
rect 13126 8394 13186 8470
rect 15377 8467 15443 8470
rect 15745 8394 15811 8397
rect 13126 8392 15811 8394
rect 13126 8336 15750 8392
rect 15806 8336 15811 8392
rect 13126 8334 15811 8336
rect 10317 8331 10383 8334
rect 12985 8331 13051 8334
rect 15745 8331 15811 8334
rect 7557 8258 7623 8261
rect 10133 8258 10199 8261
rect 7557 8256 10199 8258
rect 7557 8200 7562 8256
rect 7618 8200 10138 8256
rect 10194 8200 10199 8256
rect 7557 8198 10199 8200
rect 7557 8195 7623 8198
rect 10133 8195 10199 8198
rect 11605 8258 11671 8261
rect 11605 8256 17786 8258
rect 11605 8200 11610 8256
rect 11666 8200 17786 8256
rect 11605 8198 17786 8200
rect 11605 8195 11671 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 7005 8122 7071 8125
rect 7281 8122 7347 8125
rect 7005 8120 7347 8122
rect 7005 8064 7010 8120
rect 7066 8064 7286 8120
rect 7342 8064 7347 8120
rect 7005 8062 7347 8064
rect 7005 8059 7071 8062
rect 7281 8059 7347 8062
rect 0 7986 480 8016
rect 4061 7986 4127 7989
rect 17585 7986 17651 7989
rect 0 7984 4127 7986
rect 0 7928 4066 7984
rect 4122 7928 4127 7984
rect 0 7926 4127 7928
rect 0 7896 480 7926
rect 4061 7923 4127 7926
rect 4294 7984 17651 7986
rect 4294 7928 17590 7984
rect 17646 7928 17651 7984
rect 4294 7926 17651 7928
rect 17726 7986 17786 8198
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 17726 7926 27538 7986
rect 2865 7850 2931 7853
rect 4294 7850 4354 7926
rect 17585 7923 17651 7926
rect 2865 7848 4354 7850
rect 2865 7792 2870 7848
rect 2926 7792 4354 7848
rect 2865 7790 4354 7792
rect 4797 7850 4863 7853
rect 14917 7850 14983 7853
rect 4797 7848 14983 7850
rect 4797 7792 4802 7848
rect 4858 7792 14922 7848
rect 14978 7792 14983 7848
rect 4797 7790 14983 7792
rect 2865 7787 2931 7790
rect 4797 7787 4863 7790
rect 14917 7787 14983 7790
rect 1209 7714 1275 7717
rect 5257 7714 5323 7717
rect 1209 7712 5323 7714
rect 1209 7656 1214 7712
rect 1270 7656 5262 7712
rect 5318 7656 5323 7712
rect 1209 7654 5323 7656
rect 1209 7651 1275 7654
rect 5257 7651 5323 7654
rect 7281 7714 7347 7717
rect 11605 7714 11671 7717
rect 7281 7712 11671 7714
rect 7281 7656 7286 7712
rect 7342 7656 11610 7712
rect 11666 7656 11671 7712
rect 7281 7654 11671 7656
rect 7281 7651 7347 7654
rect 11605 7651 11671 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 6177 7578 6243 7581
rect 14181 7578 14247 7581
rect 6177 7576 14247 7578
rect 6177 7520 6182 7576
rect 6238 7520 14186 7576
rect 14242 7520 14247 7576
rect 6177 7518 14247 7520
rect 6177 7515 6243 7518
rect 14181 7515 14247 7518
rect 3509 7442 3575 7445
rect 10777 7442 10843 7445
rect 3509 7440 10843 7442
rect 3509 7384 3514 7440
rect 3570 7384 10782 7440
rect 10838 7384 10843 7440
rect 3509 7382 10843 7384
rect 3509 7379 3575 7382
rect 10777 7379 10843 7382
rect 15469 7442 15535 7445
rect 19517 7442 19583 7445
rect 15469 7440 19583 7442
rect 15469 7384 15474 7440
rect 15530 7384 19522 7440
rect 19578 7384 19583 7440
rect 15469 7382 19583 7384
rect 15469 7379 15535 7382
rect 19517 7379 19583 7382
rect 0 7306 480 7336
rect 8385 7306 8451 7309
rect 0 7304 8451 7306
rect 0 7248 8390 7304
rect 8446 7248 8451 7304
rect 0 7246 8451 7248
rect 0 7216 480 7246
rect 8385 7243 8451 7246
rect 9489 7306 9555 7309
rect 18045 7306 18111 7309
rect 9489 7304 18111 7306
rect 9489 7248 9494 7304
rect 9550 7248 18050 7304
rect 18106 7248 18111 7304
rect 9489 7246 18111 7248
rect 9489 7243 9555 7246
rect 18045 7243 18111 7246
rect 1577 7170 1643 7173
rect 3509 7170 3575 7173
rect 1577 7168 3575 7170
rect 1577 7112 1582 7168
rect 1638 7112 3514 7168
rect 3570 7112 3575 7168
rect 1577 7110 3575 7112
rect 1577 7107 1643 7110
rect 3509 7107 3575 7110
rect 3693 7170 3759 7173
rect 7373 7170 7439 7173
rect 3693 7168 7439 7170
rect 3693 7112 3698 7168
rect 3754 7112 7378 7168
rect 7434 7112 7439 7168
rect 3693 7110 7439 7112
rect 3693 7107 3759 7110
rect 7373 7107 7439 7110
rect 10685 7170 10751 7173
rect 12709 7170 12775 7173
rect 10685 7168 12775 7170
rect 10685 7112 10690 7168
rect 10746 7112 12714 7168
rect 12770 7112 12775 7168
rect 10685 7110 12775 7112
rect 10685 7107 10751 7110
rect 12709 7107 12775 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 27478 7064 27538 7926
rect 2497 7034 2563 7037
rect 3233 7034 3299 7037
rect 7005 7034 7071 7037
rect 2497 7032 3066 7034
rect 2497 6976 2502 7032
rect 2558 6976 3066 7032
rect 2497 6974 3066 6976
rect 2497 6971 2563 6974
rect 3006 6762 3066 6974
rect 3233 7032 7071 7034
rect 3233 6976 3238 7032
rect 3294 6976 7010 7032
rect 7066 6976 7071 7032
rect 3233 6974 7071 6976
rect 27478 6974 28000 7064
rect 3233 6971 3299 6974
rect 7005 6971 7071 6974
rect 27520 6944 28000 6974
rect 3601 6898 3667 6901
rect 8753 6898 8819 6901
rect 3601 6896 8819 6898
rect 3601 6840 3606 6896
rect 3662 6840 8758 6896
rect 8814 6840 8819 6896
rect 3601 6838 8819 6840
rect 3601 6835 3667 6838
rect 8753 6835 8819 6838
rect 10961 6898 11027 6901
rect 15561 6898 15627 6901
rect 10961 6896 15627 6898
rect 10961 6840 10966 6896
rect 11022 6840 15566 6896
rect 15622 6840 15627 6896
rect 10961 6838 15627 6840
rect 10961 6835 11027 6838
rect 15561 6835 15627 6838
rect 3693 6762 3759 6765
rect 3006 6760 3759 6762
rect 3006 6704 3698 6760
rect 3754 6704 3759 6760
rect 3006 6702 3759 6704
rect 3693 6699 3759 6702
rect 4153 6762 4219 6765
rect 5165 6762 5231 6765
rect 8293 6762 8359 6765
rect 4153 6760 8359 6762
rect 4153 6704 4158 6760
rect 4214 6704 5170 6760
rect 5226 6704 8298 6760
rect 8354 6704 8359 6760
rect 4153 6702 8359 6704
rect 4153 6699 4219 6702
rect 5165 6699 5231 6702
rect 8293 6699 8359 6702
rect 18045 6762 18111 6765
rect 27613 6762 27679 6765
rect 18045 6760 27679 6762
rect 18045 6704 18050 6760
rect 18106 6704 27618 6760
rect 27674 6704 27679 6760
rect 18045 6702 27679 6704
rect 18045 6699 18111 6702
rect 27613 6699 27679 6702
rect 0 6626 480 6656
rect 3785 6626 3851 6629
rect 0 6624 3851 6626
rect 0 6568 3790 6624
rect 3846 6568 3851 6624
rect 0 6566 3851 6568
rect 0 6536 480 6566
rect 3785 6563 3851 6566
rect 8017 6626 8083 6629
rect 11237 6626 11303 6629
rect 8017 6624 11303 6626
rect 8017 6568 8022 6624
rect 8078 6568 11242 6624
rect 11298 6568 11303 6624
rect 8017 6566 11303 6568
rect 8017 6563 8083 6566
rect 11237 6563 11303 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 2129 6490 2195 6493
rect 5073 6490 5139 6493
rect 2129 6488 5139 6490
rect 2129 6432 2134 6488
rect 2190 6432 5078 6488
rect 5134 6432 5139 6488
rect 2129 6430 5139 6432
rect 2129 6427 2195 6430
rect 5073 6427 5139 6430
rect 17902 6428 17908 6492
rect 17972 6490 17978 6492
rect 18321 6490 18387 6493
rect 17972 6488 18387 6490
rect 17972 6432 18326 6488
rect 18382 6432 18387 6488
rect 17972 6430 18387 6432
rect 17972 6428 17978 6430
rect 18321 6427 18387 6430
rect 6361 6354 6427 6357
rect 7373 6354 7439 6357
rect 18505 6354 18571 6357
rect 6361 6352 18571 6354
rect 6361 6296 6366 6352
rect 6422 6296 7378 6352
rect 7434 6296 18510 6352
rect 18566 6296 18571 6352
rect 6361 6294 18571 6296
rect 6361 6291 6427 6294
rect 7373 6291 7439 6294
rect 18505 6291 18571 6294
rect 1393 6218 1459 6221
rect 6913 6218 6979 6221
rect 1393 6216 6979 6218
rect 1393 6160 1398 6216
rect 1454 6160 6918 6216
rect 6974 6160 6979 6216
rect 1393 6158 6979 6160
rect 1393 6155 1459 6158
rect 6913 6155 6979 6158
rect 7189 6218 7255 6221
rect 19333 6218 19399 6221
rect 7189 6216 19399 6218
rect 7189 6160 7194 6216
rect 7250 6160 19338 6216
rect 19394 6160 19399 6216
rect 7189 6158 19399 6160
rect 7189 6155 7255 6158
rect 19333 6155 19399 6158
rect 0 6082 480 6112
rect 1761 6082 1827 6085
rect 0 6080 1827 6082
rect 0 6024 1766 6080
rect 1822 6024 1827 6080
rect 0 6022 1827 6024
rect 0 5992 480 6022
rect 1761 6019 1827 6022
rect 2957 6082 3023 6085
rect 4797 6082 4863 6085
rect 2957 6080 4863 6082
rect 2957 6024 2962 6080
rect 3018 6024 4802 6080
rect 4858 6024 4863 6080
rect 2957 6022 4863 6024
rect 2957 6019 3023 6022
rect 4797 6019 4863 6022
rect 5073 6082 5139 6085
rect 10133 6082 10199 6085
rect 5073 6080 10199 6082
rect 5073 6024 5078 6080
rect 5134 6024 10138 6080
rect 10194 6024 10199 6080
rect 5073 6022 10199 6024
rect 5073 6019 5139 6022
rect 10133 6019 10199 6022
rect 11881 6082 11947 6085
rect 13997 6082 14063 6085
rect 11881 6080 14063 6082
rect 11881 6024 11886 6080
rect 11942 6024 14002 6080
rect 14058 6024 14063 6080
rect 11881 6022 14063 6024
rect 11881 6019 11947 6022
rect 13997 6019 14063 6022
rect 16481 6082 16547 6085
rect 19425 6082 19491 6085
rect 16481 6080 19491 6082
rect 16481 6024 16486 6080
rect 16542 6024 19430 6080
rect 19486 6024 19491 6080
rect 16481 6022 19491 6024
rect 16481 6019 16547 6022
rect 19425 6019 19491 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 2313 5946 2379 5949
rect 7281 5946 7347 5949
rect 2313 5944 7347 5946
rect 2313 5888 2318 5944
rect 2374 5888 7286 5944
rect 7342 5888 7347 5944
rect 2313 5886 7347 5888
rect 2313 5883 2379 5886
rect 7281 5883 7347 5886
rect 14549 5946 14615 5949
rect 18689 5946 18755 5949
rect 14549 5944 18755 5946
rect 14549 5888 14554 5944
rect 14610 5888 18694 5944
rect 18750 5888 18755 5944
rect 14549 5886 18755 5888
rect 14549 5883 14615 5886
rect 18689 5883 18755 5886
rect 4613 5810 4679 5813
rect 6494 5810 6500 5812
rect 4613 5808 6500 5810
rect 4613 5752 4618 5808
rect 4674 5752 6500 5808
rect 4613 5750 6500 5752
rect 4613 5747 4679 5750
rect 6494 5748 6500 5750
rect 6564 5748 6570 5812
rect 6821 5810 6887 5813
rect 9765 5810 9831 5813
rect 6821 5808 9831 5810
rect 6821 5752 6826 5808
rect 6882 5752 9770 5808
rect 9826 5752 9831 5808
rect 6821 5750 9831 5752
rect 6821 5747 6887 5750
rect 9765 5747 9831 5750
rect 9949 5810 10015 5813
rect 20989 5810 21055 5813
rect 9949 5808 21055 5810
rect 9949 5752 9954 5808
rect 10010 5752 20994 5808
rect 21050 5752 21055 5808
rect 9949 5750 21055 5752
rect 9949 5747 10015 5750
rect 20989 5747 21055 5750
rect 4061 5674 4127 5677
rect 7833 5674 7899 5677
rect 4061 5672 7899 5674
rect 4061 5616 4066 5672
rect 4122 5616 7838 5672
rect 7894 5616 7899 5672
rect 4061 5614 7899 5616
rect 4061 5611 4127 5614
rect 7833 5611 7899 5614
rect 8017 5674 8083 5677
rect 9673 5674 9739 5677
rect 20345 5674 20411 5677
rect 8017 5672 20411 5674
rect 8017 5616 8022 5672
rect 8078 5616 9678 5672
rect 9734 5616 20350 5672
rect 20406 5616 20411 5672
rect 8017 5614 20411 5616
rect 8017 5611 8083 5614
rect 9673 5611 9739 5614
rect 20345 5611 20411 5614
rect 2773 5540 2839 5541
rect 2773 5536 2820 5540
rect 2884 5538 2890 5540
rect 11513 5538 11579 5541
rect 12157 5538 12223 5541
rect 14641 5538 14707 5541
rect 2773 5480 2778 5536
rect 2773 5476 2820 5480
rect 2884 5478 2930 5538
rect 11513 5536 14707 5538
rect 11513 5480 11518 5536
rect 11574 5480 12162 5536
rect 12218 5480 14646 5536
rect 14702 5480 14707 5536
rect 11513 5478 14707 5480
rect 2884 5476 2890 5478
rect 2773 5475 2839 5476
rect 11513 5475 11579 5478
rect 12157 5475 12223 5478
rect 14641 5475 14707 5478
rect 15377 5538 15443 5541
rect 19425 5538 19491 5541
rect 15377 5536 19491 5538
rect 15377 5480 15382 5536
rect 15438 5480 19430 5536
rect 19486 5480 19491 5536
rect 15377 5478 19491 5480
rect 15377 5475 15443 5478
rect 19425 5475 19491 5478
rect 5610 5472 5930 5473
rect 0 5402 480 5432
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 6085 5404 6151 5405
rect 6085 5402 6132 5404
rect 0 5342 4906 5402
rect 6040 5400 6132 5402
rect 6040 5344 6090 5400
rect 6040 5342 6132 5344
rect 0 5312 480 5342
rect 4846 5266 4906 5342
rect 6085 5340 6132 5342
rect 6196 5340 6202 5404
rect 6729 5402 6795 5405
rect 11513 5402 11579 5405
rect 13537 5402 13603 5405
rect 6729 5400 11579 5402
rect 6729 5344 6734 5400
rect 6790 5344 11518 5400
rect 11574 5344 11579 5400
rect 6729 5342 11579 5344
rect 6085 5339 6151 5340
rect 6729 5339 6795 5342
rect 11513 5339 11579 5342
rect 11654 5400 13603 5402
rect 11654 5344 13542 5400
rect 13598 5344 13603 5400
rect 11654 5342 13603 5344
rect 11513 5266 11579 5269
rect 4846 5264 11579 5266
rect 4846 5208 11518 5264
rect 11574 5208 11579 5264
rect 4846 5206 11579 5208
rect 11513 5203 11579 5206
rect 1945 5130 2011 5133
rect 2681 5130 2747 5133
rect 1945 5128 2747 5130
rect 1945 5072 1950 5128
rect 2006 5072 2686 5128
rect 2742 5072 2747 5128
rect 1945 5070 2747 5072
rect 1945 5067 2011 5070
rect 2681 5067 2747 5070
rect 3233 5130 3299 5133
rect 4153 5130 4219 5133
rect 3233 5128 4219 5130
rect 3233 5072 3238 5128
rect 3294 5072 4158 5128
rect 4214 5072 4219 5128
rect 3233 5070 4219 5072
rect 3233 5067 3299 5070
rect 4153 5067 4219 5070
rect 4613 5130 4679 5133
rect 11654 5130 11714 5342
rect 13537 5339 13603 5342
rect 16389 5402 16455 5405
rect 22461 5402 22527 5405
rect 16389 5400 22527 5402
rect 16389 5344 16394 5400
rect 16450 5344 22466 5400
rect 22522 5344 22527 5400
rect 16389 5342 22527 5344
rect 16389 5339 16455 5342
rect 22461 5339 22527 5342
rect 11789 5266 11855 5269
rect 13629 5266 13695 5269
rect 11789 5264 13695 5266
rect 11789 5208 11794 5264
rect 11850 5208 13634 5264
rect 13690 5208 13695 5264
rect 11789 5206 13695 5208
rect 11789 5203 11855 5206
rect 13629 5203 13695 5206
rect 4613 5128 11714 5130
rect 4613 5072 4618 5128
rect 4674 5072 11714 5128
rect 4613 5070 11714 5072
rect 18597 5130 18663 5133
rect 20713 5132 20779 5133
rect 20662 5130 20668 5132
rect 18597 5128 20178 5130
rect 18597 5072 18602 5128
rect 18658 5072 20178 5128
rect 18597 5070 20178 5072
rect 20622 5070 20668 5130
rect 20732 5128 20779 5132
rect 20774 5072 20779 5128
rect 4613 5067 4679 5070
rect 18597 5067 18663 5070
rect 13077 4994 13143 4997
rect 15929 4994 15995 4997
rect 13077 4992 15995 4994
rect 13077 4936 13082 4992
rect 13138 4936 15934 4992
rect 15990 4936 15995 4992
rect 13077 4934 15995 4936
rect 20118 4994 20178 5070
rect 20662 5068 20668 5070
rect 20732 5068 20779 5072
rect 20713 5067 20779 5068
rect 27061 4994 27127 4997
rect 20118 4992 27127 4994
rect 20118 4936 27066 4992
rect 27122 4936 27127 4992
rect 20118 4934 27127 4936
rect 13077 4931 13143 4934
rect 15929 4931 15995 4934
rect 27061 4931 27127 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 10869 4858 10935 4861
rect 12433 4858 12499 4861
rect 18321 4858 18387 4861
rect 10869 4856 18387 4858
rect 10869 4800 10874 4856
rect 10930 4800 12438 4856
rect 12494 4800 18326 4856
rect 18382 4800 18387 4856
rect 10869 4798 18387 4800
rect 10869 4795 10935 4798
rect 12433 4795 12499 4798
rect 18321 4795 18387 4798
rect 0 4722 480 4752
rect 3877 4722 3943 4725
rect 0 4720 3943 4722
rect 0 4664 3882 4720
rect 3938 4664 3943 4720
rect 0 4662 3943 4664
rect 0 4632 480 4662
rect 3877 4659 3943 4662
rect 5441 4722 5507 4725
rect 14273 4722 14339 4725
rect 5441 4720 14339 4722
rect 5441 4664 5446 4720
rect 5502 4664 14278 4720
rect 14334 4664 14339 4720
rect 5441 4662 14339 4664
rect 5441 4659 5507 4662
rect 14273 4659 14339 4662
rect 14641 4722 14707 4725
rect 19609 4722 19675 4725
rect 14641 4720 19675 4722
rect 14641 4664 14646 4720
rect 14702 4664 19614 4720
rect 19670 4664 19675 4720
rect 14641 4662 19675 4664
rect 14641 4659 14707 4662
rect 19609 4659 19675 4662
rect 2497 4586 2563 4589
rect 3969 4586 4035 4589
rect 19885 4586 19951 4589
rect 2497 4584 19951 4586
rect 2497 4528 2502 4584
rect 2558 4528 3974 4584
rect 4030 4528 19890 4584
rect 19946 4528 19951 4584
rect 2497 4526 19951 4528
rect 2497 4523 2563 4526
rect 3969 4523 4035 4526
rect 19885 4523 19951 4526
rect 18505 4450 18571 4453
rect 21081 4450 21147 4453
rect 18505 4448 21147 4450
rect 18505 4392 18510 4448
rect 18566 4392 21086 4448
rect 21142 4392 21147 4448
rect 18505 4390 21147 4392
rect 18505 4387 18571 4390
rect 21081 4387 21147 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 2589 4314 2655 4317
rect 5441 4314 5507 4317
rect 11329 4314 11395 4317
rect 2589 4312 5507 4314
rect 2589 4256 2594 4312
rect 2650 4256 5446 4312
rect 5502 4256 5507 4312
rect 2589 4254 5507 4256
rect 2589 4251 2655 4254
rect 5441 4251 5507 4254
rect 6686 4312 11395 4314
rect 6686 4256 11334 4312
rect 11390 4256 11395 4312
rect 6686 4254 11395 4256
rect 0 4178 480 4208
rect 6686 4178 6746 4254
rect 11329 4251 11395 4254
rect 11513 4314 11579 4317
rect 12617 4314 12683 4317
rect 11513 4312 12683 4314
rect 11513 4256 11518 4312
rect 11574 4256 12622 4312
rect 12678 4256 12683 4312
rect 11513 4254 12683 4256
rect 11513 4251 11579 4254
rect 12617 4251 12683 4254
rect 17677 4314 17743 4317
rect 19425 4314 19491 4317
rect 17677 4312 19491 4314
rect 17677 4256 17682 4312
rect 17738 4256 19430 4312
rect 19486 4256 19491 4312
rect 17677 4254 19491 4256
rect 17677 4251 17743 4254
rect 19425 4251 19491 4254
rect 21449 4178 21515 4181
rect 0 4118 6746 4178
rect 6870 4176 21515 4178
rect 6870 4120 21454 4176
rect 21510 4120 21515 4176
rect 6870 4118 21515 4120
rect 0 4088 480 4118
rect 6453 4042 6519 4045
rect 6870 4042 6930 4118
rect 21449 4115 21515 4118
rect 6453 4040 6930 4042
rect 6453 3984 6458 4040
rect 6514 3984 6930 4040
rect 6453 3982 6930 3984
rect 15561 4042 15627 4045
rect 20621 4042 20687 4045
rect 21633 4042 21699 4045
rect 15561 4040 20178 4042
rect 15561 3984 15566 4040
rect 15622 3984 20178 4040
rect 15561 3982 20178 3984
rect 6453 3979 6519 3982
rect 15561 3979 15627 3982
rect 2589 3906 2655 3909
rect 7097 3906 7163 3909
rect 8293 3906 8359 3909
rect 9673 3906 9739 3909
rect 2589 3904 6378 3906
rect 2589 3848 2594 3904
rect 2650 3848 6378 3904
rect 2589 3846 6378 3848
rect 2589 3843 2655 3846
rect 657 3770 723 3773
rect 6177 3770 6243 3773
rect 657 3768 6243 3770
rect 657 3712 662 3768
rect 718 3712 6182 3768
rect 6238 3712 6243 3768
rect 657 3710 6243 3712
rect 6318 3770 6378 3846
rect 7097 3904 9739 3906
rect 7097 3848 7102 3904
rect 7158 3848 8298 3904
rect 8354 3848 9678 3904
rect 9734 3848 9739 3904
rect 7097 3846 9739 3848
rect 7097 3843 7163 3846
rect 8293 3843 8359 3846
rect 9673 3843 9739 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 7649 3770 7715 3773
rect 6318 3768 7715 3770
rect 6318 3712 7654 3768
rect 7710 3712 7715 3768
rect 6318 3710 7715 3712
rect 657 3707 723 3710
rect 6177 3707 6243 3710
rect 7649 3707 7715 3710
rect 1393 3634 1459 3637
rect 5717 3634 5783 3637
rect 8201 3634 8267 3637
rect 12709 3634 12775 3637
rect 1393 3632 5642 3634
rect 1393 3576 1398 3632
rect 1454 3576 5642 3632
rect 1393 3574 5642 3576
rect 1393 3571 1459 3574
rect 0 3498 480 3528
rect 3509 3498 3575 3501
rect 0 3496 3575 3498
rect 0 3440 3514 3496
rect 3570 3440 3575 3496
rect 0 3438 3575 3440
rect 5582 3498 5642 3574
rect 5717 3632 8267 3634
rect 5717 3576 5722 3632
rect 5778 3576 8206 3632
rect 8262 3576 8267 3632
rect 5717 3574 8267 3576
rect 5717 3571 5783 3574
rect 8201 3571 8267 3574
rect 10182 3632 12775 3634
rect 10182 3576 12714 3632
rect 12770 3576 12775 3632
rect 10182 3574 12775 3576
rect 7833 3498 7899 3501
rect 5582 3496 7899 3498
rect 5582 3440 7838 3496
rect 7894 3440 7899 3496
rect 5582 3438 7899 3440
rect 0 3408 480 3438
rect 3509 3435 3575 3438
rect 7833 3435 7899 3438
rect 9029 3498 9095 3501
rect 10182 3498 10242 3574
rect 12709 3571 12775 3574
rect 13261 3634 13327 3637
rect 20118 3634 20178 3982
rect 20621 4040 21699 4042
rect 20621 3984 20626 4040
rect 20682 3984 21638 4040
rect 21694 3984 21699 4040
rect 20621 3982 21699 3984
rect 20621 3979 20687 3982
rect 21633 3979 21699 3982
rect 26509 3634 26575 3637
rect 13261 3632 19810 3634
rect 13261 3576 13266 3632
rect 13322 3576 19810 3632
rect 13261 3574 19810 3576
rect 20118 3632 26575 3634
rect 20118 3576 26514 3632
rect 26570 3576 26575 3632
rect 20118 3574 26575 3576
rect 13261 3571 13327 3574
rect 13353 3498 13419 3501
rect 9029 3496 10242 3498
rect 9029 3440 9034 3496
rect 9090 3440 10242 3496
rect 9029 3438 10242 3440
rect 10366 3496 13419 3498
rect 10366 3440 13358 3496
rect 13414 3440 13419 3496
rect 10366 3438 13419 3440
rect 9029 3435 9095 3438
rect 2497 3362 2563 3365
rect 4153 3362 4219 3365
rect 2497 3360 4219 3362
rect 2497 3304 2502 3360
rect 2558 3304 4158 3360
rect 4214 3304 4219 3360
rect 2497 3302 4219 3304
rect 2497 3299 2563 3302
rect 4153 3299 4219 3302
rect 9305 3362 9371 3365
rect 10366 3362 10426 3438
rect 13353 3435 13419 3438
rect 14825 3498 14891 3501
rect 19609 3498 19675 3501
rect 14825 3496 19675 3498
rect 14825 3440 14830 3496
rect 14886 3440 19614 3496
rect 19670 3440 19675 3496
rect 14825 3438 19675 3440
rect 19750 3498 19810 3574
rect 26509 3571 26575 3574
rect 23657 3498 23723 3501
rect 19750 3496 23723 3498
rect 19750 3440 23662 3496
rect 23718 3440 23723 3496
rect 19750 3438 23723 3440
rect 14825 3435 14891 3438
rect 19609 3435 19675 3438
rect 23657 3435 23723 3438
rect 9305 3360 10426 3362
rect 9305 3304 9310 3360
rect 9366 3304 10426 3360
rect 9305 3302 10426 3304
rect 12433 3362 12499 3365
rect 12709 3362 12775 3365
rect 12433 3360 12775 3362
rect 12433 3304 12438 3360
rect 12494 3304 12714 3360
rect 12770 3304 12775 3360
rect 12433 3302 12775 3304
rect 9305 3299 9371 3302
rect 12433 3299 12499 3302
rect 12709 3299 12775 3302
rect 19241 3362 19307 3365
rect 19241 3360 23490 3362
rect 19241 3304 19246 3360
rect 19302 3304 23490 3360
rect 19241 3302 23490 3304
rect 19241 3299 19307 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 6177 3226 6243 3229
rect 14273 3226 14339 3229
rect 16205 3226 16271 3229
rect 22369 3226 22435 3229
rect 6177 3224 14842 3226
rect 6177 3168 6182 3224
rect 6238 3168 14278 3224
rect 14334 3168 14842 3224
rect 6177 3166 14842 3168
rect 6177 3163 6243 3166
rect 14273 3163 14339 3166
rect 2313 3090 2379 3093
rect 4613 3090 4679 3093
rect 2313 3088 4679 3090
rect 2313 3032 2318 3088
rect 2374 3032 4618 3088
rect 4674 3032 4679 3088
rect 2313 3030 4679 3032
rect 2313 3027 2379 3030
rect 4613 3027 4679 3030
rect 9305 3090 9371 3093
rect 12433 3090 12499 3093
rect 9305 3088 12499 3090
rect 9305 3032 9310 3088
rect 9366 3032 12438 3088
rect 12494 3032 12499 3088
rect 9305 3030 12499 3032
rect 14782 3090 14842 3166
rect 16205 3224 22435 3226
rect 16205 3168 16210 3224
rect 16266 3168 22374 3224
rect 22430 3168 22435 3224
rect 16205 3166 22435 3168
rect 16205 3163 16271 3166
rect 22369 3163 22435 3166
rect 17861 3090 17927 3093
rect 14782 3088 17927 3090
rect 14782 3032 17866 3088
rect 17922 3032 17927 3088
rect 14782 3030 17927 3032
rect 23430 3090 23490 3302
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 24853 3090 24919 3093
rect 23430 3088 24919 3090
rect 23430 3032 24858 3088
rect 24914 3032 24919 3088
rect 23430 3030 24919 3032
rect 9305 3027 9371 3030
rect 12433 3027 12499 3030
rect 17861 3027 17927 3030
rect 24853 3027 24919 3030
rect 2037 2954 2103 2957
rect 6545 2954 6611 2957
rect 2037 2952 6611 2954
rect 2037 2896 2042 2952
rect 2098 2896 6550 2952
rect 6606 2896 6611 2952
rect 2037 2894 6611 2896
rect 2037 2891 2103 2894
rect 6545 2891 6611 2894
rect 11421 2954 11487 2957
rect 18137 2954 18203 2957
rect 11421 2952 18203 2954
rect 11421 2896 11426 2952
rect 11482 2896 18142 2952
rect 18198 2896 18203 2952
rect 11421 2894 18203 2896
rect 11421 2891 11487 2894
rect 18137 2891 18203 2894
rect 18965 2954 19031 2957
rect 22185 2954 22251 2957
rect 18965 2952 22251 2954
rect 18965 2896 18970 2952
rect 19026 2896 22190 2952
rect 22246 2896 22251 2952
rect 18965 2894 22251 2896
rect 18965 2891 19031 2894
rect 22185 2891 22251 2894
rect 0 2818 480 2848
rect 8569 2818 8635 2821
rect 0 2816 8635 2818
rect 0 2760 8574 2816
rect 8630 2760 8635 2816
rect 0 2758 8635 2760
rect 0 2728 480 2758
rect 8569 2755 8635 2758
rect 10869 2818 10935 2821
rect 19241 2818 19307 2821
rect 10869 2816 19307 2818
rect 10869 2760 10874 2816
rect 10930 2760 19246 2816
rect 19302 2760 19307 2816
rect 10869 2758 19307 2760
rect 10869 2755 10935 2758
rect 19241 2755 19307 2758
rect 20345 2818 20411 2821
rect 22093 2818 22159 2821
rect 20345 2816 22159 2818
rect 20345 2760 20350 2816
rect 20406 2760 22098 2816
rect 22154 2760 22159 2816
rect 20345 2758 22159 2760
rect 20345 2755 20411 2758
rect 22093 2755 22159 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 2865 2682 2931 2685
rect 3182 2682 3188 2684
rect 2865 2680 3188 2682
rect 2865 2624 2870 2680
rect 2926 2624 3188 2680
rect 2865 2622 3188 2624
rect 2865 2619 2931 2622
rect 3182 2620 3188 2622
rect 3252 2620 3258 2684
rect 3509 2682 3575 2685
rect 8385 2682 8451 2685
rect 3509 2680 8451 2682
rect 3509 2624 3514 2680
rect 3570 2624 8390 2680
rect 8446 2624 8451 2680
rect 3509 2622 8451 2624
rect 3509 2619 3575 2622
rect 8385 2619 8451 2622
rect 13813 2682 13879 2685
rect 18321 2682 18387 2685
rect 13813 2680 18387 2682
rect 13813 2624 13818 2680
rect 13874 2624 18326 2680
rect 18382 2624 18387 2680
rect 13813 2622 18387 2624
rect 13813 2619 13879 2622
rect 18321 2619 18387 2622
rect 10041 2546 10107 2549
rect 11145 2546 11211 2549
rect 10041 2544 11211 2546
rect 10041 2488 10046 2544
rect 10102 2488 11150 2544
rect 11206 2488 11211 2544
rect 10041 2486 11211 2488
rect 10041 2483 10107 2486
rect 11145 2483 11211 2486
rect 14181 2546 14247 2549
rect 17677 2546 17743 2549
rect 14181 2544 17743 2546
rect 14181 2488 14186 2544
rect 14242 2488 17682 2544
rect 17738 2488 17743 2544
rect 14181 2486 17743 2488
rect 14181 2483 14247 2486
rect 17677 2483 17743 2486
rect 17861 2546 17927 2549
rect 21265 2546 21331 2549
rect 17861 2544 21331 2546
rect 17861 2488 17866 2544
rect 17922 2488 21270 2544
rect 21326 2488 21331 2544
rect 17861 2486 21331 2488
rect 17861 2483 17927 2486
rect 21265 2483 21331 2486
rect 3325 2410 3391 2413
rect 10777 2410 10843 2413
rect 3325 2408 10843 2410
rect 3325 2352 3330 2408
rect 3386 2352 10782 2408
rect 10838 2352 10843 2408
rect 3325 2350 10843 2352
rect 3325 2347 3391 2350
rect 10777 2347 10843 2350
rect 14365 2410 14431 2413
rect 25405 2410 25471 2413
rect 14365 2408 25471 2410
rect 14365 2352 14370 2408
rect 14426 2352 25410 2408
rect 25466 2352 25471 2408
rect 14365 2350 25471 2352
rect 14365 2347 14431 2350
rect 25405 2347 25471 2350
rect 0 2274 480 2304
rect 1577 2274 1643 2277
rect 0 2272 1643 2274
rect 0 2216 1582 2272
rect 1638 2216 1643 2272
rect 0 2214 1643 2216
rect 0 2184 480 2214
rect 1577 2211 1643 2214
rect 3141 2274 3207 2277
rect 5349 2274 5415 2277
rect 3141 2272 5415 2274
rect 3141 2216 3146 2272
rect 3202 2216 5354 2272
rect 5410 2216 5415 2272
rect 3141 2214 5415 2216
rect 3141 2211 3207 2214
rect 5349 2211 5415 2214
rect 5993 2274 6059 2277
rect 14549 2274 14615 2277
rect 5993 2272 14615 2274
rect 5993 2216 5998 2272
rect 6054 2216 14554 2272
rect 14610 2216 14615 2272
rect 5993 2214 14615 2216
rect 5993 2211 6059 2214
rect 14549 2211 14615 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 3785 2002 3851 2005
rect 14181 2002 14247 2005
rect 3785 2000 14247 2002
rect 3785 1944 3790 2000
rect 3846 1944 14186 2000
rect 14242 1944 14247 2000
rect 3785 1942 14247 1944
rect 3785 1939 3851 1942
rect 14181 1939 14247 1942
rect 14641 2002 14707 2005
rect 18045 2002 18111 2005
rect 14641 2000 18111 2002
rect 14641 1944 14646 2000
rect 14702 1944 18050 2000
rect 18106 1944 18111 2000
rect 14641 1942 18111 1944
rect 14641 1939 14707 1942
rect 18045 1939 18111 1942
rect 4521 1866 4587 1869
rect 1166 1864 4587 1866
rect 1166 1808 4526 1864
rect 4582 1808 4587 1864
rect 1166 1806 4587 1808
rect 0 1594 480 1624
rect 1166 1594 1226 1806
rect 4521 1803 4587 1806
rect 2497 1730 2563 1733
rect 19977 1730 20043 1733
rect 24025 1732 24091 1733
rect 2497 1728 20043 1730
rect 2497 1672 2502 1728
rect 2558 1672 19982 1728
rect 20038 1672 20043 1728
rect 2497 1670 20043 1672
rect 2497 1667 2563 1670
rect 19977 1667 20043 1670
rect 23974 1668 23980 1732
rect 24044 1730 24091 1732
rect 24044 1728 24136 1730
rect 24086 1672 24136 1728
rect 24044 1670 24136 1672
rect 24044 1668 24091 1670
rect 24025 1667 24091 1668
rect 0 1534 1226 1594
rect 1393 1594 1459 1597
rect 3325 1594 3391 1597
rect 1393 1592 3391 1594
rect 1393 1536 1398 1592
rect 1454 1536 3330 1592
rect 3386 1536 3391 1592
rect 1393 1534 3391 1536
rect 0 1504 480 1534
rect 1393 1531 1459 1534
rect 3325 1531 3391 1534
rect 3601 1594 3667 1597
rect 6085 1594 6151 1597
rect 3601 1592 6151 1594
rect 3601 1536 3606 1592
rect 3662 1536 6090 1592
rect 6146 1536 6151 1592
rect 3601 1534 6151 1536
rect 3601 1531 3667 1534
rect 6085 1531 6151 1534
rect 13169 1594 13235 1597
rect 14733 1594 14799 1597
rect 19885 1594 19951 1597
rect 13169 1592 19951 1594
rect 13169 1536 13174 1592
rect 13230 1536 14738 1592
rect 14794 1536 19890 1592
rect 19946 1536 19951 1592
rect 13169 1534 19951 1536
rect 13169 1531 13235 1534
rect 14733 1531 14799 1534
rect 19885 1531 19951 1534
rect 4061 1458 4127 1461
rect 11513 1458 11579 1461
rect 4061 1456 11579 1458
rect 4061 1400 4066 1456
rect 4122 1400 11518 1456
rect 11574 1400 11579 1456
rect 4061 1398 11579 1400
rect 4061 1395 4127 1398
rect 11513 1395 11579 1398
rect 17861 1458 17927 1461
rect 24209 1458 24275 1461
rect 17861 1456 24275 1458
rect 17861 1400 17866 1456
rect 17922 1400 24214 1456
rect 24270 1400 24275 1456
rect 17861 1398 24275 1400
rect 17861 1395 17927 1398
rect 24209 1395 24275 1398
rect 6269 1322 6335 1325
rect 19425 1322 19491 1325
rect 6269 1320 19491 1322
rect 6269 1264 6274 1320
rect 6330 1264 19430 1320
rect 19486 1264 19491 1320
rect 6269 1262 19491 1264
rect 6269 1259 6335 1262
rect 19425 1259 19491 1262
rect 3969 1186 4035 1189
rect 10041 1186 10107 1189
rect 3969 1184 10107 1186
rect 3969 1128 3974 1184
rect 4030 1128 10046 1184
rect 10102 1128 10107 1184
rect 3969 1126 10107 1128
rect 3969 1123 4035 1126
rect 10041 1123 10107 1126
rect 4613 1050 4679 1053
rect 21817 1050 21883 1053
rect 4613 1048 21883 1050
rect 4613 992 4618 1048
rect 4674 992 21822 1048
rect 21878 992 21883 1048
rect 4613 990 21883 992
rect 4613 987 4679 990
rect 21817 987 21883 990
rect 0 914 480 944
rect 9673 914 9739 917
rect 20529 914 20595 917
rect 0 912 9739 914
rect 0 856 9678 912
rect 9734 856 9739 912
rect 0 854 9739 856
rect 0 824 480 854
rect 9673 851 9739 854
rect 9814 912 20595 914
rect 9814 856 20534 912
rect 20590 856 20595 912
rect 9814 854 20595 856
rect 4153 778 4219 781
rect 9814 778 9874 854
rect 20529 851 20595 854
rect 4153 776 9874 778
rect 4153 720 4158 776
rect 4214 720 9874 776
rect 4153 718 9874 720
rect 10041 778 10107 781
rect 22185 778 22251 781
rect 10041 776 22251 778
rect 10041 720 10046 776
rect 10102 720 22190 776
rect 22246 720 22251 776
rect 10041 718 22251 720
rect 4153 715 4219 718
rect 10041 715 10107 718
rect 22185 715 22251 718
rect 2589 642 2655 645
rect 20253 642 20319 645
rect 2589 640 20319 642
rect 2589 584 2594 640
rect 2650 584 20258 640
rect 20314 584 20319 640
rect 2589 582 20319 584
rect 2589 579 2655 582
rect 20253 579 20319 582
rect 0 370 480 400
rect 4061 370 4127 373
rect 0 368 4127 370
rect 0 312 4066 368
rect 4122 312 4127 368
rect 0 310 4127 312
rect 0 280 480 310
rect 4061 307 4127 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 6500 12608 6564 12612
rect 6500 12552 6550 12608
rect 6550 12552 6564 12608
rect 6500 12548 6564 12552
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 6132 9148 6196 9212
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 3188 8332 3252 8396
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 17908 6428 17972 6492
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 6500 5748 6564 5812
rect 2820 5536 2884 5540
rect 2820 5480 2834 5536
rect 2834 5480 2884 5536
rect 2820 5476 2884 5480
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 6132 5400 6196 5404
rect 6132 5344 6146 5400
rect 6146 5344 6196 5400
rect 6132 5340 6196 5344
rect 20668 5128 20732 5132
rect 20668 5072 20718 5128
rect 20718 5072 20732 5128
rect 20668 5068 20732 5072
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 3188 2620 3252 2684
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 23980 1728 24044 1732
rect 23980 1672 24030 1728
rect 24030 1672 24044 1728
rect 23980 1668 24044 1672
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 6499 12612 6565 12613
rect 6499 12548 6500 12612
rect 6564 12548 6565 12612
rect 6499 12547 6565 12548
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 6131 9212 6197 9213
rect 6131 9148 6132 9212
rect 6196 9148 6197 9212
rect 6131 9147 6197 9148
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 3187 8396 3253 8397
rect 3187 8332 3188 8396
rect 3252 8332 3253 8396
rect 3187 8331 3253 8332
rect 2819 5540 2885 5541
rect 2819 5476 2820 5540
rect 2884 5476 2885 5540
rect 2819 5475 2885 5476
rect 2822 5218 2882 5475
rect 3190 2685 3250 8331
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 6134 6578 6194 9147
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 6134 5405 6194 6342
rect 6502 5813 6562 12547
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 6499 5812 6565 5813
rect 6499 5748 6500 5812
rect 6564 5748 6565 5812
rect 6499 5747 6565 5748
rect 6131 5404 6197 5405
rect 6131 5340 6132 5404
rect 6196 5340 6197 5404
rect 6131 5339 6197 5340
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 3187 2684 3253 2685
rect 3187 2620 3188 2684
rect 3252 2620 3253 2684
rect 3187 2619 3253 2620
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 6502 1818 6562 5747
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 2734 4982 2970 5218
rect 6046 6342 6282 6578
rect 17822 6492 18058 6578
rect 17822 6428 17908 6492
rect 17908 6428 17972 6492
rect 17972 6428 18058 6492
rect 17822 6342 18058 6428
rect 20582 5132 20818 5218
rect 20582 5068 20668 5132
rect 20668 5068 20732 5132
rect 20732 5068 20818 5132
rect 20582 4982 20818 5068
rect 6414 1582 6650 1818
rect 23894 1732 24130 1818
rect 23894 1668 23980 1732
rect 23980 1668 24044 1732
rect 24044 1668 24130 1732
rect 23894 1582 24130 1668
<< metal5 >>
rect 6004 6578 18100 6620
rect 6004 6342 6046 6578
rect 6282 6342 17822 6578
rect 18058 6342 18100 6578
rect 6004 6300 18100 6342
rect 2692 5218 20860 5260
rect 2692 4982 2734 5218
rect 2970 4982 20582 5218
rect 20818 4982 20860 5218
rect 2692 4940 20860 4982
rect 6372 1818 24172 1860
rect 6372 1582 6414 1818
rect 6650 1582 23894 1818
rect 24130 1582 24172 1818
rect 6372 1540 24172 1582
use scs8hd_fill_2  FILLER_1_8 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__S tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_conb_1  _049_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_7.mux_l2_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_25
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_21
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_7.scs8hd_dfxbp_1_2_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_55 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6164 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_48
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_54
timestamp 1586364061
transform 1 0 6072 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_58
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_88
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_86
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_82
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_11.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_111
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _073_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_115
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_115
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_119
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_11.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_146
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _074_
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_150
timestamp 1586364061
transform 1 0 14904 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_169
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_173
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_179
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_203
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _083_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20792 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_track_33.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_223
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _078_
timestamp 1586364061
transform 1 0 21252 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_224
timestamp 1586364061
transform 1 0 21712 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_231
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _077_
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _076_
timestamp 1586364061
transform 1 0 22448 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_236
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_0_240 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_conb_1  _051_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_253
timestamp 1586364061
transform 1 0 24380 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _088_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_248 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23920 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_257
timestamp 1586364061
transform 1 0 24748 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_260
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_272
timestamp 1586364061
transform 1 0 26128 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_276
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use scs8hd_conb_1  _033_
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_7.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_12
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_50
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_61
timestamp 1586364061
transform 1 0 6716 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_78
timestamp 1586364061
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _072_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_82
timestamp 1586364061
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_86
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_101
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_15.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_124
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_128
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_19.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_152
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_160
timestamp 1586364061
transform 1 0 15824 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_164
timestamp 1586364061
transform 1 0 16192 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_2  _075_
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_187
timestamp 1586364061
transform 1 0 18308 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_191
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _079_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_203
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_207
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_2  _086_
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 21804 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_219
timestamp 1586364061
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_223
timestamp 1586364061
transform 1 0 21620 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_231
timestamp 1586364061
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_243
timestamp 1586364061
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_255
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_267
timestamp 1586364061
transform 1 0 25668 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_7.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_23
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 1786 592
use scs8hd_buf_4  mux_left_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_68
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_72
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_99
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_15.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 1786 592
use scs8hd_buf_4  mux_left_track_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_120
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_129
timestamp 1586364061
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_133
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_157
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16284 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_161
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_174
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_178
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18768 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_182
timestamp 1586364061
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_190
timestamp 1586364061
transform 1 0 18584 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_194
timestamp 1586364061
transform 1 0 18952 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_198
timestamp 1586364061
transform 1 0 19320 0 1 3808
box -38 -48 314 592
use scs8hd_buf_2  _080_
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_203
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_211
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_215
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _052_
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 314 592
use scs8hd_buf_2  _084_
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_223
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_227
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_3_234
timestamp 1586364061
transform 1 0 22632 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_242
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_conb_1  _032_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_7.mux_l1_in_3_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_3_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_49
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_45
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_58
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_11.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11316 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_15.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_122
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_126
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15548 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_139
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_147
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_19.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16928 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_170
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_193
timestamp 1586364061
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_197
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _082_
timestamp 1586364061
transform 1 0 19596 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _087_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20148 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_205
timestamp 1586364061
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_209
timestamp 1586364061
transform 1 0 20332 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_219
timestamp 1586364061
transform 1 0 21252 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_223
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_235
timestamp 1586364061
transform 1 0 22724 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_259
timestamp 1586364061
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_271
timestamp 1586364061
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_10
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_2_
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_23
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _071_
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_44
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_52
timestamp 1586364061
transform 1 0 5888 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6900 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_72
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_76
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _067_
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_117
timestamp 1586364061
transform 1 0 11868 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _065_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_131
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_158
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_19.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_162
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_19.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_19.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_210
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_218
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_230
timestamp 1586364061
transform 1 0 22264 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_242
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _070_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_12
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_10
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 1786 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_35
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_49
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_52
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_75
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _069_
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 1786 592
use scs8hd_buf_4  mux_left_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_99
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_104
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_103
timestamp 1586364061
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_21.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1786 592
use scs8hd_mux2_2  mux_left_track_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_126
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_130
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_143
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_146
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_147
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_152
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_151
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_21.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_21.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15824 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_173
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_169
timestamp 1586364061
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_175
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_169
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_19.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17572 0 -1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_21.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_198
timestamp 1586364061
transform 1 0 19320 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_207
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_203
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_215
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_203
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_227
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_239
timestamp 1586364061
transform 1 0 23092 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_243
timestamp 1586364061
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_conb_1  _030_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_55
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_59
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_2  _068_
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_71
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_75
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_99
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_13.mux_l3_in_0_
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_103
timestamp 1586364061
transform 1 0 10580 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_13.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _090_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_148
timestamp 1586364061
transform 1 0 14720 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_21.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_162
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _053_
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_185
timestamp 1586364061
transform 1 0 18124 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_189
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_196
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_200
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_212
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_32
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_55
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_13.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_96
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_23.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_129
timestamp 1586364061
transform 1 0 12972 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_21.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_23.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13892 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_148
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_152
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_165
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_169
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_173
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_177
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _050_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_181
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_187
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_191
timestamp 1586364061
transform 1 0 18676 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_227
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_239
timestamp 1586364061
transform 1 0 23092 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_8
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_10_40
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_60
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_78
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_82
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_86
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_90
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_99
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_103
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_23.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_121
timestamp 1586364061
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_140
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_148
timestamp 1586364061
transform 1 0 14720 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _028_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_157
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_23.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_161
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_184
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_208 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_3_
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 866 592
use scs8hd_buf_4  mux_left_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_9
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_13
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_26
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_30
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 590 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_3_
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_70
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_87
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_104
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_23.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _027_
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_162
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_166
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_181
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_11
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_47
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_51
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _061_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_87
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_101
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_23.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_131
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 314 592
use scs8hd_buf_2  _093_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_158
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _091_
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15824 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_162
timestamp 1586364061
transform 1 0 16008 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_170
timestamp 1586364061
transform 1 0 16744 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_4  mux_left_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_11
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 590 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_29
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_25
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _066_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_14_40
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4968 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_57
timestamp 1586364061
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_53
timestamp 1586364061
transform 1 0 5980 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_67
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_buf_4  mux_left_track_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 590 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_71
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _062_
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_87
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10120 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_105
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_111
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use scs8hd_conb_1  _031_
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_115
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _059_
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_137
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_134
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_130
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 1786 592
use scs8hd_buf_2  _092_
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_157
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_140
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_2  _089_
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_161
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_169
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_175
timestamp 1586364061
transform 1 0 17204 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_181
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_187
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_199
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1472 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_13
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_17
timestamp 1586364061
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 1786 592
use scs8hd_buf_2  _063_
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_44
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_52
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_56
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_4_
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_60
timestamp 1586364061
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_73
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 1786 592
use scs8hd_conb_1  _029_
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_100
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_104
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 12512 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_174
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_182
timestamp 1586364061
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4140 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_21
timestamp 1586364061
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_25
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_42
timestamp 1586364061
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_63
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_74
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13524 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_133
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_149
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_173
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_185
timestamp 1586364061
transform 1 0 18124 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_197
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_209
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_conb_1  _045_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 1786 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_6
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_10
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_33
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_37
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_41
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_81
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_85
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_88
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _046_
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_105
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_116
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 1786 592
use scs8hd_buf_4  mux_bottom_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_146
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_151
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_202
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_214
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_226
timestamp 1586364061
transform 1 0 21896 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_17_238
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4232 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_43
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_47
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use scs8hd_conb_1  _048_
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_70
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_78
timestamp 1586364061
transform 1 0 8280 0 -1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_5_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_82
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_86
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_3_
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_136
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_140
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_144
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_175
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_187
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_2  _081_
timestamp 1586364061
transform 1 0 19504 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_204
timestamp 1586364061
transform 1 0 19872 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_212
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _064_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_28
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_24
timestamp 1586364061
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_41
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_45
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_45
timestamp 1586364061
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _058_
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 406 592
use scs8hd_buf_2  _056_
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_59
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_76
timestamp 1586364061
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_72
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_79
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_86
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_99
timestamp 1586364061
transform 1 0 10212 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_96
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_100
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10304 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 866 592
use scs8hd_decap_6  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_113
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_127
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_148
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_139
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_160
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_164
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_177
timestamp 1586364061
transform 1 0 17388 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_4  mux_bottom_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_188
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_191
timestamp 1586364061
transform 1 0 18676 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_195
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_215
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_207
timestamp 1586364061
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_213
timestamp 1586364061
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_227
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_239
timestamp 1586364061
transform 1 0 23092 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_243
timestamp 1586364061
transform 1 0 23460 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_14
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _054_
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_41
timestamp 1586364061
transform 1 0 4876 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_45
timestamp 1586364061
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_81
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_85
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_93
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_101
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_146
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_165
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_169
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_181
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 1932 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_11
timestamp 1586364061
transform 1 0 2116 0 -1 14688
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_51
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_60
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use scs8hd_conb_1  _043_
timestamp 1586364061
transform 1 0 9752 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10212 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_90
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_97
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_101
timestamp 1586364061
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_124
timestamp 1586364061
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_128
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_2  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_158
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_162
timestamp 1586364061
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_182
timestamp 1586364061
transform 1 0 17848 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_194
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_2  _060_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_17
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_28
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_32
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_45
timestamp 1586364061
transform 1 0 5244 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_49
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_76
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_80
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_84
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12512 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_133
timestamp 1586364061
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_137
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_141
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_145
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_149
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_172
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_176
timestamp 1586364061
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 18216 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 18584 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_180
timestamp 1586364061
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_188
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_192
timestamp 1586364061
transform 1 0 18768 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_204
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_216
timestamp 1586364061
transform 1 0 20976 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_228
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_buf_2  _055_
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 406 592
use scs8hd_buf_2  _057_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 2300 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_11
timestamp 1586364061
transform 1 0 2116 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use scs8hd_conb_1  _041_
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_24_39
timestamp 1586364061
transform 1 0 4692 0 -1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_43
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_87
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11592 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_112
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_116
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_126
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_132
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_150
timestamp 1586364061
transform 1 0 14904 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 774 592
use scs8hd_buf_2  _085_
timestamp 1586364061
transform 1 0 18400 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_180
timestamp 1586364061
transform 1 0 17664 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_192
timestamp 1586364061
transform 1 0 18768 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_204
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_212
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l1_in_2_
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_18
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _044_
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_22
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_33
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_36
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_40
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_32.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _042_
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_101
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_105
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_112
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_116
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13340 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_131
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16652 0 1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_166
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_6  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_13
timestamp 1586364061
transform 1 0 2300 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_11
timestamp 1586364061
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 2300 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_24
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_20
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_32
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_46
timestamp 1586364061
transform 1 0 5336 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_42
timestamp 1586364061
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_32.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 5520 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_57
timestamp 1586364061
transform 1 0 6348 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_61
timestamp 1586364061
transform 1 0 6716 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_89
timestamp 1586364061
transform 1 0 9292 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_85
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_81
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l1_in_3_
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_111
timestamp 1586364061
transform 1 0 11316 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_136
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_127
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 130 592
use scs8hd_conb_1  _047_
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_149
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_153
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_175
timestamp 1586364061
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_160
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_164
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_168
timestamp 1586364061
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_187
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_180
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_199
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_11
timestamp 1586364061
transform 1 0 2116 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_36
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_28_42
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_32.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_62
timestamp 1586364061
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_66
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_79
timestamp 1586364061
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_83
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_87
timestamp 1586364061
transform 1 0 9108 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 10212 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 12052 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11684 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_101
timestamp 1586364061
transform 1 0 10396 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_113
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_121
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_139
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_143
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_147
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_167
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_179
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_191
timestamp 1586364061
transform 1 0 18676 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_203
timestamp 1586364061
transform 1 0 19780 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_211
timestamp 1586364061
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_conb_1  _037_
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_14
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_18
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _038_
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_41
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_45
timestamp 1586364061
transform 1 0 5244 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_32.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_75
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_79
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_6_
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_84
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l1_in_2_
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_track_16.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_149
timestamp 1586364061
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_153
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_166
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_182
timestamp 1586364061
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_29_216
timestamp 1586364061
transform 1 0 20976 0 1 17952
box -38 -48 314 592
use scs8hd_buf_4  mux_top_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21252 0 1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_225
timestamp 1586364061
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_229
timestamp 1586364061
transform 1 0 22172 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_241
timestamp 1586364061
transform 1 0 23276 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_mux2_2  mux_top_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_11
timestamp 1586364061
transform 1 0 2116 0 -1 19040
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 590 592
use scs8hd_mux2_2  mux_top_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6348 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_51
timestamp 1586364061
transform 1 0 5796 0 -1 19040
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_72
timestamp 1586364061
transform 1 0 7728 0 -1 19040
box -38 -48 1142 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_87
timestamp 1586364061
transform 1 0 9108 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_conb_1  _035_
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_113
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_16.mux_l1_in_3_
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_167
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_179
timestamp 1586364061
transform 1 0 17572 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_191
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_203
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_211
timestamp 1586364061
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_3_
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_21
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_25
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_38
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_42
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_46
timestamp 1586364061
transform 1 0 5336 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5520 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_54
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_50
timestamp 1586364061
transform 1 0 5704 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 406 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 8924 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_81
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_142
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_146
timestamp 1586364061
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_166
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_170
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_174
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_182
timestamp 1586364061
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_198
timestamp 1586364061
transform 1 0 19320 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 1142 592
use scs8hd_buf_2  _097_
timestamp 1586364061
transform 1 0 22264 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_222
timestamp 1586364061
transform 1 0 21528 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_234
timestamp 1586364061
transform 1 0 22632 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_238
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_11
timestamp 1586364061
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use scs8hd_conb_1  _034_
timestamp 1586364061
transform 1 0 1840 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 2300 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 2668 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4140 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3036 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6440 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_42
timestamp 1586364061
transform 1 0 4968 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_46
timestamp 1586364061
transform 1 0 5336 0 -1 20128
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7084 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_60
timestamp 1586364061
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 130 592
use scs8hd_conb_1  _036_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_96
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11132 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_100
timestamp 1586364061
transform 1 0 10304 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_104
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_107
timestamp 1586364061
transform 1 0 10948 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 13432 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_128
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 15640 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14904 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16192 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 16008 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_160
timestamp 1586364061
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19136 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_32_183
timestamp 1586364061
transform 1 0 17940 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_195
timestamp 1586364061
transform 1 0 19044 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 1564 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 1840 0 -1 21216
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 1472 0 1 20128
box -38 -48 866 592
use scs8hd_decap_4  FILLER_34_17
timestamp 1586364061
transform 1 0 2668 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_17
timestamp 1586364061
transform 1 0 2668 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_13
timestamp 1586364061
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_28
timestamp 1586364061
transform 1 0 3680 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_23
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3496 0 -1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 4232 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_30
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_34
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4600 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_36
timestamp 1586364061
transform 1 0 4416 0 -1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_47
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_40
timestamp 1586364061
transform 1 0 4784 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7176 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8372 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_60
timestamp 1586364061
transform 1 0 6624 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_64
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_77
timestamp 1586364061
transform 1 0 8188 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_81
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_85
timestamp 1586364061
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9292 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 8740 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_91
timestamp 1586364061
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_102
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_106
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_112
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_120
timestamp 1586364061
transform 1 0 12144 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_16.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_133
timestamp 1586364061
transform 1 0 13340 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_138
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_132
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 13156 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_4  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_146
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_142
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_152
timestamp 1586364061
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_149
timestamp 1586364061
transform 1 0 14812 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14904 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 15640 0 -1 21216
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_33_169
timestamp 1586364061
transform 1 0 16652 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_177
timestamp 1586364061
transform 1 0 17388 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_4  mux_top_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_181
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_190
timestamp 1586364061
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_194
timestamp 1586364061
transform 1 0 18952 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_189
timestamp 1586364061
transform 1 0 18492 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_206
timestamp 1586364061
transform 1 0 20056 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_214
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_217
timestamp 1586364061
transform 1 0 21068 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_201
timestamp 1586364061
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_229
timestamp 1586364061
transform 1 0 22172 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_219
timestamp 1586364061
transform 1 0 21252 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_231
timestamp 1586364061
transform 1 0 22356 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_241
timestamp 1586364061
transform 1 0 23276 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_243
timestamp 1586364061
transform 1 0 23460 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_255
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_34_267
timestamp 1586364061
transform 1 0 25668 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_18
timestamp 1586364061
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 3496 0 1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 3312 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_22
timestamp 1586364061
transform 1 0 3128 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_45
timestamp 1586364061
transform 1 0 5244 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_49
timestamp 1586364061
transform 1 0 5612 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_71
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_79
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 406 592
use scs8hd_mux2_2  mux_top_track_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 8832 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_83
timestamp 1586364061
transform 1 0 8740 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_99
timestamp 1586364061
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_112
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_6_
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 13800 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_136
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 14904 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 14720 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14352 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_140
timestamp 1586364061
transform 1 0 13984 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_146
timestamp 1586364061
transform 1 0 14536 0 1 21216
box -38 -48 222 592
use scs8hd_conb_1  _040_
timestamp 1586364061
transform 1 0 16468 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 16928 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15916 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 16284 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_163
timestamp 1586364061
transform 1 0 16100 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_170
timestamp 1586364061
transform 1 0 16744 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_174
timestamp 1586364061
transform 1 0 17112 0 1 21216
box -38 -48 774 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 18124 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 18676 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_182
timestamp 1586364061
transform 1 0 17848 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_189
timestamp 1586364061
transform 1 0 18492 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_193
timestamp 1586364061
transform 1 0 18860 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_205
timestamp 1586364061
transform 1 0 19964 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_217
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_229
timestamp 1586364061
transform 1 0 22172 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_35_241
timestamp 1586364061
transform 1 0 23276 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_mux2_2  mux_top_track_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 1840 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_7
timestamp 1586364061
transform 1 0 1748 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_10
timestamp 1586364061
transform 1 0 2024 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_36
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 406 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5060 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4876 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_40
timestamp 1586364061
transform 1 0 4784 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_52
timestamp 1586364061
transform 1 0 5888 0 -1 22304
box -38 -48 774 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6624 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_69
timestamp 1586364061
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_73
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_77
timestamp 1586364061
transform 1 0 8188 0 -1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9936 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_85
timestamp 1586364061
transform 1 0 8924 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_98
timestamp 1586364061
transform 1 0 10120 0 -1 22304
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_5_
timestamp 1586364061
transform 1 0 13156 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_123
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_127
timestamp 1586364061
transform 1 0 12788 0 -1 22304
box -38 -48 406 592
use scs8hd_mux2_2  mux_top_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_140
timestamp 1586364061
transform 1 0 13984 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_144
timestamp 1586364061
transform 1 0 14352 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_150
timestamp 1586364061
transform 1 0 14904 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_2  _096_
timestamp 1586364061
transform 1 0 16836 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 16284 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_163
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_167
timestamp 1586364061
transform 1 0 16468 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_175
timestamp 1586364061
transform 1 0 17204 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_187
timestamp 1586364061
transform 1 0 18308 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_199
timestamp 1586364061
transform 1 0 19412 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_36_211
timestamp 1586364061
transform 1 0 20516 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2300 0 1 22304
box -38 -48 1786 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_9
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_32
timestamp 1586364061
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_36
timestamp 1586364061
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4784 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_49
timestamp 1586364061
transform 1 0 5612 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7176 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6992 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_79
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_83
timestamp 1586364061
transform 1 0 8740 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_89
timestamp 1586364061
transform 1 0 9292 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12052 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11684 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 10948 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_105
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_109
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_117
timestamp 1586364061
transform 1 0 11868 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 1786 592
use scs8hd_buf_4  mux_top_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_121
timestamp 1586364061
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_129
timestamp 1586364061
transform 1 0 12972 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_133
timestamp 1586364061
transform 1 0 13340 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_156
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_160
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_168
timestamp 1586364061
transform 1 0 16560 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_173
timestamp 1586364061
transform 1 0 17020 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 18216 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_181
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_188
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_200
timestamp 1586364061
transform 1 0 19504 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_212
timestamp 1586364061
transform 1 0 20608 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 21804 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_224
timestamp 1586364061
transform 1 0 21712 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_227
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_239
timestamp 1586364061
transform 1 0 23092 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_243
timestamp 1586364061
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 1932 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_11
timestamp 1586364061
transform 1 0 2116 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4324 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4692 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_37
timestamp 1586364061
transform 1 0 4508 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_3_
timestamp 1586364061
transform 1 0 5520 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5060 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_41
timestamp 1586364061
transform 1 0 4876 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_45
timestamp 1586364061
transform 1 0 5244 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_57
timestamp 1586364061
transform 1 0 6348 0 -1 23392
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7084 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_61
timestamp 1586364061
transform 1 0 6716 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_64
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_98
timestamp 1586364061
transform 1 0 10120 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12052 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 10304 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_111
timestamp 1586364061
transform 1 0 11316 0 -1 23392
box -38 -48 774 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13064 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_128
timestamp 1586364061
transform 1 0 12880 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_132
timestamp 1586364061
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 16836 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_38_163
timestamp 1586364061
transform 1 0 16100 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_38_175
timestamp 1586364061
transform 1 0 17204 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 17940 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_187
timestamp 1586364061
transform 1 0 18308 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_199
timestamp 1586364061
transform 1 0 19412 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_38_211
timestamp 1586364061
transform 1 0 20516 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 21804 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_223
timestamp 1586364061
transform 1 0 21620 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_229
timestamp 1586364061
transform 1 0 22172 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_241
timestamp 1586364061
transform 1 0 23276 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_253
timestamp 1586364061
transform 1 0 24380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_265
timestamp 1586364061
transform 1 0 25484 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_273
timestamp 1586364061
transform 1 0 26220 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1472 0 -1 24480
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 866 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2760 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_12
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_16
timestamp 1586364061
transform 1 0 2576 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2944 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4324 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_23
timestamp 1586364061
transform 1 0 3220 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_47
timestamp 1586364061
transform 1 0 5428 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_43
timestamp 1586364061
transform 1 0 5060 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5244 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5612 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4876 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_50
timestamp 1586364061
transform 1 0 5704 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_55
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5796 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5980 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_66
timestamp 1586364061
transform 1 0 7176 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_62
timestamp 1586364061
transform 1 0 6808 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6992 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_79
timestamp 1586364061
transform 1 0 8372 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_75
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_71
timestamp 1586364061
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7544 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 10028 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 590 592
use scs8hd_decap_8  FILLER_40_83
timestamp 1586364061
transform 1 0 8740 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_91
timestamp 1586364061
transform 1 0 9476 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_6  FILLER_40_99
timestamp 1586364061
transform 1 0 10212 0 -1 24480
box -38 -48 590 592
use scs8hd_conb_1  _039_
timestamp 1586364061
transform 1 0 10856 0 1 23392
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 10672 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_109
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_113
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_124
timestamp 1586364061
transform 1 0 12512 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_40_136
timestamp 1586364061
transform 1 0 13616 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_146
timestamp 1586364061
transform 1 0 14536 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13892 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_156
timestamp 1586364061
transform 1 0 15456 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_152
timestamp 1586364061
transform 1 0 15088 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14904 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_158
timestamp 1586364061
transform 1 0 15640 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_4  mux_top_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15548 0 1 23392
box -38 -48 590 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_163
timestamp 1586364061
transform 1 0 16100 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_168
timestamp 1586364061
transform 1 0 16560 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_170
timestamp 1586364061
transform 1 0 16744 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_194
timestamp 1586364061
transform 1 0 18952 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_197
timestamp 1586364061
transform 1 0 19228 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_193
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 18492 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_182
timestamp 1586364061
transform 1 0 17848 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_204
timestamp 1586364061
transform 1 0 19872 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_205
timestamp 1586364061
transform 1 0 19964 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 19412 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 19596 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 19504 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_212
timestamp 1586364061
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_217
timestamp 1586364061
transform 1 0 21068 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_209
timestamp 1586364061
transform 1 0 20332 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 20700 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 21252 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_221
timestamp 1586364061
transform 1 0 21436 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_229
timestamp 1586364061
transform 1 0 22172 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_233
timestamp 1586364061
transform 1 0 22540 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_241
timestamp 1586364061
transform 1 0 23276 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 1564 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_7
timestamp 1586364061
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_11
timestamp 1586364061
transform 1 0 2116 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_19
timestamp 1586364061
transform 1 0 2852 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 3956 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3772 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3036 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_23
timestamp 1586364061
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5336 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5704 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_40
timestamp 1586364061
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_44
timestamp 1586364061
transform 1 0 5152 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_48
timestamp 1586364061
transform 1 0 5520 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_52
timestamp 1586364061
transform 1 0 5888 0 1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_41_58
timestamp 1586364061
transform 1 0 6440 0 1 24480
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7176 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 8188 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6992 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_75
timestamp 1586364061
transform 1 0 8004 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_79
timestamp 1586364061
transform 1 0 8372 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 10028 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 9844 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 8556 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_83
timestamp 1586364061
transform 1 0 8740 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_87
timestamp 1586364061
transform 1 0 9108 0 1 24480
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 11040 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 11408 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_106
timestamp 1586364061
transform 1 0 10856 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 406 592
use scs8hd_buf_4  mux_top_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12972 0 1 24480
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12788 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _095_
timestamp 1586364061
transform 1 0 15364 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 13892 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 14812 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_141
timestamp 1586364061
transform 1 0 14076 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_151
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 15916 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_163
timestamp 1586364061
transform 1 0 16100 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_175
timestamp 1586364061
transform 1 0 17204 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4324 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 7544 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7176 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_42_68
timestamp 1586364061
transform 1 0 7360 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_79
timestamp 1586364061
transform 1 0 8372 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 10028 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_91
timestamp 1586364061
transform 1 0 9476 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_42_99
timestamp 1586364061
transform 1 0 10212 0 -1 25568
box -38 -48 590 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_4_
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_8  FILLER_42_114
timestamp 1586364061
transform 1 0 11592 0 -1 25568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_122
timestamp 1586364061
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _094_
timestamp 1586364061
transform 1 0 13892 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_143
timestamp 1586364061
transform 1 0 14260 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_34_
port 0 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_35_
port 1 nsew default input
rlabel metal2 s 1214 0 1270 480 6 bottom_left_grid_pin_36_
port 2 nsew default input
rlabel metal2 s 1766 0 1822 480 6 bottom_left_grid_pin_37_
port 3 nsew default input
rlabel metal2 s 2318 0 2374 480 6 bottom_left_grid_pin_38_
port 4 nsew default input
rlabel metal2 s 2870 0 2926 480 6 bottom_left_grid_pin_39_
port 5 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_40_
port 6 nsew default input
rlabel metal2 s 3882 0 3938 480 6 bottom_left_grid_pin_41_
port 7 nsew default input
rlabel metal2 s 25962 0 26018 480 6 bottom_right_grid_pin_1_
port 8 nsew default input
rlabel metal3 s 0 25712 480 25832 6 ccff_head
port 9 nsew default input
rlabel metal3 s 0 26256 480 26376 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 12928 480 13048 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 21904 480 22024 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 22448 480 22568 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 23128 480 23248 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 23808 480 23928 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 24352 480 24472 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 25032 480 25152 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 15512 480 15632 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 16736 480 16856 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 17416 480 17536 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 18096 480 18216 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 18640 480 18760 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 6536 480 6656 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 7216 480 7336 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 7896 480 8016 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 9120 480 9240 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 11704 480 11824 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 1504 480 1624 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 2184 480 2304 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 2728 480 2848 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 4088 480 4208 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 4632 480 4752 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 5312 480 5432 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 5992 480 6112 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal2 s 4434 0 4490 480 6 chany_bottom_in[0]
port 51 nsew default input
rlabel metal2 s 9862 0 9918 480 6 chany_bottom_in[10]
port 52 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[11]
port 53 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[12]
port 54 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chany_bottom_in[13]
port 55 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[14]
port 56 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[15]
port 57 nsew default input
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_in[16]
port 58 nsew default input
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_in[17]
port 59 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[18]
port 60 nsew default input
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_in[19]
port 61 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[1]
port 62 nsew default input
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_in[2]
port 63 nsew default input
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_in[3]
port 64 nsew default input
rlabel metal2 s 6642 0 6698 480 6 chany_bottom_in[4]
port 65 nsew default input
rlabel metal2 s 7194 0 7250 480 6 chany_bottom_in[5]
port 66 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[6]
port 67 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[7]
port 68 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chany_bottom_in[8]
port 69 nsew default input
rlabel metal2 s 9310 0 9366 480 6 chany_bottom_in[9]
port 70 nsew default input
rlabel metal2 s 15198 0 15254 480 6 chany_bottom_out[0]
port 71 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 chany_bottom_out[10]
port 72 nsew default tristate
rlabel metal2 s 21178 0 21234 480 6 chany_bottom_out[11]
port 73 nsew default tristate
rlabel metal2 s 21638 0 21694 480 6 chany_bottom_out[12]
port 74 nsew default tristate
rlabel metal2 s 22190 0 22246 480 6 chany_bottom_out[13]
port 75 nsew default tristate
rlabel metal2 s 22742 0 22798 480 6 chany_bottom_out[14]
port 76 nsew default tristate
rlabel metal2 s 23294 0 23350 480 6 chany_bottom_out[15]
port 77 nsew default tristate
rlabel metal2 s 23846 0 23902 480 6 chany_bottom_out[16]
port 78 nsew default tristate
rlabel metal2 s 24398 0 24454 480 6 chany_bottom_out[17]
port 79 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 chany_bottom_out[18]
port 80 nsew default tristate
rlabel metal2 s 25410 0 25466 480 6 chany_bottom_out[19]
port 81 nsew default tristate
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_out[1]
port 82 nsew default tristate
rlabel metal2 s 16302 0 16358 480 6 chany_bottom_out[2]
port 83 nsew default tristate
rlabel metal2 s 16854 0 16910 480 6 chany_bottom_out[3]
port 84 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[4]
port 85 nsew default tristate
rlabel metal2 s 17866 0 17922 480 6 chany_bottom_out[5]
port 86 nsew default tristate
rlabel metal2 s 18418 0 18474 480 6 chany_bottom_out[6]
port 87 nsew default tristate
rlabel metal2 s 18970 0 19026 480 6 chany_bottom_out[7]
port 88 nsew default tristate
rlabel metal2 s 19522 0 19578 480 6 chany_bottom_out[8]
port 89 nsew default tristate
rlabel metal2 s 20074 0 20130 480 6 chany_bottom_out[9]
port 90 nsew default tristate
rlabel metal2 s 4526 27520 4582 28000 6 chany_top_in[0]
port 91 nsew default input
rlabel metal2 s 10046 27520 10102 28000 6 chany_top_in[10]
port 92 nsew default input
rlabel metal2 s 10598 27520 10654 28000 6 chany_top_in[11]
port 93 nsew default input
rlabel metal2 s 11150 27520 11206 28000 6 chany_top_in[12]
port 94 nsew default input
rlabel metal2 s 11702 27520 11758 28000 6 chany_top_in[13]
port 95 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_in[14]
port 96 nsew default input
rlabel metal2 s 12806 27520 12862 28000 6 chany_top_in[15]
port 97 nsew default input
rlabel metal2 s 13358 27520 13414 28000 6 chany_top_in[16]
port 98 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[17]
port 99 nsew default input
rlabel metal2 s 14370 27520 14426 28000 6 chany_top_in[18]
port 100 nsew default input
rlabel metal2 s 14922 27520 14978 28000 6 chany_top_in[19]
port 101 nsew default input
rlabel metal2 s 5078 27520 5134 28000 6 chany_top_in[1]
port 102 nsew default input
rlabel metal2 s 5630 27520 5686 28000 6 chany_top_in[2]
port 103 nsew default input
rlabel metal2 s 6182 27520 6238 28000 6 chany_top_in[3]
port 104 nsew default input
rlabel metal2 s 6734 27520 6790 28000 6 chany_top_in[4]
port 105 nsew default input
rlabel metal2 s 7286 27520 7342 28000 6 chany_top_in[5]
port 106 nsew default input
rlabel metal2 s 7838 27520 7894 28000 6 chany_top_in[6]
port 107 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[7]
port 108 nsew default input
rlabel metal2 s 8942 27520 8998 28000 6 chany_top_in[8]
port 109 nsew default input
rlabel metal2 s 9494 27520 9550 28000 6 chany_top_in[9]
port 110 nsew default input
rlabel metal2 s 15474 27520 15530 28000 6 chany_top_out[0]
port 111 nsew default tristate
rlabel metal2 s 20994 27520 21050 28000 6 chany_top_out[10]
port 112 nsew default tristate
rlabel metal2 s 21546 27520 21602 28000 6 chany_top_out[11]
port 113 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[12]
port 114 nsew default tristate
rlabel metal2 s 22650 27520 22706 28000 6 chany_top_out[13]
port 115 nsew default tristate
rlabel metal2 s 23202 27520 23258 28000 6 chany_top_out[14]
port 116 nsew default tristate
rlabel metal2 s 23754 27520 23810 28000 6 chany_top_out[15]
port 117 nsew default tristate
rlabel metal2 s 24306 27520 24362 28000 6 chany_top_out[16]
port 118 nsew default tristate
rlabel metal2 s 24858 27520 24914 28000 6 chany_top_out[17]
port 119 nsew default tristate
rlabel metal2 s 25410 27520 25466 28000 6 chany_top_out[18]
port 120 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[19]
port 121 nsew default tristate
rlabel metal2 s 16026 27520 16082 28000 6 chany_top_out[1]
port 122 nsew default tristate
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[2]
port 123 nsew default tristate
rlabel metal2 s 17130 27520 17186 28000 6 chany_top_out[3]
port 124 nsew default tristate
rlabel metal2 s 17682 27520 17738 28000 6 chany_top_out[4]
port 125 nsew default tristate
rlabel metal2 s 18234 27520 18290 28000 6 chany_top_out[5]
port 126 nsew default tristate
rlabel metal2 s 18786 27520 18842 28000 6 chany_top_out[6]
port 127 nsew default tristate
rlabel metal2 s 19338 27520 19394 28000 6 chany_top_out[7]
port 128 nsew default tristate
rlabel metal2 s 19890 27520 19946 28000 6 chany_top_out[8]
port 129 nsew default tristate
rlabel metal2 s 20442 27520 20498 28000 6 chany_top_out[9]
port 130 nsew default tristate
rlabel metal3 s 27520 6944 28000 7064 6 left_top_grid_pin_42_
port 131 nsew default input
rlabel metal3 s 0 26936 480 27056 6 left_top_grid_pin_43_
port 132 nsew default input
rlabel metal2 s 27066 27520 27122 28000 6 left_top_grid_pin_44_
port 133 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_45_
port 134 nsew default input
rlabel metal2 s 26514 0 26570 480 6 left_top_grid_pin_46_
port 135 nsew default input
rlabel metal2 s 27066 0 27122 480 6 left_top_grid_pin_47_
port 136 nsew default input
rlabel metal2 s 27618 27520 27674 28000 6 left_top_grid_pin_48_
port 137 nsew default input
rlabel metal3 s 27520 20952 28000 21072 6 left_top_grid_pin_49_
port 138 nsew default input
rlabel metal2 s 27618 0 27674 480 6 prog_clk
port 139 nsew default input
rlabel metal2 s 202 27520 258 28000 6 top_left_grid_pin_34_
port 140 nsew default input
rlabel metal2 s 662 27520 718 28000 6 top_left_grid_pin_35_
port 141 nsew default input
rlabel metal2 s 1214 27520 1270 28000 6 top_left_grid_pin_36_
port 142 nsew default input
rlabel metal2 s 1766 27520 1822 28000 6 top_left_grid_pin_37_
port 143 nsew default input
rlabel metal2 s 2318 27520 2374 28000 6 top_left_grid_pin_38_
port 144 nsew default input
rlabel metal2 s 2870 27520 2926 28000 6 top_left_grid_pin_39_
port 145 nsew default input
rlabel metal2 s 3422 27520 3478 28000 6 top_left_grid_pin_40_
port 146 nsew default input
rlabel metal2 s 3974 27520 4030 28000 6 top_left_grid_pin_41_
port 147 nsew default input
rlabel metal2 s 26514 27520 26570 28000 6 top_right_grid_pin_1_
port 148 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 149 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
