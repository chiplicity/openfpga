* NGSPICE file created from grid_clb.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_sdfxbp_1 abstract view
.subckt scs8hd_sdfxbp_1 CLK D Q QN SCD SCE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_1 abstract view
.subckt scs8hd_or2_1 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_clkbuf_16 abstract view
.subckt scs8hd_clkbuf_16 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_clkbuf_1 abstract view
.subckt scs8hd_clkbuf_1 A X vgnd vpwr
.ends

.subckt grid_clb Test_en bottom_width_0_height_0__pin_16_ bottom_width_0_height_0__pin_17_
+ bottom_width_0_height_0__pin_18_ bottom_width_0_height_0__pin_19_ bottom_width_0_height_0__pin_20_
+ bottom_width_0_height_0__pin_21_ bottom_width_0_height_0__pin_22_ bottom_width_0_height_0__pin_23_
+ bottom_width_0_height_0__pin_24_ bottom_width_0_height_0__pin_25_ bottom_width_0_height_0__pin_26_
+ bottom_width_0_height_0__pin_27_ bottom_width_0_height_0__pin_28_ bottom_width_0_height_0__pin_29_
+ bottom_width_0_height_0__pin_30_ bottom_width_0_height_0__pin_31_ bottom_width_0_height_0__pin_42_lower
+ bottom_width_0_height_0__pin_42_upper bottom_width_0_height_0__pin_43_lower bottom_width_0_height_0__pin_43_upper
+ bottom_width_0_height_0__pin_44_lower bottom_width_0_height_0__pin_44_upper bottom_width_0_height_0__pin_45_lower
+ bottom_width_0_height_0__pin_45_upper bottom_width_0_height_0__pin_46_lower bottom_width_0_height_0__pin_46_upper
+ bottom_width_0_height_0__pin_47_lower bottom_width_0_height_0__pin_47_upper bottom_width_0_height_0__pin_48_lower
+ bottom_width_0_height_0__pin_48_upper bottom_width_0_height_0__pin_49_lower bottom_width_0_height_0__pin_49_upper
+ bottom_width_0_height_0__pin_50_ bottom_width_0_height_0__pin_51_ ccff_head ccff_tail
+ clk left_width_0_height_0__pin_52_ prog_clk right_width_0_height_0__pin_0_ right_width_0_height_0__pin_10_
+ right_width_0_height_0__pin_11_ right_width_0_height_0__pin_12_ right_width_0_height_0__pin_13_
+ right_width_0_height_0__pin_14_ right_width_0_height_0__pin_15_ right_width_0_height_0__pin_1_
+ right_width_0_height_0__pin_2_ right_width_0_height_0__pin_34_lower right_width_0_height_0__pin_34_upper
+ right_width_0_height_0__pin_35_lower right_width_0_height_0__pin_35_upper right_width_0_height_0__pin_36_lower
+ right_width_0_height_0__pin_36_upper right_width_0_height_0__pin_37_lower right_width_0_height_0__pin_37_upper
+ right_width_0_height_0__pin_38_lower right_width_0_height_0__pin_38_upper right_width_0_height_0__pin_39_lower
+ right_width_0_height_0__pin_39_upper right_width_0_height_0__pin_3_ right_width_0_height_0__pin_40_lower
+ right_width_0_height_0__pin_40_upper right_width_0_height_0__pin_41_lower right_width_0_height_0__pin_41_upper
+ right_width_0_height_0__pin_4_ right_width_0_height_0__pin_5_ right_width_0_height_0__pin_6_
+ right_width_0_height_0__pin_7_ right_width_0_height_0__pin_8_ right_width_0_height_0__pin_9_
+ top_width_0_height_0__pin_32_ top_width_0_height_0__pin_33_ vpwr vgnd
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_277 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _62_/HI
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_406 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _36_/HI
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_43_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_239 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_5_332 vgnd vpwr scs8hd_decap_4
XFILLER_36_269 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_8_181 vpwr vgnd scs8hd_fill_2
XFILLER_59_306 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_39 vgnd vpwr scs8hd_decap_12
XFILLER_42_239 vgnd vpwr scs8hd_decap_6
XFILLER_27_225 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_6_118 vgnd vpwr scs8hd_decap_8
XFILLER_10_125 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_58_383 vgnd vpwr scs8hd_decap_12
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_41_250 vpwr vgnd scs8hd_fill_2
XFILLER_33_239 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_162 vpwr vgnd scs8hd_fill_2
XFILLER_64_397 vgnd vpwr scs8hd_decap_6
XFILLER_64_342 vgnd vpwr scs8hd_decap_12
X_66_ bottom_width_0_height_0__pin_44_lower bottom_width_0_height_0__pin_44_upper
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1_0_clk/X ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XFILLER_59_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_272 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ right_width_0_height_0__pin_4_ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_15_217 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_23_31 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ bottom_width_0_height_0__pin_29_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_2_154 vpwr vgnd scs8hd_fill_2
XFILLER_61_367 vgnd vpwr scs8hd_decap_4
XFILLER_9_33 vgnd vpwr scs8hd_fill_1
XFILLER_9_66 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_272 vgnd vpwr scs8hd_decap_3
XFILLER_50_3 vgnd vpwr scs8hd_decap_12
XFILLER_56_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_331 vgnd vpwr scs8hd_decap_12
XFILLER_52_301 vgnd vpwr scs8hd_decap_4
XFILLER_52_312 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
X_49_ _49_/HI _49_/LO vgnd vpwr scs8hd_conb_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_43_301 vpwr vgnd scs8hd_fill_2
XFILLER_28_320 vpwr vgnd scs8hd_fill_2
XFILLER_18_53 vpwr vgnd scs8hd_fill_2
XPHY_554 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_543 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_532 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_521 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_510 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_253 vpwr vgnd scs8hd_fill_2
XFILLER_7_268 vpwr vgnd scs8hd_fill_2
XFILLER_11_297 vpwr vgnd scs8hd_fill_2
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_301 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_40_337 vgnd vpwr scs8hd_decap_12
XFILLER_25_367 vgnd vpwr scs8hd_decap_12
XFILLER_20_76 vpwr vgnd scs8hd_fill_2
XFILLER_20_32 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_62 vgnd vpwr scs8hd_decap_12
XFILLER_45_51 vgnd vpwr scs8hd_decap_8
XFILLER_16_356 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XPHY_395 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_384 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_373 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_362 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_351 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_337 vpwr vgnd scs8hd_fill_2
XPHY_340 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_89 vgnd vpwr scs8hd_fill_1
XFILLER_39_404 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_245 vgnd vpwr scs8hd_decap_12
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_17_109 vgnd vpwr scs8hd_fill_1
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_21_392 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _35_/HI vgnd vpwr scs8hd_diode_2
XFILLER_13_348 vpwr vgnd scs8hd_fill_2
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_385 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_215 vgnd vpwr scs8hd_decap_12
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_64 vgnd vpwr scs8hd_fill_1
XFILLER_13_123 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_5_355 vpwr vgnd scs8hd_fill_2
XFILLER_9_127 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_36_215 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_27_259 vgnd vpwr scs8hd_decap_4
XFILLER_27_237 vgnd vpwr scs8hd_fill_1
XFILLER_50_295 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XFILLER_2_369 vpwr vgnd scs8hd_fill_2
XFILLER_58_395 vpwr vgnd scs8hd_fill_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_226 vpwr vgnd scs8hd_fill_2
XFILLER_18_215 vpwr vgnd scs8hd_fill_2
XFILLER_53_62 vgnd vpwr scs8hd_decap_12
XFILLER_53_51 vgnd vpwr scs8hd_decap_8
XFILLER_41_273 vgnd vpwr scs8hd_decap_3
XFILLER_5_174 vgnd vpwr scs8hd_decap_3
XFILLER_49_362 vpwr vgnd scs8hd_fill_2
XFILLER_64_354 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
X_65_ bottom_width_0_height_0__pin_43_lower bottom_width_0_height_0__pin_43_upper
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_32_262 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_159 vgnd vpwr scs8hd_decap_12
XFILLER_55_343 vgnd vpwr scs8hd_decap_4
XFILLER_55_310 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_23_240 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_2_111 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ bottom_width_0_height_0__pin_28_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_64_94 vgnd vpwr scs8hd_decap_12
XFILLER_46_398 vgnd vpwr scs8hd_decap_8
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_43_3 vgnd vpwr scs8hd_decap_12
XFILLER_56_129 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_376 vpwr vgnd scs8hd_fill_2
XFILLER_37_343 vgnd vpwr scs8hd_decap_3
X_48_ _48_/HI _48_/LO vgnd vpwr scs8hd_conb_1
XFILLER_52_346 vpwr vgnd scs8hd_fill_2
XFILLER_52_324 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_500 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_55_184 vgnd vpwr scs8hd_decap_12
XFILLER_28_398 vgnd vpwr scs8hd_decap_8
XFILLER_18_65 vpwr vgnd scs8hd_fill_2
XFILLER_18_43 vgnd vpwr scs8hd_fill_1
XFILLER_18_32 vgnd vpwr scs8hd_decap_4
XPHY_555 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_544 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_533 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_522 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_511 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_214 vgnd vpwr scs8hd_fill_1
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
XFILLER_11_221 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
XFILLER_19_332 vpwr vgnd scs8hd_fill_2
XFILLER_61_110 vgnd vpwr scs8hd_decap_12
XFILLER_34_379 vgnd vpwr scs8hd_decap_12
XFILLER_34_346 vgnd vpwr scs8hd_decap_8
XFILLER_34_335 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_52_154 vgnd vpwr scs8hd_decap_12
XFILLER_40_349 vgnd vpwr scs8hd_decap_8
XFILLER_33_390 vgnd vpwr scs8hd_decap_12
XFILLER_25_379 vgnd vpwr scs8hd_decap_12
XFILLER_20_88 vgnd vpwr scs8hd_decap_4
XFILLER_4_206 vpwr vgnd scs8hd_fill_2
XFILLER_45_74 vgnd vpwr scs8hd_decap_12
XFILLER_43_110 vgnd vpwr scs8hd_decap_12
XPHY_352 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_341 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_330 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_28_162 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_313 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_61_62 vgnd vpwr scs8hd_decap_12
XFILLER_61_51 vgnd vpwr scs8hd_decap_8
XPHY_396 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_385 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_374 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_363 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_162 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_257 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_316 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_99 vpwr vgnd scs8hd_fill_2
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ bottom_width_0_height_0__pin_18_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_48_202 vgnd vpwr scs8hd_decap_12
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
XFILLER_16_154 vgnd vpwr scs8hd_decap_12
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_257 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_227 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_157 vgnd vpwr scs8hd_decap_12
XFILLER_22_146 vgnd vpwr scs8hd_decap_6
XFILLER_10_319 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_290 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_8
XFILLER_53_260 vgnd vpwr scs8hd_decap_12
XFILLER_26_43 vpwr vgnd scs8hd_fill_2
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_5_301 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_208 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_205 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_35_293 vgnd vpwr scs8hd_decap_12
XFILLER_35_282 vpwr vgnd scs8hd_fill_2
XFILLER_10_116 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ right_width_0_height_0__pin_1_ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_56 vgnd vpwr scs8hd_decap_6
XFILLER_2_337 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_18_205 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_5_131 vpwr vgnd scs8hd_fill_2
XFILLER_5_197 vpwr vgnd scs8hd_fill_2
XFILLER_64_311 vgnd vpwr scs8hd_decap_12
XFILLER_49_341 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_392 vgnd vpwr scs8hd_decap_12
X_64_ bottom_width_0_height_0__pin_42_lower bottom_width_0_height_0__pin_42_upper
+ vgnd vpwr scs8hd_buf_2
XFILLER_64_366 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_285 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _61_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ top_width_0_height_0__pin_33_ vgnd vpwr scs8hd_diode_2
XFILLER_11_403 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_145 vgnd vpwr scs8hd_fill_1
XFILLER_46_333 vgnd vpwr scs8hd_decap_3
XFILLER_61_347 vpwr vgnd scs8hd_fill_2
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_57 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XFILLER_49_171 vgnd vpwr scs8hd_decap_12
X_47_ _47_/HI _47_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_52_369 vpwr vgnd scs8hd_fill_2
XFILLER_20_211 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_534 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_523 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_512 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_501 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_55_196 vgnd vpwr scs8hd_decap_12
XFILLER_43_358 vpwr vgnd scs8hd_fill_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_377 vgnd vpwr scs8hd_decap_12
XFILLER_18_88 vpwr vgnd scs8hd_fill_2
XPHY_556 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_545 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_380 vpwr vgnd scs8hd_fill_2
XFILLER_7_226 vgnd vpwr scs8hd_decap_4
XFILLER_11_233 vgnd vpwr scs8hd_fill_1
XFILLER_59_62 vgnd vpwr scs8hd_decap_12
XFILLER_59_51 vgnd vpwr scs8hd_decap_8
XFILLER_46_141 vgnd vpwr scs8hd_decap_12
XFILLER_34_325 vgnd vpwr scs8hd_decap_4
XFILLER_19_355 vgnd vpwr scs8hd_decap_4
XFILLER_42_391 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_281 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_57_406 vgnd vpwr scs8hd_fill_1
XFILLER_29_119 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_166 vgnd vpwr scs8hd_decap_12
XFILLER_40_317 vpwr vgnd scs8hd_fill_2
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_25_347 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0_0_clk/X ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_402 vgnd vpwr scs8hd_fill_1
XFILLER_48_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_28_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_45_86 vgnd vpwr scs8hd_decap_12
XPHY_386 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_375 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_364 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_353 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_306 vgnd vpwr scs8hd_decap_12
XPHY_342 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_331 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_28_185 vpwr vgnd scs8hd_fill_2
XPHY_320 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_16_325 vgnd vpwr scs8hd_decap_8
XFILLER_61_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_397 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_36 vgnd vpwr scs8hd_decap_12
XFILLER_6_58 vgnd vpwr scs8hd_decap_4
XFILLER_6_69 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_262 vpwr vgnd scs8hd_fill_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_22_306 vgnd vpwr scs8hd_fill_1
XFILLER_22_328 vpwr vgnd scs8hd_fill_2
XFILLER_57_269 vgnd vpwr scs8hd_decap_12
XFILLER_13_306 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ bottom_width_0_height_0__pin_17_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_166 vgnd vpwr scs8hd_decap_12
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_361 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_398 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _48_/HI
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_49_lower vgnd vpwr scs8hd_mux2_1
XFILLER_54_239 vgnd vpwr scs8hd_decap_12
XFILLER_47_280 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_169 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_280 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ bottom_width_0_height_0__pin_29_ vgnd vpwr scs8hd_diode_2
XFILLER_53_272 vgnd vpwr scs8hd_decap_12
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_103 vpwr vgnd scs8hd_fill_2
XFILLER_13_158 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
X_80_ right_width_0_height_0__pin_41_lower right_width_0_height_0__pin_41_upper vgnd
+ vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1_0_clk/X ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_26 vpwr vgnd scs8hd_fill_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_44_272 vgnd vpwr scs8hd_fill_1
XFILLER_12_191 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_390 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_23_401 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_316 vpwr vgnd scs8hd_fill_2
XFILLER_58_320 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_53_86 vgnd vpwr scs8hd_decap_12
XFILLER_41_297 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_64_323 vgnd vpwr scs8hd_decap_12
XFILLER_49_386 vpwr vgnd scs8hd_fill_2
X_63_ _63_/HI _63_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_378 vpwr vgnd scs8hd_fill_2
XFILLER_55_367 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_23_286 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_46_312 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XFILLER_64_63 vgnd vpwr scs8hd_decap_12
XFILLER_46_389 vgnd vpwr scs8hd_decap_8
XFILLER_9_36 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_52_337 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_356 vgnd vpwr scs8hd_decap_4
XFILLER_37_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
X_46_ _46_/HI _46_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_245 vgnd vpwr scs8hd_decap_12
XFILLER_20_223 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _47_/HI ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
XFILLER_28_356 vgnd vpwr scs8hd_decap_12
XPHY_557 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_546 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_535 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_524 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_513 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_502 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_392 vgnd vpwr scs8hd_decap_12
XFILLER_43_337 vpwr vgnd scs8hd_fill_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_28_389 vgnd vpwr scs8hd_decap_8
XFILLER_50_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_245 vgnd vpwr scs8hd_decap_8
XFILLER_59_74 vgnd vpwr scs8hd_decap_12
XFILLER_61_123 vgnd vpwr scs8hd_decap_12
XFILLER_19_389 vgnd vpwr scs8hd_decap_12
XFILLER_19_367 vgnd vpwr scs8hd_decap_3
XFILLER_19_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_52_178 vgnd vpwr scs8hd_decap_12
XFILLER_1_81 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _56_/HI vgnd vpwr scs8hd_diode_2
XFILLER_20_68 vgnd vpwr scs8hd_decap_6
XFILLER_20_46 vgnd vpwr scs8hd_decap_12
XFILLER_43_123 vgnd vpwr scs8hd_decap_12
XFILLER_29_99 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_61_86 vgnd vpwr scs8hd_decap_12
XFILLER_45_98 vgnd vpwr scs8hd_decap_12
XPHY_398 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_387 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_376 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_365 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_354 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_343 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_318 vgnd vpwr scs8hd_decap_12
XPHY_332 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_321 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_310 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_230 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ bottom_width_0_height_0__pin_23_ vgnd vpwr scs8hd_diode_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_6_48 vgnd vpwr scs8hd_fill_1
XFILLER_3_285 vpwr vgnd scs8hd_fill_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XFILLER_15_381 vgnd vpwr scs8hd_decap_12
XFILLER_30_340 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_362 vpwr vgnd scs8hd_fill_2
XFILLER_21_340 vpwr vgnd scs8hd_fill_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ bottom_width_0_height_0__pin_16_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_48_215 vgnd vpwr scs8hd_decap_12
XFILLER_0_299 vgnd vpwr scs8hd_decap_4
XFILLER_0_244 vpwr vgnd scs8hd_fill_2
XFILLER_16_178 vgnd vpwr scs8hd_decap_4
XFILLER_16_145 vgnd vpwr scs8hd_decap_8
XFILLER_16_112 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_159 vgnd vpwr scs8hd_fill_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_333 vgnd vpwr scs8hd_decap_3
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_373 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_62_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_115 vgnd vpwr scs8hd_decap_6
XFILLER_7_91 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_284 vgnd vpwr scs8hd_decap_3
XFILLER_26_67 vpwr vgnd scs8hd_fill_2
XFILLER_26_56 vgnd vpwr scs8hd_decap_8
XFILLER_13_115 vgnd vpwr scs8hd_fill_1
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_21_192 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_137 vpwr vgnd scs8hd_fill_2
XFILLER_13_148 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _63_/HI ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_229 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_328 vpwr vgnd scs8hd_fill_2
XFILLER_58_398 vgnd vpwr scs8hd_decap_8
XFILLER_58_332 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_295 vgnd vpwr scs8hd_decap_12
XFILLER_26_240 vpwr vgnd scs8hd_fill_2
XFILLER_53_98 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_5_111 vgnd vpwr scs8hd_decap_3
XFILLER_64_335 vgnd vpwr scs8hd_decap_6
XFILLER_49_398 vpwr vgnd scs8hd_fill_2
X_62_ _62_/HI _62_/LO vgnd vpwr scs8hd_conb_1
XFILLER_17_240 vpwr vgnd scs8hd_fill_2
XFILLER_32_210 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_81 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_23_298 vgnd vpwr scs8hd_decap_6
XFILLER_23_68 vpwr vgnd scs8hd_fill_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_48_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ right_width_0_height_0__pin_6_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_2_169 vpwr vgnd scs8hd_fill_2
XFILLER_2_158 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ccff_tail vgnd vpwr scs8hd_diode_2
XFILLER_46_346 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _57_/HI
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_36_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_75 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_276 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_49_184 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_64_187 vgnd vpwr scs8hd_decap_12
XFILLER_52_305 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
X_45_ _45_/HI _45_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_257 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_55_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_28_368 vgnd vpwr scs8hd_decap_4
XFILLER_28_335 vgnd vpwr scs8hd_fill_1
XFILLER_18_57 vgnd vpwr scs8hd_decap_4
XPHY_558 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_547 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_536 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_525 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_514 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_503 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XFILLER_11_257 vpwr vgnd scs8hd_fill_2
XFILLER_50_44 vgnd vpwr scs8hd_decap_12
XFILLER_7_217 vgnd vpwr scs8hd_fill_1
XFILLER_59_86 vgnd vpwr scs8hd_decap_12
XFILLER_61_135 vgnd vpwr scs8hd_decap_12
XFILLER_46_154 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_42_371 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _55_/HI vgnd vpwr scs8hd_diode_2
XFILLER_6_261 vgnd vpwr scs8hd_decap_8
XFILLER_6_294 vpwr vgnd scs8hd_fill_2
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_25_316 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_190 vgnd vpwr scs8hd_decap_12
XFILLER_20_58 vgnd vpwr scs8hd_decap_4
XFILLER_20_36 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_404 vgnd vpwr scs8hd_decap_3
XFILLER_43_135 vgnd vpwr scs8hd_decap_12
XFILLER_28_154 vgnd vpwr scs8hd_decap_8
XPHY_300 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_61_98 vgnd vpwr scs8hd_decap_12
XPHY_399 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_388 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_377 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_366 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_355 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_344 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_333 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_322 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_311 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_110 vpwr vgnd scs8hd_fill_2
XFILLER_3_297 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_42_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_15_371 vpwr vgnd scs8hd_fill_2
XFILLER_15_393 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_30_396 vgnd vpwr scs8hd_fill_1
XFILLER_30_374 vpwr vgnd scs8hd_fill_2
XANTENNA_clkbuf_0_clk_A clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_25_135 vgnd vpwr scs8hd_decap_12
XFILLER_25_102 vpwr vgnd scs8hd_fill_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ bottom_width_0_height_0__pin_26_ vgnd vpwr scs8hd_diode_2
XFILLER_63_208 vgnd vpwr scs8hd_decap_12
XFILLER_56_32 vgnd vpwr scs8hd_decap_12
XFILLER_48_227 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_385 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_62_263 vgnd vpwr scs8hd_decap_12
XFILLER_30_182 vgnd vpwr scs8hd_decap_4
XFILLER_30_160 vgnd vpwr scs8hd_fill_1
XFILLER_30_193 vpwr vgnd scs8hd_fill_2
XFILLER_7_81 vpwr vgnd scs8hd_fill_2
XFILLER_45_208 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_12
XFILLER_5_315 vpwr vgnd scs8hd_fill_2
XFILLER_5_359 vpwr vgnd scs8hd_fill_2
XFILLER_36_219 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_44_285 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_131 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_35_241 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XFILLER_58_300 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_26_274 vgnd vpwr scs8hd_fill_1
XFILLER_26_263 vgnd vpwr scs8hd_decap_3
XFILLER_49_333 vpwr vgnd scs8hd_fill_2
X_61_ _61_/HI _61_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_255 vgnd vpwr scs8hd_decap_4
XFILLER_32_244 vpwr vgnd scs8hd_fill_2
XFILLER_20_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_55_358 vpwr vgnd scs8hd_fill_2
XFILLER_55_347 vgnd vpwr scs8hd_fill_1
XFILLER_55_314 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_71 vgnd vpwr scs8hd_fill_1
XFILLER_4_93 vpwr vgnd scs8hd_fill_2
XFILLER_63_391 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_141 vgnd vpwr scs8hd_decap_12
XFILLER_48_44 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ right_width_0_height_0__pin_5_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_2_148 vpwr vgnd scs8hd_fill_2
XFILLER_2_115 vpwr vgnd scs8hd_fill_2
XFILLER_64_87 vgnd vpwr scs8hd_decap_6
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
XFILLER_61_306 vgnd vpwr scs8hd_decap_12
XFILLER_46_369 vgnd vpwr scs8hd_fill_1
XFILLER_46_325 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1_0_clk/X ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_27 vgnd vpwr scs8hd_decap_6
XFILLER_14_233 vgnd vpwr scs8hd_decap_6
XFILLER_14_288 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_49_196 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_170 vgnd vpwr scs8hd_decap_3
X_44_ _44_/HI _44_/LO vgnd vpwr scs8hd_conb_1
XFILLER_64_199 vgnd vpwr scs8hd_decap_12
XFILLER_60_383 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_269 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_43_306 vgnd vpwr scs8hd_decap_4
XFILLER_18_69 vpwr vgnd scs8hd_fill_2
XFILLER_18_36 vgnd vpwr scs8hd_fill_1
XPHY_559 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_548 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_537 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_526 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_515 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_504 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_11_203 vpwr vgnd scs8hd_fill_2
XFILLER_11_225 vgnd vpwr scs8hd_decap_8
XFILLER_11_236 vpwr vgnd scs8hd_fill_2
XFILLER_50_56 vgnd vpwr scs8hd_decap_12
XFILLER_59_98 vgnd vpwr scs8hd_decap_12
XFILLER_19_336 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _45_/HI vgnd vpwr scs8hd_diode_2
XFILLER_61_147 vgnd vpwr scs8hd_decap_12
XFILLER_46_166 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_306 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_361 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_68 vgnd vpwr scs8hd_fill_1
XFILLER_43_147 vgnd vpwr scs8hd_decap_12
XPHY_334 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_323 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_312 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_301 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_16_317 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_389 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_378 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_367 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_356 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_345 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_70 vgnd vpwr scs8hd_decap_4
XFILLER_19_166 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_147 vgnd vpwr scs8hd_decap_12
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1_0_clk/X ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XFILLER_21_353 vpwr vgnd scs8hd_fill_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XFILLER_56_44 vgnd vpwr scs8hd_decap_12
XFILLER_48_239 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_120 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_302 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_91 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_clkbuf_1_0_0_clk_A clkbuf_0_clk/X vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ bottom_width_0_height_0__pin_20_ vgnd vpwr scs8hd_diode_2
XFILLER_38_250 vgnd vpwr scs8hd_decap_12
XFILLER_53_297 vpwr vgnd scs8hd_fill_2
XFILLER_53_220 vgnd vpwr scs8hd_decap_12
XFILLER_41_404 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_68 vgnd vpwr scs8hd_decap_12
XFILLER_5_338 vpwr vgnd scs8hd_fill_2
XFILLER_44_264 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ bottom_width_0_height_0__pin_31_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_or2_1
XFILLER_8_154 vpwr vgnd scs8hd_fill_2
XFILLER_12_183 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_165 vgnd vpwr scs8hd_decap_8
XFILLER_27_209 vgnd vpwr scs8hd_decap_4
XFILLER_50_267 vpwr vgnd scs8hd_fill_2
XFILLER_50_245 vgnd vpwr scs8hd_fill_1
XFILLER_35_286 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XFILLER_58_312 vgnd vpwr scs8hd_fill_1
XFILLER_58_356 vgnd vpwr scs8hd_decap_6
XFILLER_41_278 vpwr vgnd scs8hd_fill_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_5_135 vpwr vgnd scs8hd_fill_2
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_64_304 vgnd vpwr scs8hd_decap_6
XFILLER_49_345 vgnd vpwr scs8hd_fill_1
XFILLER_49_301 vpwr vgnd scs8hd_fill_2
X_60_ _60_/HI _60_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_330 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_297 vpwr vgnd scs8hd_fill_2
XFILLER_17_264 vgnd vpwr scs8hd_decap_12
XFILLER_17_220 vpwr vgnd scs8hd_fill_2
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_289 vpwr vgnd scs8hd_fill_2
XFILLER_32_267 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_326 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_278 vpwr vgnd scs8hd_fill_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ right_width_0_height_0__pin_4_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_48_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
XFILLER_61_318 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_46_359 vpwr vgnd scs8hd_fill_2
XFILLER_0_19 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_70 vpwr vgnd scs8hd_fill_2
XFILLER_13_92 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_64_156 vgnd vpwr scs8hd_decap_12
XFILLER_37_348 vpwr vgnd scs8hd_fill_2
X_43_ _43_/HI _43_/LO vgnd vpwr scs8hd_conb_1
XFILLER_60_395 vpwr vgnd scs8hd_fill_2
XFILLER_45_392 vgnd vpwr scs8hd_decap_12
XFILLER_20_215 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_9_271 vpwr vgnd scs8hd_fill_2
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XPHY_516 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_505 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_55_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XPHY_549 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_538 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_527 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_362 vpwr vgnd scs8hd_fill_2
XFILLER_50_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_359 vgnd vpwr scs8hd_fill_1
XFILLER_19_315 vpwr vgnd scs8hd_fill_2
XFILLER_61_159 vgnd vpwr scs8hd_decap_12
XFILLER_46_178 vgnd vpwr scs8hd_decap_12
XFILLER_42_340 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_230 vpwr vgnd scs8hd_fill_2
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_43_159 vgnd vpwr scs8hd_decap_12
XPHY_368 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_357 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_346 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_335 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_324 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_28_189 vpwr vgnd scs8hd_fill_2
XPHY_313 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_302 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_379 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_4
XFILLER_59_281 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_178 vgnd vpwr scs8hd_decap_3
XFILLER_19_123 vgnd vpwr scs8hd_decap_3
XFILLER_30_398 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_159 vgnd vpwr scs8hd_fill_1
XFILLER_21_321 vgnd vpwr scs8hd_decap_4
XFILLER_21_310 vgnd vpwr scs8hd_decap_4
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_56_251 vgnd vpwr scs8hd_decap_12
XFILLER_56_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _40_/HI vgnd vpwr scs8hd_diode_2
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_325 vgnd vpwr scs8hd_decap_8
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_70 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_398 vgnd vpwr scs8hd_decap_8
XFILLER_47_240 vpwr vgnd scs8hd_fill_2
XFILLER_62_276 vgnd vpwr scs8hd_decap_12
XFILLER_47_284 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_7_391 vgnd vpwr scs8hd_decap_12
XFILLER_53_232 vgnd vpwr scs8hd_decap_12
XFILLER_38_262 vgnd vpwr scs8hd_decap_12
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_107 vgnd vpwr scs8hd_decap_8
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_19 vgnd vpwr scs8hd_fill_1
XFILLER_29_251 vgnd vpwr scs8hd_fill_1
XFILLER_17_402 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_177 vpwr vgnd scs8hd_fill_2
XFILLER_12_151 vpwr vgnd scs8hd_fill_2
XFILLER_12_162 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _38_/HI
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_4_361 vpwr vgnd scs8hd_fill_2
XFILLER_50_202 vgnd vpwr scs8hd_decap_12
XFILLER_35_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_210 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_158 vpwr vgnd scs8hd_fill_2
XFILLER_57_390 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_224 vgnd vpwr scs8hd_decap_8
XFILLER_32_213 vgnd vpwr scs8hd_fill_1
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XFILLER_40_290 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_51 vgnd vpwr scs8hd_decap_3
XFILLER_23_213 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _37_/HI
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_42_lower vgnd vpwr scs8hd_mux2_1
XFILLER_23_268 vpwr vgnd scs8hd_fill_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_154 vgnd vpwr scs8hd_decap_12
XFILLER_48_68 vgnd vpwr scs8hd_decap_12
XFILLER_46_316 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_64_56 vgnd vpwr scs8hd_decap_6
XFILLER_54_360 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_14_202 vgnd vpwr scs8hd_decap_12
XFILLER_14_224 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_82 vpwr vgnd scs8hd_fill_2
XFILLER_49_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_64_168 vgnd vpwr scs8hd_decap_12
XFILLER_52_308 vpwr vgnd scs8hd_fill_2
X_42_ _42_/HI _42_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_290 vgnd vpwr scs8hd_decap_12
XFILLER_9_294 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_327 vgnd vpwr scs8hd_decap_8
XFILLER_28_316 vpwr vgnd scs8hd_fill_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_539 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_528 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_517 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_506 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_55_135 vgnd vpwr scs8hd_decap_12
XFILLER_51_341 vpwr vgnd scs8hd_fill_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_404 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_190 vgnd vpwr scs8hd_decap_12
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_30 vpwr vgnd scs8hd_fill_2
XFILLER_52_105 vgnd vpwr scs8hd_decap_12
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
XFILLER_1_85 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_51_171 vgnd vpwr scs8hd_decap_12
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XPHY_369 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_358 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_347 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_336 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_325 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_314 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_303 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_341 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_234 vpwr vgnd scs8hd_fill_2
XFILLER_3_289 vpwr vgnd scs8hd_fill_2
XFILLER_10_83 vgnd vpwr scs8hd_decap_8
XFILLER_59_293 vgnd vpwr scs8hd_decap_12
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_135 vpwr vgnd scs8hd_fill_2
XFILLER_19_92 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_30_344 vgnd vpwr scs8hd_decap_4
XFILLER_30_322 vgnd vpwr scs8hd_decap_12
XFILLER_30_300 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ bottom_width_0_height_0__pin_17_ vgnd vpwr scs8hd_diode_2
XFILLER_57_208 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_33_193 vpwr vgnd scs8hd_fill_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XFILLER_21_388 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_56_263 vgnd vpwr scs8hd_decap_12
XFILLER_56_68 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_337 vgnd vpwr scs8hd_decap_12
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_311 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_208 vgnd vpwr scs8hd_decap_12
XFILLER_62_288 vgnd vpwr scs8hd_decap_12
XFILLER_50_406 vgnd vpwr scs8hd_fill_1
Xclkbuf_0_clk clk clkbuf_0_clk/X vgnd vpwr scs8hd_clkbuf_16
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_30_152 vgnd vpwr scs8hd_fill_1
XFILLER_38_296 vpwr vgnd scs8hd_fill_2
XFILLER_38_274 vgnd vpwr scs8hd_fill_1
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_406 vgnd vpwr scs8hd_fill_1
XFILLER_29_274 vpwr vgnd scs8hd_fill_2
XFILLER_8_145 vpwr vgnd scs8hd_fill_2
XFILLER_4_340 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_35_233 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1_0_clk/X ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_406 vgnd vpwr scs8hd_fill_1
XFILLER_5_104 vgnd vpwr scs8hd_decap_3
XFILLER_49_358 vpwr vgnd scs8hd_fill_2
XFILLER_49_325 vgnd vpwr scs8hd_decap_8
XFILLER_32_236 vgnd vpwr scs8hd_decap_6
XFILLER_55_306 vpwr vgnd scs8hd_fill_2
XFILLER_4_63 vpwr vgnd scs8hd_fill_2
XFILLER_4_85 vgnd vpwr scs8hd_decap_4
XFILLER_23_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_291 vgnd vpwr scs8hd_decap_12
XFILLER_23_258 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_58_166 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_306 vgnd vpwr scs8hd_fill_1
X_41_ _41_/HI _41_/LO vgnd vpwr scs8hd_conb_1
XFILLER_64_125 vgnd vpwr scs8hd_decap_12
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_240 vpwr vgnd scs8hd_fill_2
XFILLER_55_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ right_width_0_height_0__pin_11_ vgnd vpwr scs8hd_diode_2
XFILLER_18_39 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XPHY_529 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_518 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_507 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_331 vgnd vpwr scs8hd_decap_4
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_217 vpwr vgnd scs8hd_fill_2
XFILLER_50_15 vgnd vpwr scs8hd_decap_12
XFILLER_34_309 vgnd vpwr scs8hd_fill_1
XANTENNA__64__A bottom_width_0_height_0__pin_42_lower vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
XFILLER_24_60 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ bottom_width_0_height_0__pin_19_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_or2_1
XFILLER_6_210 vgnd vpwr scs8hd_decap_4
XFILLER_6_276 vgnd vpwr scs8hd_decap_3
XFILLER_6_298 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_294 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1_0_clk/X ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_52_117 vgnd vpwr scs8hd_decap_12
XFILLER_18_361 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XFILLER_45_59 vpwr vgnd scs8hd_fill_2
XFILLER_45_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_359 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_348 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_337 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_326 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_315 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_304 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_353 vpwr vgnd scs8hd_fill_2
XFILLER_3_213 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
XFILLER_30_312 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_378 vgnd vpwr scs8hd_decap_12
XFILLER_30_367 vpwr vgnd scs8hd_fill_2
XFILLER_30_334 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_106 vgnd vpwr scs8hd_decap_12
XFILLER_21_367 vpwr vgnd scs8hd_fill_2
XFILLER_21_301 vpwr vgnd scs8hd_fill_2
XFILLER_15_29 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XFILLER_0_238 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_decap_3
XFILLER_24_172 vgnd vpwr scs8hd_decap_3
XFILLER_24_150 vgnd vpwr scs8hd_decap_3
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_194 vgnd vpwr scs8hd_decap_3
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_349 vgnd vpwr scs8hd_decap_12
XFILLER_12_323 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_21_50 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_297 vpwr vgnd scs8hd_fill_2
XFILLER_47_264 vpwr vgnd scs8hd_fill_2
XFILLER_47_220 vgnd vpwr scs8hd_decap_12
XFILLER_35_404 vgnd vpwr scs8hd_decap_3
XFILLER_46_80 vgnd vpwr scs8hd_decap_12
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_161 vgnd vpwr scs8hd_decap_12
XFILLER_30_186 vgnd vpwr scs8hd_fill_1
XFILLER_7_85 vgnd vpwr scs8hd_decap_4
XFILLER_53_289 vgnd vpwr scs8hd_decap_6
XFILLER_53_245 vgnd vpwr scs8hd_decap_12
XFILLER_38_286 vgnd vpwr scs8hd_fill_1
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_5_319 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA__72__A bottom_width_0_height_0__pin_50_ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_4_330 vpwr vgnd scs8hd_fill_2
XFILLER_4_374 vpwr vgnd scs8hd_fill_2
XFILLER_4_396 vgnd vpwr scs8hd_fill_1
XFILLER_50_215 vgnd vpwr scs8hd_decap_12
XFILLER_35_212 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ bottom_width_0_height_0__pin_50_ vgnd vpwr scs8hd_diode_2
XFILLER_58_315 vgnd vpwr scs8hd_decap_3
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_53_59 vpwr vgnd scs8hd_fill_2
XFILLER_53_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_116 vgnd vpwr scs8hd_decap_4
XFILLER_5_127 vpwr vgnd scs8hd_fill_2
XFILLER_49_348 vgnd vpwr scs8hd_fill_1
XANTENNA__67__A bottom_width_0_height_0__pin_45_lower vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_259 vgnd vpwr scs8hd_fill_1
XFILLER_4_171 vgnd vpwr scs8hd_decap_3
XFILLER_4_193 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_381 vgnd vpwr scs8hd_decap_12
XFILLER_23_204 vgnd vpwr scs8hd_decap_3
XFILLER_48_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_119 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_58_178 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_392 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_62 vgnd vpwr scs8hd_decap_4
XFILLER_13_95 vgnd vpwr scs8hd_decap_8
XFILLER_49_123 vgnd vpwr scs8hd_decap_12
X_40_ _40_/HI _40_/LO vgnd vpwr scs8hd_conb_1
XFILLER_64_137 vgnd vpwr scs8hd_decap_12
XFILLER_54_80 vgnd vpwr scs8hd_decap_12
XFILLER_45_362 vpwr vgnd scs8hd_fill_2
XFILLER_45_340 vpwr vgnd scs8hd_fill_2
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
XFILLER_60_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_55_159 vgnd vpwr scs8hd_decap_12
XPHY_519 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_508 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_376 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_384 vpwr vgnd scs8hd_fill_2
XFILLER_11_207 vgnd vpwr scs8hd_decap_4
XFILLER_50_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_7 vpwr vgnd scs8hd_fill_2
XFILLER_42_321 vpwr vgnd scs8hd_fill_2
XFILLER_27_362 vgnd vpwr scs8hd_decap_4
XANTENNA__80__A right_width_0_height_0__pin_41_lower vgnd vpwr scs8hd_diode_2
XFILLER_42_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_72 vgnd vpwr scs8hd_fill_1
XFILLER_6_222 vpwr vgnd scs8hd_fill_2
XFILLER_10_240 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ right_width_0_height_0__pin_14_ vgnd vpwr scs8hd_diode_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
XFILLER_52_129 vgnd vpwr scs8hd_decap_12
XFILLER_33_365 vgnd vpwr scs8hd_fill_1
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XFILLER_45_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_316 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_305 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_61_59 vpwr vgnd scs8hd_fill_2
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XFILLER_51_184 vgnd vpwr scs8hd_decap_12
XPHY_349 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_338 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_327 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_398 vgnd vpwr scs8hd_decap_8
XFILLER_24_365 vgnd vpwr scs8hd_decap_3
XFILLER_3_258 vpwr vgnd scs8hd_fill_2
XANTENNA__75__A right_width_0_height_0__pin_36_lower vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_118 vgnd vpwr scs8hd_decap_4
XFILLER_33_184 vgnd vpwr scs8hd_decap_4
XFILLER_21_357 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_56_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_56_276 vgnd vpwr scs8hd_decap_12
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_335 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_202 vgnd vpwr scs8hd_decap_12
XFILLER_47_276 vpwr vgnd scs8hd_fill_2
XFILLER_47_232 vpwr vgnd scs8hd_fill_2
XFILLER_62_80 vgnd vpwr scs8hd_decap_12
XFILLER_30_154 vgnd vpwr scs8hd_decap_6
XPHY_4 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_257 vgnd vpwr scs8hd_fill_1
XFILLER_38_276 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_21_132 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _60_/HI
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_39_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_202 vgnd vpwr scs8hd_decap_12
XFILLER_29_287 vgnd vpwr scs8hd_decap_12
XFILLER_29_254 vgnd vpwr scs8hd_decap_12
XFILLER_29_243 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_16_84 vpwr vgnd scs8hd_fill_2
XFILLER_16_51 vpwr vgnd scs8hd_fill_2
XFILLER_12_154 vgnd vpwr scs8hd_decap_8
XFILLER_12_187 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_8_158 vgnd vpwr scs8hd_decap_4
XFILLER_50_227 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_27 vgnd vpwr scs8hd_decap_12
XFILLER_26_268 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_367 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _49_/HI
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_48_lower vgnd vpwr scs8hd_mux2_1
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
XFILLER_4_76 vgnd vpwr scs8hd_decap_3
XFILLER_63_330 vgnd vpwr scs8hd_decap_12
XFILLER_48_393 vgnd vpwr scs8hd_decap_4
XFILLER_16_290 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_48_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _43_/HI vgnd vpwr scs8hd_diode_2
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
XFILLER_54_352 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_282 vgnd vpwr scs8hd_decap_12
XFILLER_13_74 vpwr vgnd scs8hd_fill_2
XANTENNA__78__A right_width_0_height_0__pin_39_lower vgnd vpwr scs8hd_diode_2
XFILLER_1_142 vpwr vgnd scs8hd_fill_2
XFILLER_64_149 vgnd vpwr scs8hd_decap_6
XFILLER_49_135 vgnd vpwr scs8hd_decap_12
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_175 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_60_300 vgnd vpwr scs8hd_decap_12
XFILLER_55_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_220 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_63_171 vgnd vpwr scs8hd_decap_12
XFILLER_51_300 vpwr vgnd scs8hd_fill_2
XFILLER_48_190 vgnd vpwr scs8hd_decap_12
XFILLER_36_396 vgnd vpwr scs8hd_fill_1
XPHY_509 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_388 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_59_59 vpwr vgnd scs8hd_fill_2
XFILLER_59_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _57_/HI vgnd vpwr scs8hd_diode_2
XFILLER_46_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_319 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_42_344 vgnd vpwr scs8hd_fill_1
XFILLER_27_341 vpwr vgnd scs8hd_fill_2
XFILLER_24_40 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_24_84 vgnd vpwr scs8hd_decap_8
XFILLER_6_234 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_11 vgnd vpwr scs8hd_decap_8
XFILLER_60_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_105 vgnd vpwr scs8hd_decap_12
XFILLER_45_39 vgnd vpwr scs8hd_decap_12
XPHY_339 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_328 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_317 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_306 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_333 vgnd vpwr scs8hd_decap_3
XFILLER_24_311 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_61_27 vgnd vpwr scs8hd_decap_12
XFILLER_51_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_226 vpwr vgnd scs8hd_fill_2
XFILLER_62_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ right_width_0_height_0__pin_8_ vgnd vpwr scs8hd_diode_2
XFILLER_19_62 vpwr vgnd scs8hd_fill_2
XFILLER_15_300 vgnd vpwr scs8hd_decap_3
XFILLER_42_141 vgnd vpwr scs8hd_decap_12
XFILLER_27_193 vpwr vgnd scs8hd_fill_2
XFILLER_15_333 vpwr vgnd scs8hd_fill_2
XFILLER_15_377 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_53_406 vgnd vpwr scs8hd_fill_1
XFILLER_21_336 vpwr vgnd scs8hd_fill_2
XFILLER_21_314 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_0_218 vgnd vpwr scs8hd_fill_1
XFILLER_56_288 vgnd vpwr scs8hd_decap_12
XFILLER_56_27 vgnd vpwr scs8hd_decap_4
XFILLER_44_406 vgnd vpwr scs8hd_fill_1
XFILLER_29_403 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XPHY_103 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_74 vpwr vgnd scs8hd_fill_2
XFILLER_20_380 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1_0_clk/X ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XPHY_5 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_11_391 vgnd vpwr scs8hd_decap_12
XFILLER_26_406 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_29_299 vgnd vpwr scs8hd_decap_6
XFILLER_29_266 vgnd vpwr scs8hd_decap_6
XFILLER_29_233 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_406 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ right_width_0_height_0__pin_7_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_or2_1
XFILLER_16_74 vpwr vgnd scs8hd_fill_2
XFILLER_12_122 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_50_239 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_26_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_206 vgnd vpwr scs8hd_decap_4
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_25_280 vpwr vgnd scs8hd_fill_2
XFILLER_17_236 vpwr vgnd scs8hd_fill_2
XFILLER_40_272 vgnd vpwr scs8hd_decap_3
XFILLER_40_250 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_342 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_16_280 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
XFILLER_22_294 vgnd vpwr scs8hd_decap_12
XFILLER_22_250 vpwr vgnd scs8hd_fill_2
XFILLER_13_86 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_106 vgnd vpwr scs8hd_decap_12
XFILLER_49_147 vgnd vpwr scs8hd_decap_12
XFILLER_60_356 vgnd vpwr scs8hd_decap_6
XFILLER_60_312 vgnd vpwr scs8hd_decap_12
XFILLER_54_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_298 vpwr vgnd scs8hd_fill_2
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_51_345 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_331 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ bottom_width_0_height_0__pin_50_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_42_367 vpwr vgnd scs8hd_fill_2
XFILLER_27_375 vgnd vpwr scs8hd_decap_12
XFILLER_6_202 vpwr vgnd scs8hd_fill_2
XFILLER_6_257 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_89 vgnd vpwr scs8hd_decap_4
XFILLER_33_367 vpwr vgnd scs8hd_fill_2
XFILLER_28_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_61_39 vgnd vpwr scs8hd_decap_12
XPHY_329 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_318 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_307 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_389 vgnd vpwr scs8hd_decap_8
XFILLER_24_345 vgnd vpwr scs8hd_decap_4
XFILLER_59_220 vgnd vpwr scs8hd_decap_12
XFILLER_47_404 vgnd vpwr scs8hd_decap_3
XFILLER_3_238 vgnd vpwr scs8hd_decap_4
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_139 vpwr vgnd scs8hd_fill_2
XFILLER_19_96 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XFILLER_30_359 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_356 vgnd vpwr scs8hd_decap_8
XFILLER_15_367 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_293 vpwr vgnd scs8hd_fill_2
XFILLER_2_271 vpwr vgnd scs8hd_fill_2
XFILLER_33_197 vgnd vpwr scs8hd_decap_4
XFILLER_18_161 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _52_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_126 vgnd vpwr scs8hd_decap_3
XPHY_115 vgnd vpwr scs8hd_decap_3
XPHY_104 vgnd vpwr scs8hd_decap_3
XFILLER_24_142 vgnd vpwr scs8hd_decap_8
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_337 vgnd vpwr scs8hd_decap_12
XFILLER_62_215 vgnd vpwr scs8hd_decap_12
XFILLER_30_112 vgnd vpwr scs8hd_decap_12
XPHY_6 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_62_93 vgnd vpwr scs8hd_decap_12
XFILLER_30_189 vpwr vgnd scs8hd_fill_2
XFILLER_7_44 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_61_281 vgnd vpwr scs8hd_decap_12
XFILLER_21_167 vgnd vpwr scs8hd_decap_12
XFILLER_29_245 vgnd vpwr scs8hd_decap_6
XFILLER_44_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_149 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_311 vpwr vgnd scs8hd_fill_2
XFILLER_4_344 vpwr vgnd scs8hd_fill_2
XFILLER_35_237 vgnd vpwr scs8hd_decap_4
XFILLER_35_248 vgnd vpwr scs8hd_decap_4
XPHY_490 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_215 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ bottom_width_0_height_0__pin_26_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_1_358 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_43_62 vgnd vpwr scs8hd_decap_12
XFILLER_43_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_74 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_403 vgnd vpwr scs8hd_decap_4
XFILLER_4_67 vpwr vgnd scs8hd_fill_2
XFILLER_4_89 vgnd vpwr scs8hd_fill_1
XFILLER_4_163 vpwr vgnd scs8hd_fill_2
XFILLER_63_354 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_362 vpwr vgnd scs8hd_fill_2
XFILLER_54_398 vgnd vpwr scs8hd_decap_8
XFILLER_22_240 vgnd vpwr scs8hd_decap_8
XFILLER_14_229 vpwr vgnd scs8hd_fill_2
XFILLER_6_406 vgnd vpwr scs8hd_fill_1
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_64_118 vgnd vpwr scs8hd_decap_6
XFILLER_49_159 vgnd vpwr scs8hd_decap_12
XFILLER_45_332 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_324 vgnd vpwr scs8hd_decap_12
XFILLER_13_262 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_63_184 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_402 vgnd vpwr scs8hd_decap_4
XFILLER_59_39 vgnd vpwr scs8hd_decap_12
XFILLER_46_129 vgnd vpwr scs8hd_decap_12
XFILLER_27_387 vgnd vpwr scs8hd_decap_12
XFILLER_27_310 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ right_width_0_height_0__pin_5_ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_42_379 vgnd vpwr scs8hd_decap_12
XFILLER_24_97 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_6_269 vgnd vpwr scs8hd_decap_3
XFILLER_10_276 vpwr vgnd scs8hd_fill_2
XFILLER_60_154 vgnd vpwr scs8hd_decap_12
XFILLER_45_184 vgnd vpwr scs8hd_decap_12
XFILLER_33_357 vpwr vgnd scs8hd_fill_2
XFILLER_33_302 vgnd vpwr scs8hd_fill_1
XFILLER_18_398 vgnd vpwr scs8hd_decap_8
XFILLER_18_365 vpwr vgnd scs8hd_fill_2
XFILLER_18_332 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_280 vpwr vgnd scs8hd_fill_2
XFILLER_28_129 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_51_110 vgnd vpwr scs8hd_decap_12
XPHY_319 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_308 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_357 vgnd vpwr scs8hd_decap_8
XFILLER_59_232 vgnd vpwr scs8hd_decap_12
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_19_53 vgnd vpwr scs8hd_decap_6
XFILLER_10_66 vpwr vgnd scs8hd_fill_2
XFILLER_42_154 vgnd vpwr scs8hd_decap_12
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_19_75 vpwr vgnd scs8hd_fill_2
XFILLER_51_62 vgnd vpwr scs8hd_decap_12
XFILLER_51_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_250 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_140 vpwr vgnd scs8hd_fill_2
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_202 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_209 vpwr vgnd scs8hd_fill_2
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_121 vgnd vpwr scs8hd_decap_12
XPHY_127 vgnd vpwr scs8hd_decap_3
XFILLER_24_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_349 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _35_/HI ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
XFILLER_21_87 vpwr vgnd scs8hd_fill_2
XFILLER_21_54 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_47_268 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_227 vgnd vpwr scs8hd_decap_12
XFILLER_30_124 vgnd vpwr scs8hd_decap_12
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_7_56 vgnd vpwr scs8hd_decap_3
XFILLER_7_353 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _40_/HI
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_45_lower vgnd vpwr scs8hd_mux2_1
XFILLER_46_290 vgnd vpwr scs8hd_decap_3
XFILLER_61_293 vgnd vpwr scs8hd_decap_12
XFILLER_21_179 vgnd vpwr scs8hd_decap_4
XFILLER_29_213 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_227 vgnd vpwr scs8hd_decap_12
XFILLER_16_32 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_4_334 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_378 vgnd vpwr scs8hd_decap_12
XFILLER_35_216 vpwr vgnd scs8hd_fill_2
XPHY_491 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_480 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ bottom_width_0_height_0__pin_25_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_1_326 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_17_216 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_74 vgnd vpwr scs8hd_decap_12
XFILLER_25_293 vpwr vgnd scs8hd_fill_2
XFILLER_4_131 vpwr vgnd scs8hd_fill_2
XFILLER_48_341 vgnd vpwr scs8hd_fill_1
XFILLER_0_392 vpwr vgnd scs8hd_fill_2
XFILLER_4_46 vgnd vpwr scs8hd_decap_3
XFILLER_31_274 vpwr vgnd scs8hd_fill_2
XFILLER_31_241 vgnd vpwr scs8hd_decap_3
XFILLER_58_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_352 vgnd vpwr scs8hd_decap_3
XFILLER_54_366 vpwr vgnd scs8hd_fill_2
XFILLER_22_274 vgnd vpwr scs8hd_fill_1
XFILLER_14_219 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_123 vpwr vgnd scs8hd_fill_2
XFILLER_57_171 vgnd vpwr scs8hd_decap_12
XFILLER_45_344 vgnd vpwr scs8hd_decap_3
XFILLER_9_212 vpwr vgnd scs8hd_fill_2
XFILLER_9_223 vpwr vgnd scs8hd_fill_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_3
XFILLER_9_267 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _51_/HI ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_36_300 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_196 vgnd vpwr scs8hd_decap_12
XFILLER_51_358 vpwr vgnd scs8hd_fill_2
XFILLER_36_388 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_54_141 vgnd vpwr scs8hd_decap_12
XFILLER_42_303 vgnd vpwr scs8hd_decap_3
XFILLER_39_171 vgnd vpwr scs8hd_decap_12
XFILLER_27_399 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_347 vgnd vpwr scs8hd_fill_1
XFILLER_24_32 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_49_62 vgnd vpwr scs8hd_decap_12
XFILLER_49_51 vgnd vpwr scs8hd_decap_8
XFILLER_18_344 vpwr vgnd scs8hd_fill_2
XFILLER_18_311 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_60_166 vgnd vpwr scs8hd_decap_12
XFILLER_45_196 vgnd vpwr scs8hd_decap_12
XFILLER_33_325 vpwr vgnd scs8hd_fill_2
XFILLER_53_3 vgnd vpwr scs8hd_decap_12
XFILLER_41_380 vgnd vpwr scs8hd_decap_12
X_79_ right_width_0_height_0__pin_40_lower right_width_0_height_0__pin_40_upper vgnd
+ vpwr scs8hd_buf_2
XFILLER_56_406 vgnd vpwr scs8hd_fill_1
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XFILLER_24_325 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XPHY_309 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0_0_clk/X ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ top_width_0_height_0__pin_33_ Test_en vgnd vpwr scs8hd_sdfxbp_1
XFILLER_42_166 vgnd vpwr scs8hd_decap_12
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _41_/HI vgnd vpwr scs8hd_diode_2
XFILLER_51_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_38_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_152 vgnd vpwr scs8hd_fill_1
XFILLER_33_188 vgnd vpwr scs8hd_fill_1
XFILLER_21_317 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_280 vgnd vpwr scs8hd_decap_12
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XPHY_106 vgnd vpwr scs8hd_decap_3
XFILLER_24_133 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_199 vpwr vgnd scs8hd_fill_2
XFILLER_20_394 vgnd vpwr scs8hd_decap_3
XFILLER_21_66 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_239 vgnd vpwr scs8hd_decap_12
XFILLER_47_236 vpwr vgnd scs8hd_fill_2
XFILLER_30_136 vgnd vpwr scs8hd_decap_12
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_15_133 vpwr vgnd scs8hd_fill_2
XFILLER_7_365 vgnd vpwr scs8hd_fill_1
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_247 vgnd vpwr scs8hd_fill_1
XFILLER_21_136 vgnd vpwr scs8hd_fill_1
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_203 vpwr vgnd scs8hd_fill_2
XFILLER_44_239 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_88 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_357 vpwr vgnd scs8hd_fill_2
XFILLER_57_62 vgnd vpwr scs8hd_decap_12
XFILLER_57_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _63_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_280 vpwr vgnd scs8hd_fill_2
XPHY_492 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_481 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_470 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_272 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ bottom_width_0_height_0__pin_27_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_26_206 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_34_261 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ bottom_width_0_height_0__pin_24_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _46_/HI
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_353 vgnd vpwr scs8hd_decap_6
XFILLER_43_86 vgnd vpwr scs8hd_decap_12
XFILLER_40_264 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_36 vgnd vpwr scs8hd_fill_1
XFILLER_4_176 vpwr vgnd scs8hd_fill_2
XFILLER_48_375 vpwr vgnd scs8hd_fill_2
XFILLER_63_367 vgnd vpwr scs8hd_decap_12
XFILLER_31_253 vgnd vpwr scs8hd_decap_4
XFILLER_31_220 vpwr vgnd scs8hd_fill_2
XFILLER_23_209 vpwr vgnd scs8hd_fill_2
XFILLER_58_117 vgnd vpwr scs8hd_decap_12
XFILLER_54_356 vpwr vgnd scs8hd_fill_2
XFILLER_54_323 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_389 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ right_width_0_height_0__pin_2_ vgnd vpwr scs8hd_diode_2
XFILLER_13_45 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_301 vpwr vgnd scs8hd_fill_2
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_367 vgnd vpwr scs8hd_decap_4
XFILLER_13_231 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _58_/HI
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_235 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_304 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_323 vgnd vpwr scs8hd_decap_8
XFILLER_51_337 vpwr vgnd scs8hd_fill_2
XFILLER_51_315 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_367 vgnd vpwr scs8hd_decap_6
XFILLER_27_345 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_267 vgnd vpwr scs8hd_decap_8
XFILLER_10_289 vgnd vpwr scs8hd_decap_3
XFILLER_49_74 vgnd vpwr scs8hd_decap_12
XFILLER_1_26 vpwr vgnd scs8hd_fill_2
XFILLER_60_178 vgnd vpwr scs8hd_decap_12
XFILLER_41_392 vgnd vpwr scs8hd_decap_12
XFILLER_18_389 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
X_78_ right_width_0_height_0__pin_39_lower right_width_0_height_0__pin_39_upper vgnd
+ vpwr scs8hd_buf_2
XFILLER_51_123 vgnd vpwr scs8hd_decap_12
XFILLER_24_315 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ right_width_0_height_0__pin_14_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_46 vgnd vpwr scs8hd_fill_1
XFILLER_59_245 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_153 vgnd vpwr scs8hd_fill_1
XFILLER_19_99 vpwr vgnd scs8hd_fill_2
XFILLER_42_178 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XFILLER_27_197 vpwr vgnd scs8hd_fill_2
XFILLER_27_175 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_285 vpwr vgnd scs8hd_fill_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XFILLER_18_120 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_215 vgnd vpwr scs8hd_decap_12
XPHY_129 vgnd vpwr scs8hd_decap_3
XFILLER_64_292 vgnd vpwr scs8hd_decap_12
XPHY_118 vgnd vpwr scs8hd_decap_3
XPHY_107 vgnd vpwr scs8hd_decap_3
XFILLER_21_23 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_55_281 vgnd vpwr scs8hd_decap_12
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_112 vpwr vgnd scs8hd_fill_2
XFILLER_15_123 vgnd vpwr scs8hd_decap_3
XFILLER_30_148 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_270 vgnd vpwr scs8hd_decap_3
XFILLER_29_237 vgnd vpwr scs8hd_decap_6
XFILLER_52_251 vgnd vpwr scs8hd_decap_4
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_16_78 vgnd vpwr scs8hd_decap_4
XFILLER_8_119 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _36_/HI vgnd vpwr scs8hd_diode_2
XFILLER_57_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_240 vpwr vgnd scs8hd_fill_2
XFILLER_35_229 vpwr vgnd scs8hd_fill_2
XPHY_493 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_482 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_471 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_460 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_163 vgnd vpwr scs8hd_decap_6
XFILLER_11_192 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_306 vgnd vpwr scs8hd_fill_1
XFILLER_8_90 vpwr vgnd scs8hd_fill_2
XFILLER_57_332 vgnd vpwr scs8hd_decap_4
XFILLER_57_310 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_99 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ bottom_width_0_height_0__pin_30_ vgnd vpwr scs8hd_diode_2
XFILLER_43_98 vgnd vpwr scs8hd_decap_12
XFILLER_40_276 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_100 vpwr vgnd scs8hd_fill_2
XFILLER_4_144 vpwr vgnd scs8hd_fill_2
XFILLER_48_398 vgnd vpwr scs8hd_decap_8
XFILLER_63_379 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_262 vgnd vpwr scs8hd_decap_12
XFILLER_31_287 vpwr vgnd scs8hd_fill_2
XPHY_290 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_129 vgnd vpwr scs8hd_decap_12
XFILLER_39_321 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_210 vgnd vpwr scs8hd_decap_4
XFILLER_22_276 vgnd vpwr scs8hd_decap_4
XFILLER_22_254 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_57_184 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_243 vgnd vpwr scs8hd_fill_1
XFILLER_13_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_346 vgnd vpwr scs8hd_decap_12
XFILLER_36_313 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_27_313 vpwr vgnd scs8hd_fill_2
XFILLER_27_302 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_54_154 vgnd vpwr scs8hd_decap_12
XFILLER_50_382 vgnd vpwr scs8hd_decap_12
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_206 vpwr vgnd scs8hd_fill_2
XFILLER_49_86 vgnd vpwr scs8hd_decap_12
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_45_110 vgnd vpwr scs8hd_decap_12
XFILLER_18_324 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ccff_head vgnd vpwr scs8hd_diode_2
X_77_ right_width_0_height_0__pin_38_lower right_width_0_height_0__pin_38_upper vgnd
+ vpwr scs8hd_buf_2
XFILLER_51_135 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ right_width_0_height_0__pin_13_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_390 vgnd vpwr scs8hd_decap_12
XFILLER_3_209 vpwr vgnd scs8hd_fill_2
XFILLER_59_257 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_19_23 vgnd vpwr scs8hd_fill_1
XFILLER_50_190 vgnd vpwr scs8hd_decap_12
XFILLER_51_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_242 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_227 vgnd vpwr scs8hd_decap_12
XPHY_119 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_decap_3
XFILLER_24_168 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_20_363 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_55_293 vgnd vpwr scs8hd_decap_12
XFILLER_46_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_48 vgnd vpwr scs8hd_decap_8
XFILLER_7_301 vpwr vgnd scs8hd_fill_2
XFILLER_7_323 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_11_330 vgnd vpwr scs8hd_decap_12
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_367 vgnd vpwr scs8hd_decap_12
XFILLER_53_208 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_14_190 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_315 vpwr vgnd scs8hd_fill_2
XFILLER_4_326 vpwr vgnd scs8hd_fill_2
XFILLER_57_86 vgnd vpwr scs8hd_decap_12
XFILLER_35_208 vgnd vpwr scs8hd_fill_1
XPHY_461 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_450 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_285 vpwr vgnd scs8hd_fill_2
XPHY_494 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_483 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_472 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_131 vpwr vgnd scs8hd_fill_2
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_7_197 vpwr vgnd scs8hd_fill_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_392 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XFILLER_4_167 vpwr vgnd scs8hd_fill_2
XFILLER_4_189 vpwr vgnd scs8hd_fill_2
XFILLER_48_344 vpwr vgnd scs8hd_fill_2
XFILLER_48_333 vgnd vpwr scs8hd_decap_3
XFILLER_31_233 vpwr vgnd scs8hd_fill_2
XPHY_291 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_274 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_344 vgnd vpwr scs8hd_decap_8
XFILLER_54_314 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_266 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ bottom_width_0_height_0__pin_24_ vgnd vpwr scs8hd_diode_2
XFILLER_10_406 vgnd vpwr scs8hd_fill_1
XFILLER_57_196 vgnd vpwr scs8hd_decap_12
XFILLER_54_32 vgnd vpwr scs8hd_decap_12
XFILLER_45_358 vpwr vgnd scs8hd_fill_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_200 vgnd vpwr scs8hd_decap_12
XFILLER_13_266 vgnd vpwr scs8hd_decap_12
XFILLER_48_141 vgnd vpwr scs8hd_decap_12
XFILLER_44_391 vgnd vpwr scs8hd_decap_6
XFILLER_36_358 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_281 vpwr vgnd scs8hd_fill_2
XFILLER_59_406 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_70 vpwr vgnd scs8hd_fill_2
XFILLER_39_196 vgnd vpwr scs8hd_decap_12
XFILLER_27_358 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_166 vgnd vpwr scs8hd_decap_12
XFILLER_50_394 vgnd vpwr scs8hd_decap_3
XFILLER_42_328 vgnd vpwr scs8hd_decap_8
XFILLER_42_317 vpwr vgnd scs8hd_fill_2
XFILLER_35_380 vgnd vpwr scs8hd_decap_12
XFILLER_24_68 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_218 vpwr vgnd scs8hd_fill_2
XFILLER_49_98 vgnd vpwr scs8hd_decap_12
XFILLER_18_369 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_350 vpwr vgnd scs8hd_fill_2
XFILLER_14_90 vpwr vgnd scs8hd_fill_2
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
XFILLER_5_284 vpwr vgnd scs8hd_fill_2
X_76_ right_width_0_height_0__pin_37_lower right_width_0_height_0__pin_37_upper vgnd
+ vpwr scs8hd_buf_2
XFILLER_51_147 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ right_width_0_height_0__pin_12_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_269 vgnd vpwr scs8hd_decap_12
XFILLER_27_111 vgnd vpwr scs8hd_decap_8
XFILLER_19_79 vpwr vgnd scs8hd_fill_2
XFILLER_15_306 vpwr vgnd scs8hd_fill_2
XFILLER_2_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_144 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_51_3 vgnd vpwr scs8hd_decap_12
XFILLER_64_261 vgnd vpwr scs8hd_decap_12
XFILLER_56_239 vgnd vpwr scs8hd_decap_12
X_59_ _59_/HI _59_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_93 vpwr vgnd scs8hd_fill_2
XFILLER_2_82 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_decap_3
XFILLER_32_180 vgnd vpwr scs8hd_decap_4
XFILLER_20_342 vpwr vgnd scs8hd_fill_2
XFILLER_20_386 vgnd vpwr scs8hd_decap_8
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XFILLER_46_44 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_103 vgnd vpwr scs8hd_decap_4
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XFILLER_7_379 vgnd vpwr scs8hd_decap_12
XFILLER_11_342 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_61_220 vgnd vpwr scs8hd_decap_12
XFILLER_38_239 vgnd vpwr scs8hd_decap_8
XFILLER_21_139 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_390 vgnd vpwr scs8hd_decap_6
XFILLER_29_217 vgnd vpwr scs8hd_decap_3
XFILLER_16_47 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XFILLER_20_183 vgnd vpwr scs8hd_fill_1
XFILLER_12_139 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_261 vgnd vpwr scs8hd_decap_12
XPHY_495 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_484 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_473 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_462 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_451 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_440 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_297 vpwr vgnd scs8hd_fill_2
XFILLER_43_220 vgnd vpwr scs8hd_decap_12
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ right_width_0_height_0__pin_2_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_367 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_297 vpwr vgnd scs8hd_fill_2
XFILLER_25_253 vpwr vgnd scs8hd_fill_2
XFILLER_0_396 vgnd vpwr scs8hd_decap_6
XFILLER_31_245 vpwr vgnd scs8hd_fill_2
XPHY_292 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_54_337 vgnd vpwr scs8hd_decap_4
XFILLER_39_367 vgnd vpwr scs8hd_decap_4
XFILLER_39_301 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _61_/HI
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_38_lower vgnd vpwr scs8hd_mux2_1
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_127 vpwr vgnd scs8hd_fill_2
XFILLER_1_138 vpwr vgnd scs8hd_fill_2
XFILLER_54_44 vgnd vpwr scs8hd_decap_12
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_9_216 vgnd vpwr scs8hd_decap_4
XFILLER_9_227 vgnd vpwr scs8hd_decap_8
XFILLER_13_212 vgnd vpwr scs8hd_decap_3
XFILLER_13_278 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_271 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_82 vpwr vgnd scs8hd_fill_2
XFILLER_54_178 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_392 vgnd vpwr scs8hd_decap_12
XFILLER_24_36 vgnd vpwr scs8hd_decap_4
XFILLER_10_215 vpwr vgnd scs8hd_fill_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_123 vgnd vpwr scs8hd_decap_12
XFILLER_33_329 vpwr vgnd scs8hd_fill_2
XFILLER_18_348 vpwr vgnd scs8hd_fill_2
XFILLER_18_337 vgnd vpwr scs8hd_decap_3
XFILLER_41_362 vpwr vgnd scs8hd_fill_2
X_75_ right_width_0_height_0__pin_36_lower right_width_0_height_0__pin_36_upper vgnd
+ vpwr scs8hd_buf_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XFILLER_24_307 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_159 vgnd vpwr scs8hd_decap_12
XFILLER_24_329 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_27_123 vgnd vpwr scs8hd_decap_12
XFILLER_15_329 vpwr vgnd scs8hd_fill_2
XFILLER_23_362 vpwr vgnd scs8hd_fill_2
XFILLER_23_351 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_90 vgnd vpwr scs8hd_decap_3
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XFILLER_18_178 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_44_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _51_/HI vgnd vpwr scs8hd_diode_2
XFILLER_64_273 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
X_58_ _58_/HI _58_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_6
XFILLER_20_398 vgnd vpwr scs8hd_decap_8
XFILLER_20_376 vpwr vgnd scs8hd_fill_2
XFILLER_46_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_44 vgnd vpwr scs8hd_decap_12
XFILLER_23_181 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_39 vgnd vpwr scs8hd_decap_3
XFILLER_7_347 vgnd vpwr scs8hd_decap_3
XFILLER_11_354 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_81 vgnd vpwr scs8hd_decap_8
XFILLER_61_232 vgnd vpwr scs8hd_decap_12
XFILLER_46_295 vpwr vgnd scs8hd_fill_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XFILLER_29_229 vpwr vgnd scs8hd_fill_2
XFILLER_29_207 vgnd vpwr scs8hd_decap_4
XFILLER_52_276 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_232 vgnd vpwr scs8hd_decap_6
XFILLER_28_284 vgnd vpwr scs8hd_decap_8
XFILLER_28_273 vpwr vgnd scs8hd_fill_2
XPHY_496 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_485 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_474 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_463 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_452 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_441 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_430 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_162 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_195 vpwr vgnd scs8hd_fill_2
XFILLER_34_265 vpwr vgnd scs8hd_fill_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_19_273 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ bottom_width_0_height_0__pin_21_ vgnd vpwr scs8hd_diode_2
XFILLER_8_82 vgnd vpwr scs8hd_decap_8
XFILLER_8_93 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ right_width_0_height_0__pin_1_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XFILLER_25_276 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_364 vpwr vgnd scs8hd_fill_2
XFILLER_0_342 vgnd vpwr scs8hd_decap_3
XFILLER_0_331 vgnd vpwr scs8hd_decap_3
XFILLER_31_224 vpwr vgnd scs8hd_fill_2
XFILLER_16_276 vpwr vgnd scs8hd_fill_2
XFILLER_16_232 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_257 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XPHY_293 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_49 vgnd vpwr scs8hd_decap_12
XFILLER_57_110 vgnd vpwr scs8hd_decap_12
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_54_56 vgnd vpwr scs8hd_decap_12
XFILLER_53_382 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_63_135 vgnd vpwr scs8hd_decap_12
XFILLER_48_154 vgnd vpwr scs8hd_decap_12
XFILLER_36_305 vpwr vgnd scs8hd_fill_2
XFILLER_28_90 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_183 vgnd vpwr scs8hd_fill_1
XFILLER_51_319 vgnd vpwr scs8hd_decap_12
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_35_371 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_135 vgnd vpwr scs8hd_decap_12
XFILLER_1_19 vgnd vpwr scs8hd_decap_3
XFILLER_60_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_26_360 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_5_264 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XFILLER_5_297 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
X_74_ right_width_0_height_0__pin_35_lower right_width_0_height_0__pin_35_upper vgnd
+ vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_32_385 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _53_/HI vgnd vpwr scs8hd_diode_2
XFILLER_27_135 vgnd vpwr scs8hd_decap_12
XFILLER_19_26 vpwr vgnd scs8hd_fill_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_42_105 vgnd vpwr scs8hd_decap_12
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_289 vpwr vgnd scs8hd_fill_2
XFILLER_2_267 vpwr vgnd scs8hd_fill_2
XFILLER_2_201 vpwr vgnd scs8hd_fill_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_157 vpwr vgnd scs8hd_fill_2
XFILLER_18_124 vpwr vgnd scs8hd_fill_2
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_91 vgnd vpwr scs8hd_decap_3
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_341 vpwr vgnd scs8hd_fill_2
XFILLER_49_271 vpwr vgnd scs8hd_fill_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xclkbuf_1_1_0_clk clkbuf_0_clk/X clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_clkbuf_1
XFILLER_64_230 vgnd vpwr scs8hd_decap_12
X_57_ _57_/HI _57_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_21_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_333 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ right_width_0_height_0__pin_15_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_208 vgnd vpwr scs8hd_decap_12
XFILLER_46_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ bottom_width_0_height_0__pin_27_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_or2_1
XFILLER_15_116 vgnd vpwr scs8hd_decap_4
XFILLER_62_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_7_315 vpwr vgnd scs8hd_fill_2
XFILLER_11_93 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_46_285 vgnd vpwr scs8hd_decap_3
XFILLER_25_403 vgnd vpwr scs8hd_decap_4
XFILLER_52_255 vgnd vpwr scs8hd_fill_1
XFILLER_40_406 vgnd vpwr scs8hd_fill_1
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_163 vgnd vpwr scs8hd_decap_12
XFILLER_4_307 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_406 vgnd vpwr scs8hd_fill_1
XPHY_497 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_486 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_475 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_464 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_453 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_442 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_431 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_420 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_70 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_362 vpwr vgnd scs8hd_fill_2
XFILLER_19_230 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_406 vgnd vpwr scs8hd_fill_1
XFILLER_19_296 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ right_width_0_height_0__pin_0_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_8_61 vgnd vpwr scs8hd_decap_8
XFILLER_57_336 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_40_247 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_104 vpwr vgnd scs8hd_fill_2
XFILLER_4_148 vgnd vpwr scs8hd_decap_3
XFILLER_63_306 vgnd vpwr scs8hd_decap_12
XFILLER_48_369 vgnd vpwr scs8hd_decap_4
XFILLER_48_325 vgnd vpwr scs8hd_decap_8
XFILLER_31_203 vpwr vgnd scs8hd_fill_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_81 vgnd vpwr scs8hd_decap_3
XFILLER_16_211 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_3
XPHY_294 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_54_328 vgnd vpwr scs8hd_decap_6
XFILLER_47_380 vpwr vgnd scs8hd_fill_2
XFILLER_39_358 vpwr vgnd scs8hd_fill_2
XFILLER_62_361 vgnd vpwr scs8hd_decap_12
XFILLER_30_280 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_39 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_45_306 vgnd vpwr scs8hd_decap_3
XFILLER_54_68 vgnd vpwr scs8hd_decap_12
XFILLER_53_394 vgnd vpwr scs8hd_decap_12
XFILLER_45_328 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_38_391 vgnd vpwr scs8hd_decap_6
XFILLER_13_258 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XFILLER_63_147 vgnd vpwr scs8hd_decap_12
XFILLER_48_166 vgnd vpwr scs8hd_decap_12
XFILLER_29_391 vgnd vpwr scs8hd_decap_12
XFILLER_44_372 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_262 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ccff_head ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_27_306 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_342 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_206 vgnd vpwr scs8hd_decap_8
XFILLER_45_147 vgnd vpwr scs8hd_decap_12
XFILLER_18_328 vpwr vgnd scs8hd_fill_2
XFILLER_60_117 vgnd vpwr scs8hd_decap_12
XFILLER_26_372 vgnd vpwr scs8hd_decap_12
XFILLER_5_221 vgnd vpwr scs8hd_decap_4
XFILLER_5_276 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
X_73_ right_width_0_height_0__pin_34_lower right_width_0_height_0__pin_34_upper vgnd
+ vpwr scs8hd_buf_2
XFILLER_32_331 vpwr vgnd scs8hd_fill_2
XFILLER_32_320 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_147 vgnd vpwr scs8hd_decap_6
XFILLER_19_49 vpwr vgnd scs8hd_fill_2
XFILLER_42_117 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_235 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_331 vgnd vpwr scs8hd_decap_4
XPHY_92 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_242 vgnd vpwr scs8hd_decap_6
X_56_ _56_/HI _56_/LO vgnd vpwr scs8hd_conb_1
XFILLER_24_139 vgnd vpwr scs8hd_fill_1
XFILLER_20_312 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_55_220 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_128 vgnd vpwr scs8hd_decap_3
XFILLER_62_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_161 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_7_327 vgnd vpwr scs8hd_decap_12
XFILLER_11_301 vgnd vpwr scs8hd_decap_4
XFILLER_11_367 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_19_401 vgnd vpwr scs8hd_decap_6
XFILLER_61_245 vgnd vpwr scs8hd_decap_12
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ bottom_width_0_height_0__pin_18_ vgnd vpwr scs8hd_diode_2
XFILLER_14_194 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_297 vpwr vgnd scs8hd_fill_2
XFILLER_37_275 vgnd vpwr scs8hd_fill_1
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
X_39_ _39_/HI _39_/LO vgnd vpwr scs8hd_conb_1
XFILLER_52_267 vgnd vpwr scs8hd_decap_8
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _52_/HI
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_35_lower vgnd vpwr scs8hd_mux2_1
XFILLER_20_175 vgnd vpwr scs8hd_decap_8
XFILLER_20_186 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XPHY_443 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_432 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_421 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_289 vpwr vgnd scs8hd_fill_2
XFILLER_43_245 vpwr vgnd scs8hd_fill_2
XPHY_410 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_498 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_487 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_476 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_465 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_454 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_93 vgnd vpwr scs8hd_fill_1
XFILLER_22_82 vpwr vgnd scs8hd_fill_2
Xclkbuf_1_0_0_clk clkbuf_0_clk/X clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_clkbuf_1
XFILLER_7_135 vpwr vgnd scs8hd_fill_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_142 vpwr vgnd scs8hd_fill_2
XFILLER_11_153 vgnd vpwr scs8hd_decap_3
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
XFILLER_34_234 vgnd vpwr scs8hd_decap_8
XFILLER_8_40 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_57_359 vgnd vpwr scs8hd_fill_1
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XFILLER_43_15 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_43_59 vpwr vgnd scs8hd_fill_2
XFILLER_0_311 vgnd vpwr scs8hd_fill_1
XFILLER_4_127 vpwr vgnd scs8hd_fill_2
XFILLER_63_318 vgnd vpwr scs8hd_decap_12
XFILLER_48_348 vpwr vgnd scs8hd_fill_2
XFILLER_48_337 vgnd vpwr scs8hd_decap_4
XFILLER_16_201 vpwr vgnd scs8hd_fill_2
XFILLER_31_237 vpwr vgnd scs8hd_fill_2
XPHY_295 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_71 vgnd vpwr scs8hd_decap_4
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _41_/HI
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_44_lower vgnd vpwr scs8hd_mux2_1
XFILLER_39_315 vgnd vpwr scs8hd_decap_4
XFILLER_3_182 vgnd vpwr scs8hd_fill_1
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_47_392 vgnd vpwr scs8hd_decap_12
XFILLER_22_215 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_123 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_53_362 vpwr vgnd scs8hd_fill_2
XFILLER_63_159 vgnd vpwr scs8hd_decap_12
XFILLER_48_178 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_241 vpwr vgnd scs8hd_fill_2
XFILLER_8_285 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _54_/HI vgnd vpwr scs8hd_diode_2
XFILLER_50_365 vpwr vgnd scs8hd_fill_2
XFILLER_35_362 vpwr vgnd scs8hd_fill_2
XFILLER_50_398 vgnd vpwr scs8hd_decap_8
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_2_406 vgnd vpwr scs8hd_fill_1
XFILLER_45_159 vgnd vpwr scs8hd_decap_12
XFILLER_18_307 vpwr vgnd scs8hd_fill_2
XFILLER_60_129 vgnd vpwr scs8hd_decap_12
XFILLER_41_376 vpwr vgnd scs8hd_fill_2
XFILLER_41_310 vgnd vpwr scs8hd_decap_4
XFILLER_26_384 vgnd vpwr scs8hd_decap_12
XANTENNA__70__A bottom_width_0_height_0__pin_48_lower vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
X_72_ bottom_width_0_height_0__pin_50_ bottom_width_0_height_0__pin_51_ vgnd vpwr
+ scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_362 vpwr vgnd scs8hd_fill_2
XFILLER_32_398 vgnd vpwr scs8hd_decap_8
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_51_59 vpwr vgnd scs8hd_fill_2
XFILLER_51_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_129 vgnd vpwr scs8hd_decap_12
XFILLER_23_321 vpwr vgnd scs8hd_fill_2
XFILLER_23_310 vpwr vgnd scs8hd_fill_2
XFILLER_58_251 vgnd vpwr scs8hd_decap_12
XFILLER_18_115 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_61_405 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_18_148 vgnd vpwr scs8hd_decap_4
XANTENNA__65__A bottom_width_0_height_0__pin_43_lower vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_365 vgnd vpwr scs8hd_decap_8
XPHY_93 vgnd vpwr scs8hd_decap_3
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XFILLER_14_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_49_284 vpwr vgnd scs8hd_fill_2
XFILLER_49_240 vpwr vgnd scs8hd_fill_2
X_55_ _55_/HI _55_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_97 vgnd vpwr scs8hd_decap_3
XFILLER_2_86 vgnd vpwr scs8hd_decap_4
XFILLER_2_42 vpwr vgnd scs8hd_fill_2
XFILLER_1_291 vpwr vgnd scs8hd_fill_2
XFILLER_20_346 vpwr vgnd scs8hd_fill_2
XFILLER_20_324 vgnd vpwr scs8hd_decap_3
XFILLER_17_192 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_391 vgnd vpwr scs8hd_decap_12
XFILLER_46_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_55_232 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_107 vgnd vpwr scs8hd_fill_1
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
XFILLER_23_173 vpwr vgnd scs8hd_fill_2
XFILLER_7_339 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_379 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_11_51 vgnd vpwr scs8hd_decap_4
XFILLER_46_243 vpwr vgnd scs8hd_fill_2
XFILLER_61_257 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_52_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_350 vgnd vpwr scs8hd_decap_6
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_52_202 vgnd vpwr scs8hd_decap_12
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
X_38_ _38_/HI _38_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_121 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_28_210 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_477 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_466 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_455 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_444 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_433 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_422 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_268 vpwr vgnd scs8hd_fill_2
XPHY_411 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_400 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_110 vpwr vgnd scs8hd_fill_2
XPHY_499 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_488 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_169 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ right_width_0_height_0__pin_12_ vgnd vpwr scs8hd_diode_2
XFILLER_3_331 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_202 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_57_349 vpwr vgnd scs8hd_fill_2
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XFILLER_43_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_213 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_305 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_17_50 vgnd vpwr scs8hd_decap_4
XFILLER_16_235 vpwr vgnd scs8hd_fill_2
XANTENNA__73__A right_width_0_height_0__pin_34_lower vgnd vpwr scs8hd_diode_2
XFILLER_31_249 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_296 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_54_319 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_135 vgnd vpwr scs8hd_decap_12
XFILLER_54_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ right_width_0_height_0__pin_15_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_or2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA__68__A bottom_width_0_height_0__pin_46_lower vgnd vpwr scs8hd_diode_2
XFILLER_0_175 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_190 vgnd vpwr scs8hd_decap_12
XFILLER_36_319 vpwr vgnd scs8hd_fill_2
XFILLER_29_360 vgnd vpwr scs8hd_decap_6
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
XFILLER_28_82 vgnd vpwr scs8hd_decap_8
XFILLER_60_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_220 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_31 vgnd vpwr scs8hd_fill_1
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_86 vpwr vgnd scs8hd_fill_2
XFILLER_54_105 vgnd vpwr scs8hd_decap_12
XFILLER_39_135 vgnd vpwr scs8hd_decap_12
XFILLER_50_322 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _34_/HI
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_10_219 vpwr vgnd scs8hd_fill_2
XFILLER_49_59 vpwr vgnd scs8hd_fill_2
XFILLER_49_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_53_171 vgnd vpwr scs8hd_decap_12
XFILLER_41_333 vgnd vpwr scs8hd_decap_12
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
XFILLER_26_396 vgnd vpwr scs8hd_fill_1
XFILLER_14_40 vgnd vpwr scs8hd_decap_3
XFILLER_14_62 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
X_71_ bottom_width_0_height_0__pin_49_lower bottom_width_0_height_0__pin_49_upper
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_59_208 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_51_27 vgnd vpwr scs8hd_decap_12
XFILLER_50_141 vgnd vpwr scs8hd_decap_12
XFILLER_23_344 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _39_/HI ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
XFILLER_2_215 vgnd vpwr scs8hd_fill_1
XFILLER_58_263 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_94 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_26_193 vpwr vgnd scs8hd_fill_2
XFILLER_25_50 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_14_300 vgnd vpwr scs8hd_decap_8
XFILLER_14_377 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_32 vpwr vgnd scs8hd_fill_2
XFILLER_64_211 vgnd vpwr scs8hd_decap_6
XFILLER_52_406 vgnd vpwr scs8hd_fill_1
X_54_ _54_/HI _54_/LO vgnd vpwr scs8hd_conb_1
XFILLER_17_171 vpwr vgnd scs8hd_fill_2
XFILLER_2_65 vpwr vgnd scs8hd_fill_2
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _58_/HI vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_46_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_196 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _37_/HI vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XANTENNA__76__A right_width_0_height_0__pin_37_lower vgnd vpwr scs8hd_diode_2
XFILLER_46_299 vpwr vgnd scs8hd_fill_2
XFILLER_34_406 vgnd vpwr scs8hd_fill_1
XFILLER_61_269 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
X_37_ _37_/HI _37_/LO vgnd vpwr scs8hd_conb_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_199 vgnd vpwr scs8hd_decap_12
XFILLER_57_15 vgnd vpwr scs8hd_decap_12
XFILLER_57_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_406 vgnd vpwr scs8hd_fill_1
XPHY_489 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_478 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_467 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_456 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_445 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_434 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_423 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_412 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_401 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_104 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_310 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_188 vgnd vpwr scs8hd_decap_4
XFILLER_34_269 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_97 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_57_339 vgnd vpwr scs8hd_fill_1
XFILLER_57_306 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_25_203 vpwr vgnd scs8hd_fill_2
XFILLER_43_39 vgnd vpwr scs8hd_decap_12
XFILLER_40_239 vgnd vpwr scs8hd_decap_8
XFILLER_25_236 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_368 vpwr vgnd scs8hd_fill_2
XFILLER_56_361 vgnd vpwr scs8hd_decap_6
XFILLER_56_350 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_228 vgnd vpwr scs8hd_fill_1
XPHY_297 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_286 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _55_/HI ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_4
XFILLER_3_162 vpwr vgnd scs8hd_fill_2
XFILLER_58_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_228 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_147 vgnd vpwr scs8hd_decap_12
XFILLER_54_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_217 vgnd vpwr scs8hd_decap_3
XFILLER_13_239 vpwr vgnd scs8hd_fill_2
XFILLER_0_121 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_309 vpwr vgnd scs8hd_fill_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_3
XFILLER_44_331 vgnd vpwr scs8hd_decap_3
XFILLER_44_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_232 vgnd vpwr scs8hd_decap_3
XFILLER_8_254 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_298 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_54_117 vgnd vpwr scs8hd_decap_12
XFILLER_39_147 vgnd vpwr scs8hd_decap_12
XFILLER_50_334 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_27 vgnd vpwr scs8hd_decap_12
XFILLER_41_345 vgnd vpwr scs8hd_decap_3
XFILLER_41_301 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_14_74 vpwr vgnd scs8hd_fill_2
XANTENNA__79__A right_width_0_height_0__pin_40_lower vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_268 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_404 vgnd vpwr scs8hd_decap_3
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XFILLER_17_331 vpwr vgnd scs8hd_fill_2
X_70_ bottom_width_0_height_0__pin_48_lower bottom_width_0_height_0__pin_48_upper
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_386 vpwr vgnd scs8hd_fill_2
XFILLER_51_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_389 vgnd vpwr scs8hd_decap_12
XFILLER_23_367 vgnd vpwr scs8hd_decap_3
XFILLER_2_205 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_128 vgnd vpwr scs8hd_decap_3
XFILLER_18_106 vpwr vgnd scs8hd_fill_2
XPHY_95 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_345 vgnd vpwr scs8hd_fill_1
XFILLER_14_389 vgnd vpwr scs8hd_decap_8
XFILLER_49_220 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
X_53_ _53_/HI _53_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_260 vpwr vgnd scs8hd_fill_2
XFILLER_49_297 vpwr vgnd scs8hd_fill_2
XFILLER_24_109 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_32_186 vgnd vpwr scs8hd_fill_1
XFILLER_20_359 vpwr vgnd scs8hd_fill_2
XFILLER_20_337 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_55_245 vgnd vpwr scs8hd_decap_12
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
XFILLER_23_131 vgnd vpwr scs8hd_decap_3
XFILLER_7_319 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_97 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ right_width_0_height_0__pin_9_ vgnd vpwr scs8hd_diode_2
XFILLER_52_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _32_/HI
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_41_lower vgnd vpwr scs8hd_mux2_1
XFILLER_6_396 vgnd vpwr scs8hd_fill_1
XFILLER_37_245 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
X_36_ _36_/HI _36_/LO vgnd vpwr scs8hd_conb_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_52_215 vgnd vpwr scs8hd_decap_12
XFILLER_37_267 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_145 vpwr vgnd scs8hd_fill_2
XFILLER_57_27 vgnd vpwr scs8hd_decap_12
XPHY_479 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_468 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_457 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_446 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_435 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_424 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_413 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_402 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_127 vpwr vgnd scs8hd_fill_2
XFILLER_22_74 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vgnd vpwr scs8hd_decap_6
XFILLER_19_234 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_32 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _62_/HI vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_303 vgnd vpwr scs8hd_fill_1
XFILLER_0_336 vgnd vpwr scs8hd_decap_3
XFILLER_31_207 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _32_/HI vgnd vpwr scs8hd_diode_2
XFILLER_16_215 vpwr vgnd scs8hd_fill_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XPHY_298 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_287 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_174 vpwr vgnd scs8hd_fill_2
XFILLER_47_340 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_62_398 vgnd vpwr scs8hd_decap_8
XFILLER_30_262 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_284 vpwr vgnd scs8hd_fill_2
XFILLER_57_159 vgnd vpwr scs8hd_decap_12
XFILLER_53_332 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_273 vgnd vpwr scs8hd_fill_1
XFILLER_5_406 vgnd vpwr scs8hd_fill_1
XFILLER_28_73 vgnd vpwr scs8hd_decap_6
XFILLER_44_398 vgnd vpwr scs8hd_decap_8
XFILLER_44_343 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_159 vgnd vpwr scs8hd_decap_12
XFILLER_5_66 vpwr vgnd scs8hd_fill_2
XFILLER_5_99 vgnd vpwr scs8hd_decap_3
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_54_129 vgnd vpwr scs8hd_decap_12
XFILLER_35_376 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_49_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_53_184 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_26_398 vgnd vpwr scs8hd_decap_8
XFILLER_26_332 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _39_/HI vgnd vpwr scs8hd_diode_2
XFILLER_5_236 vpwr vgnd scs8hd_fill_2
XFILLER_14_97 vgnd vpwr scs8hd_decap_8
XFILLER_49_402 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
XFILLER_17_354 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_335 vgnd vpwr scs8hd_fill_1
XFILLER_32_324 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ right_width_0_height_0__pin_3_ vgnd vpwr scs8hd_diode_2
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XFILLER_2_239 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_58_276 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_14_335 vgnd vpwr scs8hd_fill_1
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XFILLER_49_232 vgnd vpwr scs8hd_decap_6
XFILLER_37_405 vpwr vgnd scs8hd_fill_2
X_52_ _52_/HI _52_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_17_184 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_361 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_55_257 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ right_width_0_height_0__pin_3_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_or2_1
XFILLER_23_121 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_46_202 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_121 vgnd vpwr scs8hd_decap_4
XFILLER_14_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
X_35_ _35_/HI _35_/LO vgnd vpwr scs8hd_conb_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_227 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_57_39 vgnd vpwr scs8hd_decap_12
XFILLER_28_202 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_425 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_414 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_403 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_469 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_458 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_447 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_436 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_53 vgnd vpwr scs8hd_decap_8
XFILLER_11_146 vgnd vpwr scs8hd_decap_4
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
XFILLER_22_86 vgnd vpwr scs8hd_decap_6
XFILLER_3_301 vpwr vgnd scs8hd_fill_2
XFILLER_3_367 vgnd vpwr scs8hd_decap_4
XFILLER_42_271 vpwr vgnd scs8hd_fill_2
XFILLER_27_290 vpwr vgnd scs8hd_fill_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_249 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_205 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XPHY_299 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_288 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_300 vgnd vpwr scs8hd_decap_12
XFILLER_58_93 vgnd vpwr scs8hd_decap_12
XFILLER_47_363 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_62_377 vgnd vpwr scs8hd_decap_12
XFILLER_30_274 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_344 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_263 vgnd vpwr scs8hd_fill_1
XFILLER_21_241 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_105 vgnd vpwr scs8hd_decap_12
XFILLER_44_366 vgnd vpwr scs8hd_decap_4
XFILLER_29_352 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_78 vpwr vgnd scs8hd_fill_2
XFILLER_8_267 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_141 vgnd vpwr scs8hd_decap_12
XFILLER_47_171 vgnd vpwr scs8hd_decap_12
XFILLER_35_355 vgnd vpwr scs8hd_decap_4
XFILLER_35_344 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ bottom_width_0_height_0__pin_31_ vgnd vpwr scs8hd_diode_2
XFILLER_50_369 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _34_/HI vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_196 vgnd vpwr scs8hd_decap_12
XFILLER_41_358 vpwr vgnd scs8hd_fill_2
XFILLER_41_325 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_44_141 vgnd vpwr scs8hd_decap_12
XFILLER_32_358 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_406 vgnd vpwr scs8hd_fill_1
XFILLER_27_119 vgnd vpwr scs8hd_decap_3
XFILLER_50_166 vgnd vpwr scs8hd_decap_12
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_358 vpwr vgnd scs8hd_fill_2
XFILLER_46_406 vgnd vpwr scs8hd_fill_1
XFILLER_58_288 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ right_width_0_height_0__pin_6_ vgnd vpwr scs8hd_diode_2
XFILLER_26_152 vgnd vpwr scs8hd_fill_1
XPHY_42 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_75 vpwr vgnd scs8hd_fill_2
XFILLER_22_380 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_49_288 vgnd vpwr scs8hd_decap_3
X_51_ _51_/HI _51_/LO vgnd vpwr scs8hd_conb_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_1_295 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_28_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_55_269 vgnd vpwr scs8hd_decap_12
XFILLER_23_177 vpwr vgnd scs8hd_fill_2
XFILLER_11_306 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_46_258 vgnd vpwr scs8hd_decap_12
XFILLER_46_247 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_361 vgnd vpwr scs8hd_decap_12
XFILLER_6_398 vgnd vpwr scs8hd_decap_8
XFILLER_52_239 vgnd vpwr scs8hd_decap_12
XFILLER_45_280 vpwr vgnd scs8hd_fill_2
X_34_ _34_/HI _34_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ bottom_width_0_height_0__pin_22_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_125 vgnd vpwr scs8hd_fill_1
XFILLER_9_170 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_247 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_250 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XPHY_459 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_448 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_437 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_426 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_415 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_404 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_114 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_98 vgnd vpwr scs8hd_decap_12
XFILLER_22_32 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_158 vpwr vgnd scs8hd_fill_2
XFILLER_3_335 vpwr vgnd scs8hd_fill_2
XFILLER_47_62 vgnd vpwr scs8hd_decap_12
XFILLER_47_51 vgnd vpwr scs8hd_decap_8
XFILLER_34_206 vgnd vpwr scs8hd_decap_8
XFILLER_19_203 vpwr vgnd scs8hd_fill_2
XFILLER_8_78 vpwr vgnd scs8hd_fill_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_390 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1_0_clk/X ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ bottom_width_0_height_0__pin_50_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XFILLER_18_280 vpwr vgnd scs8hd_fill_2
XFILLER_33_283 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_342 vpwr vgnd scs8hd_fill_2
XFILLER_17_54 vgnd vpwr scs8hd_fill_1
XFILLER_16_239 vpwr vgnd scs8hd_fill_2
XFILLER_16_228 vgnd vpwr scs8hd_decap_4
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XPHY_289 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_132 vgnd vpwr scs8hd_decap_3
XFILLER_3_110 vpwr vgnd scs8hd_fill_2
XFILLER_62_389 vgnd vpwr scs8hd_decap_8
XFILLER_62_312 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_220 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_301 vgnd vpwr scs8hd_decap_4
XFILLER_38_364 vpwr vgnd scs8hd_fill_2
XFILLER_53_378 vpwr vgnd scs8hd_fill_2
XFILLER_53_367 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_297 vpwr vgnd scs8hd_fill_2
XFILLER_48_117 vgnd vpwr scs8hd_decap_12
XFILLER_0_113 vpwr vgnd scs8hd_fill_2
XFILLER_0_179 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_323 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_253 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_35_312 vpwr vgnd scs8hd_fill_2
XFILLER_50_337 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_367 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_356 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_205 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XFILLER_29_161 vpwr vgnd scs8hd_fill_2
XFILLER_17_301 vpwr vgnd scs8hd_fill_2
XFILLER_55_62 vgnd vpwr scs8hd_decap_12
XFILLER_55_51 vgnd vpwr scs8hd_decap_8
XFILLER_32_337 vpwr vgnd scs8hd_fill_2
XFILLER_40_381 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_271 vpwr vgnd scs8hd_fill_2
XFILLER_23_304 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_178 vgnd vpwr scs8hd_decap_12
XFILLER_23_348 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_98 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_decap_3
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_54 vpwr vgnd scs8hd_fill_2
XPHY_43 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XFILLER_14_337 vpwr vgnd scs8hd_fill_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_49_267 vpwr vgnd scs8hd_fill_2
XFILLER_49_245 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_17_153 vgnd vpwr scs8hd_decap_12
XFILLER_2_69 vpwr vgnd scs8hd_fill_2
X_50_ _50_/HI _50_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_329 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_175 vpwr vgnd scs8hd_fill_2
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_63_281 vgnd vpwr scs8hd_decap_12
XFILLER_23_123 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_11_318 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ right_width_0_height_0__pin_0_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _38_/HI vgnd vpwr scs8hd_diode_2
XFILLER_11_89 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_46_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _44_/HI
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_47_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_145 vpwr vgnd scs8hd_fill_2
XFILLER_6_366 vgnd vpwr scs8hd_decap_12
XFILLER_10_373 vgnd vpwr scs8hd_decap_12
X_33_ _33_/HI _33_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ bottom_width_0_height_0__pin_21_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_60_251 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_215 vgnd vpwr scs8hd_decap_3
XFILLER_51_284 vgnd vpwr scs8hd_decap_3
XPHY_449 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_438 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_427 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_416 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_405 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_108 vgnd vpwr scs8hd_decap_12
XFILLER_59_362 vpwr vgnd scs8hd_fill_2
XFILLER_3_358 vpwr vgnd scs8hd_fill_2
XFILLER_63_51 vgnd vpwr scs8hd_decap_8
XFILLER_47_74 vgnd vpwr scs8hd_decap_12
XFILLER_63_62 vgnd vpwr scs8hd_decap_12
XFILLER_42_295 vpwr vgnd scs8hd_fill_2
XFILLER_6_163 vpwr vgnd scs8hd_fill_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_207 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_306 vpwr vgnd scs8hd_fill_2
XFILLER_56_398 vgnd vpwr scs8hd_decap_8
XFILLER_17_77 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XFILLER_24_295 vgnd vpwr scs8hd_decap_12
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_406 vgnd vpwr scs8hd_fill_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_166 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_62_324 vgnd vpwr scs8hd_decap_12
XFILLER_47_376 vpwr vgnd scs8hd_fill_2
XFILLER_30_210 vgnd vpwr scs8hd_fill_1
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
XFILLER_30_276 vpwr vgnd scs8hd_fill_2
XFILLER_30_232 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_357 vgnd vpwr scs8hd_decap_3
XFILLER_38_398 vgnd vpwr scs8hd_decap_8
XFILLER_38_387 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_276 vpwr vgnd scs8hd_fill_2
XFILLER_21_221 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_129 vgnd vpwr scs8hd_decap_12
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_125 vgnd vpwr scs8hd_decap_3
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_44_379 vgnd vpwr scs8hd_decap_12
XFILLER_44_302 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _48_/HI vgnd vpwr scs8hd_diode_2
XFILLER_8_258 vgnd vpwr scs8hd_decap_4
XFILLER_12_276 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_184 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_62_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_217 vpwr vgnd scs8hd_fill_2
XFILLER_14_78 vgnd vpwr scs8hd_decap_12
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_17_335 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_74 vgnd vpwr scs8hd_decap_12
XFILLER_44_154 vgnd vpwr scs8hd_decap_12
XFILLER_32_327 vpwr vgnd scs8hd_fill_2
XFILLER_32_316 vpwr vgnd scs8hd_fill_2
XFILLER_32_305 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_40_393 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_250 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XFILLER_31_382 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_209 vgnd vpwr scs8hd_decap_3
XFILLER_58_202 vgnd vpwr scs8hd_decap_12
XPHY_99 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_88 vgnd vpwr scs8hd_decap_3
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vpwr vgnd scs8hd_fill_2
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ bottom_width_0_height_0__pin_28_ vgnd vpwr scs8hd_diode_2
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_264 vpwr vgnd scs8hd_fill_2
XFILLER_64_249 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_17_165 vgnd vpwr scs8hd_decap_4
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XFILLER_32_168 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_63_293 vgnd vpwr scs8hd_decap_12
XFILLER_48_290 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_61_208 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_46_227 vgnd vpwr scs8hd_decap_12
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_14_168 vgnd vpwr scs8hd_decap_3
XFILLER_6_356 vgnd vpwr scs8hd_fill_1
XFILLER_6_378 vgnd vpwr scs8hd_decap_12
XFILLER_10_385 vgnd vpwr scs8hd_decap_12
X_32_ _32_/HI _32_/LO vgnd vpwr scs8hd_conb_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ bottom_width_0_height_0__pin_20_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_60_263 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_149 vgnd vpwr scs8hd_decap_4
XFILLER_20_116 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_208 vgnd vpwr scs8hd_decap_12
XFILLER_28_227 vgnd vpwr scs8hd_decap_8
XFILLER_51_296 vpwr vgnd scs8hd_fill_2
XPHY_439 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_428 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_417 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_406 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_315 vpwr vgnd scs8hd_fill_2
XFILLER_59_341 vpwr vgnd scs8hd_fill_2
XFILLER_19_238 vgnd vpwr scs8hd_decap_6
XFILLER_63_74 vgnd vpwr scs8hd_decap_12
XFILLER_47_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_175 vpwr vgnd scs8hd_fill_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_296 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_56_300 vgnd vpwr scs8hd_decap_8
XFILLER_56_333 vgnd vpwr scs8hd_fill_1
XFILLER_17_23 vpwr vgnd scs8hd_fill_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _42_/HI vgnd vpwr scs8hd_diode_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_3_178 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_171 vgnd vpwr scs8hd_decap_12
XFILLER_47_388 vpwr vgnd scs8hd_fill_2
XFILLER_47_355 vpwr vgnd scs8hd_fill_2
XFILLER_47_344 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _59_/HI vgnd vpwr scs8hd_diode_2
XFILLER_30_244 vpwr vgnd scs8hd_fill_2
XFILLER_15_296 vpwr vgnd scs8hd_fill_2
XFILLER_30_288 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _53_/HI
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_34_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_56_141 vgnd vpwr scs8hd_decap_12
XFILLER_29_333 vpwr vgnd scs8hd_fill_2
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_204 vpwr vgnd scs8hd_fill_2
XFILLER_8_237 vpwr vgnd scs8hd_fill_2
XFILLER_12_288 vgnd vpwr scs8hd_decap_4
XFILLER_62_166 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ right_width_0_height_0__pin_10_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_47_196 vgnd vpwr scs8hd_decap_12
XFILLER_7_281 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_406 vgnd vpwr scs8hd_fill_1
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_41_306 vpwr vgnd scs8hd_fill_2
XFILLER_34_391 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_49_406 vgnd vpwr scs8hd_fill_1
XFILLER_55_86 vgnd vpwr scs8hd_decap_12
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_17_358 vpwr vgnd scs8hd_fill_2
XFILLER_17_325 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_44_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_391 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_240 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_295 vpwr vgnd scs8hd_fill_2
XFILLER_23_317 vpwr vgnd scs8hd_fill_2
XFILLER_23_306 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_394 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_23 vgnd vpwr scs8hd_decap_3
XFILLER_2_38 vpwr vgnd scs8hd_fill_2
XFILLER_2_27 vpwr vgnd scs8hd_fill_2
XFILLER_1_287 vpwr vgnd scs8hd_fill_2
XFILLER_1_243 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_188 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_9_365 vgnd vpwr scs8hd_fill_1
XFILLER_49_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_136 vpwr vgnd scs8hd_fill_2
XFILLER_23_103 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_294 vgnd vpwr scs8hd_fill_1
XFILLER_46_239 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_125 vgnd vpwr scs8hd_fill_1
XFILLER_52_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0_0_clk/X ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XFILLER_6_302 vgnd vpwr scs8hd_decap_3
XFILLER_6_324 vpwr vgnd scs8hd_fill_2
XFILLER_10_331 vgnd vpwr scs8hd_decap_4
XFILLER_6_346 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_162 vgnd vpwr scs8hd_decap_8
XFILLER_9_184 vgnd vpwr scs8hd_decap_3
XFILLER_3_92 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_51_220 vgnd vpwr scs8hd_decap_12
XPHY_407 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_261 vpwr vgnd scs8hd_fill_2
XFILLER_36_250 vpwr vgnd scs8hd_fill_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_6
XFILLER_28_206 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XPHY_429 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_418 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_386 vgnd vpwr scs8hd_decap_8
XFILLER_47_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_294 vpwr vgnd scs8hd_fill_2
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_110 vgnd vpwr scs8hd_decap_4
XFILLER_6_132 vpwr vgnd scs8hd_fill_2
XFILLER_2_382 vpwr vgnd scs8hd_fill_2
XFILLER_33_253 vgnd vpwr scs8hd_decap_4
XFILLER_21_404 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_389 vgnd vpwr scs8hd_decap_8
XFILLER_56_367 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_337 vgnd vpwr scs8hd_decap_12
XFILLER_47_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_264 vgnd vpwr scs8hd_decap_12
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_61_381 vgnd vpwr scs8hd_decap_12
XFILLER_53_326 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_289 vgnd vpwr scs8hd_decap_8
XFILLER_21_245 vgnd vpwr scs8hd_decap_12
XFILLER_44_337 vgnd vpwr scs8hd_decap_4
XFILLER_29_367 vgnd vpwr scs8hd_decap_12
XFILLER_29_356 vpwr vgnd scs8hd_fill_2
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XFILLER_52_381 vgnd vpwr scs8hd_decap_12
XFILLER_44_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ right_width_0_height_0__pin_9_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_62_178 vgnd vpwr scs8hd_decap_12
XFILLER_35_359 vgnd vpwr scs8hd_fill_1
XFILLER_35_348 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_293 vpwr vgnd scs8hd_fill_2
XFILLER_53_123 vgnd vpwr scs8hd_decap_12
XFILLER_41_329 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ bottom_width_0_height_0__pin_25_ vgnd vpwr scs8hd_diode_2
XFILLER_14_36 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_98 vgnd vpwr scs8hd_decap_12
XFILLER_44_178 vgnd vpwr scs8hd_decap_12
XFILLER_29_175 vpwr vgnd scs8hd_fill_2
XFILLER_17_348 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _46_/HI vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _42_/HI
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XFILLER_31_362 vpwr vgnd scs8hd_fill_2
XFILLER_58_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_81 vgnd vpwr scs8hd_decap_8
XFILLER_26_189 vpwr vgnd scs8hd_fill_2
XFILLER_26_112 vgnd vpwr scs8hd_decap_12
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_79 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_64_218 vgnd vpwr scs8hd_decap_12
XFILLER_57_281 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_17_112 vpwr vgnd scs8hd_fill_2
XFILLER_1_299 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_270 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _54_/HI
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_23_115 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_54_251 vgnd vpwr scs8hd_decap_12
XFILLER_39_281 vgnd vpwr scs8hd_fill_1
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_44 vgnd vpwr scs8hd_decap_12
XFILLER_22_181 vgnd vpwr scs8hd_decap_12
XFILLER_10_398 vgnd vpwr scs8hd_decap_8
XFILLER_45_240 vpwr vgnd scs8hd_fill_2
XFILLER_33_402 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_60_276 vgnd vpwr scs8hd_decap_12
XFILLER_45_284 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_71 vpwr vgnd scs8hd_fill_2
XFILLER_51_232 vgnd vpwr scs8hd_decap_12
XPHY_419 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_408 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_295 vgnd vpwr scs8hd_decap_3
XFILLER_36_273 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_7 vpwr vgnd scs8hd_fill_2
XFILLER_59_398 vpwr vgnd scs8hd_fill_2
XFILLER_59_354 vpwr vgnd scs8hd_fill_2
XFILLER_27_240 vpwr vgnd scs8hd_fill_2
XFILLER_19_207 vpwr vgnd scs8hd_fill_2
XFILLER_63_98 vgnd vpwr scs8hd_decap_12
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_173 vpwr vgnd scs8hd_fill_2
XFILLER_10_195 vpwr vgnd scs8hd_fill_2
XFILLER_12_91 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_284 vpwr vgnd scs8hd_fill_2
XFILLER_18_273 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_346 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_58_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ bottom_width_0_height_0__pin_19_ vgnd vpwr scs8hd_diode_2
XFILLER_62_349 vgnd vpwr scs8hd_decap_12
XFILLER_59_184 vgnd vpwr scs8hd_decap_12
XFILLER_55_390 vpwr vgnd scs8hd_fill_2
XFILLER_15_221 vgnd vpwr scs8hd_decap_4
XFILLER_30_224 vpwr vgnd scs8hd_fill_2
XFILLER_30_213 vgnd vpwr scs8hd_fill_1
XFILLER_15_276 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_335 vgnd vpwr scs8hd_fill_1
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_61_393 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_257 vgnd vpwr scs8hd_decap_6
XFILLER_9_70 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_117 vgnd vpwr scs8hd_decap_4
XFILLER_56_154 vgnd vpwr scs8hd_decap_12
XFILLER_29_379 vgnd vpwr scs8hd_decap_12
XFILLER_29_346 vgnd vpwr scs8hd_decap_4
XFILLER_28_79 vgnd vpwr scs8hd_fill_1
XFILLER_28_68 vgnd vpwr scs8hd_decap_3
XFILLER_60_44 vgnd vpwr scs8hd_decap_12
XFILLER_52_393 vgnd vpwr scs8hd_decap_4
XFILLER_44_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_202 vpwr vgnd scs8hd_fill_2
XFILLER_12_224 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ right_width_0_height_0__pin_8_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_371 vgnd vpwr scs8hd_decap_3
XFILLER_35_316 vpwr vgnd scs8hd_fill_2
XFILLER_53_135 vgnd vpwr scs8hd_decap_12
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_404 vgnd vpwr scs8hd_decap_3
XFILLER_5_209 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_308 vgnd vpwr scs8hd_decap_3
XFILLER_29_165 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_52_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
XFILLER_50_105 vgnd vpwr scs8hd_decap_12
XFILLER_31_341 vpwr vgnd scs8hd_fill_2
XFILLER_31_330 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_16_360 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
XFILLER_58_227 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_168 vpwr vgnd scs8hd_fill_2
XFILLER_26_124 vgnd vpwr scs8hd_decap_12
XFILLER_25_58 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XFILLER_14_308 vpwr vgnd scs8hd_fill_2
XFILLER_14_319 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XFILLER_22_363 vpwr vgnd scs8hd_fill_2
XFILLER_22_352 vpwr vgnd scs8hd_fill_2
XFILLER_1_245 vpwr vgnd scs8hd_fill_2
XFILLER_57_293 vgnd vpwr scs8hd_decap_12
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_17_179 vgnd vpwr scs8hd_decap_4
XFILLER_13_352 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_367 vgnd vpwr scs8hd_decap_12
XFILLER_55_208 vgnd vpwr scs8hd_decap_12
XFILLER_23_149 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
XFILLER_54_263 vgnd vpwr scs8hd_decap_12
XFILLER_52_56 vgnd vpwr scs8hd_decap_12
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_14_149 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_193 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_6_337 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _50_/HI vgnd vpwr scs8hd_diode_2
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_60_288 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_131 vpwr vgnd scs8hd_fill_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_193 vgnd vpwr scs8hd_decap_4
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_370 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_409 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _33_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_285 vgnd vpwr scs8hd_decap_3
XFILLER_27_263 vgnd vpwr scs8hd_fill_1
XFILLER_42_299 vpwr vgnd scs8hd_fill_2
XFILLER_30_406 vgnd vpwr scs8hd_fill_1
XFILLER_10_130 vpwr vgnd scs8hd_fill_2
XFILLER_10_141 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ top_width_0_height_0__pin_32_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
XFILLER_6_167 vgnd vpwr scs8hd_decap_3
XFILLER_10_185 vgnd vpwr scs8hd_decap_8
XFILLER_18_230 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_24_211 vgnd vpwr scs8hd_fill_1
XFILLER_17_15 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_406 vgnd vpwr scs8hd_fill_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_3_137 vgnd vpwr scs8hd_decap_4
XFILLER_59_196 vgnd vpwr scs8hd_decap_12
XFILLER_58_44 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1_0_clk/X ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _33_/HI
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_40_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_91 vgnd vpwr scs8hd_decap_12
XFILLER_15_288 vgnd vpwr scs8hd_decap_6
XFILLER_53_339 vgnd vpwr scs8hd_decap_3
XFILLER_53_306 vgnd vpwr scs8hd_decap_12
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_269 vgnd vpwr scs8hd_decap_4
XFILLER_21_225 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ bottom_width_0_height_0__pin_22_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_166 vgnd vpwr scs8hd_decap_12
XFILLER_44_306 vpwr vgnd scs8hd_fill_2
XFILLER_44_68 vgnd vpwr scs8hd_decap_12
XFILLER_37_380 vpwr vgnd scs8hd_fill_2
XFILLER_60_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_306 vgnd vpwr scs8hd_decap_4
XFILLER_43_383 vpwr vgnd scs8hd_fill_2
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XFILLER_53_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XFILLER_26_328 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _43_/HI ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_111 vgnd vpwr scs8hd_decap_8
XFILLER_4_210 vpwr vgnd scs8hd_fill_2
XFILLER_4_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
XFILLER_29_90 vgnd vpwr scs8hd_decap_3
XFILLER_50_117 vgnd vpwr scs8hd_decap_12
XFILLER_16_383 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_58_239 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0_0_clk/X ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_158 vgnd vpwr scs8hd_decap_8
XFILLER_26_136 vgnd vpwr scs8hd_decap_12
XFILLER_25_37 vpwr vgnd scs8hd_fill_2
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_235 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_302 vgnd vpwr scs8hd_decap_3
XFILLER_13_320 vgnd vpwr scs8hd_decap_12
XFILLER_13_364 vpwr vgnd scs8hd_fill_2
XFILLER_13_375 vgnd vpwr scs8hd_decap_12
XFILLER_9_379 vgnd vpwr scs8hd_decap_12
XFILLER_63_220 vgnd vpwr scs8hd_decap_12
XFILLER_51_404 vgnd vpwr scs8hd_decap_3
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
XFILLER_39_261 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_68 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_45_297 vpwr vgnd scs8hd_fill_2
XFILLER_45_264 vpwr vgnd scs8hd_fill_2
XFILLER_45_220 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_47_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_382 vgnd vpwr scs8hd_decap_12
XFILLER_51_256 vpwr vgnd scs8hd_fill_2
XFILLER_51_245 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_319 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_245 vgnd vpwr scs8hd_fill_1
XFILLER_42_267 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _59_/HI ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_6_179 vpwr vgnd scs8hd_fill_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_396 vgnd vpwr scs8hd_fill_1
XFILLER_33_223 vpwr vgnd scs8hd_fill_2
XFILLER_33_201 vgnd vpwr scs8hd_fill_1
XFILLER_18_253 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_337 vgnd vpwr scs8hd_decap_3
XFILLER_17_27 vpwr vgnd scs8hd_fill_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ top_width_0_height_0__pin_32_ vgnd vpwr scs8hd_diode_2
XFILLER_24_267 vgnd vpwr scs8hd_decap_6
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_3_105 vgnd vpwr scs8hd_decap_3
XFILLER_58_56 vgnd vpwr scs8hd_decap_12
XFILLER_47_359 vgnd vpwr scs8hd_decap_4
XFILLER_47_348 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_30_248 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_318 vgnd vpwr scs8hd_decap_6
XFILLER_38_359 vgnd vpwr scs8hd_decap_3
XFILLER_38_337 vgnd vpwr scs8hd_decap_12
XFILLER_0_41 vpwr vgnd scs8hd_fill_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_3
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_61_351 vgnd vpwr scs8hd_decap_12
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_56_178 vgnd vpwr scs8hd_decap_12
XFILLER_52_373 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _60_/HI vgnd vpwr scs8hd_diode_2
XFILLER_8_208 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_123 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_560 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_362 vpwr vgnd scs8hd_fill_2
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XFILLER_7_285 vpwr vgnd scs8hd_fill_2
XFILLER_11_270 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ bottom_width_0_height_0__pin_16_ vgnd vpwr scs8hd_diode_2
XFILLER_53_159 vgnd vpwr scs8hd_decap_12
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XFILLER_25_351 vgnd vpwr scs8hd_decap_12
XFILLER_40_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_93 vpwr vgnd scs8hd_fill_2
XFILLER_4_299 vpwr vgnd scs8hd_fill_2
XFILLER_50_129 vgnd vpwr scs8hd_decap_12
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XPHY_390 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_395 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ bottom_width_0_height_0__pin_23_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_or2_1
XFILLER_6_73 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_148 vgnd vpwr scs8hd_decap_4
XFILLER_25_27 vgnd vpwr scs8hd_decap_8
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_22_376 vpwr vgnd scs8hd_fill_2
XFILLER_22_332 vpwr vgnd scs8hd_fill_2
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_398 vgnd vpwr scs8hd_decap_8
XFILLER_1_203 vpwr vgnd scs8hd_fill_2
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_325 vgnd vpwr scs8hd_decap_12
XFILLER_13_332 vgnd vpwr scs8hd_decap_12
XFILLER_13_387 vgnd vpwr scs8hd_decap_12
XFILLER_48_262 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_63_232 vgnd vpwr scs8hd_decap_12
XFILLER_31_162 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_276 vgnd vpwr scs8hd_decap_12
XFILLER_39_284 vpwr vgnd scs8hd_fill_2
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_335 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_328 vgnd vpwr scs8hd_decap_6
XFILLER_60_202 vgnd vpwr scs8hd_decap_12
XFILLER_45_276 vpwr vgnd scs8hd_fill_2
XFILLER_45_232 vgnd vpwr scs8hd_decap_6
XFILLER_42_80 vgnd vpwr scs8hd_decap_12
XFILLER_13_162 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_30 vpwr vgnd scs8hd_fill_2
XFILLER_5_394 vgnd vpwr scs8hd_decap_12
XFILLER_36_265 vpwr vgnd scs8hd_fill_2
XFILLER_51_279 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_202 vgnd vpwr scs8hd_decap_12
XFILLER_27_298 vpwr vgnd scs8hd_fill_2
XFILLER_27_254 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_405 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_2_386 vpwr vgnd scs8hd_fill_2
XFILLER_2_320 vpwr vgnd scs8hd_fill_2
XFILLER_12_83 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_18_265 vgnd vpwr scs8hd_decap_8
XFILLER_18_276 vpwr vgnd scs8hd_fill_2
XFILLER_41_290 vgnd vpwr scs8hd_fill_1
XFILLER_33_279 vpwr vgnd scs8hd_fill_2
XFILLER_33_257 vgnd vpwr scs8hd_fill_1
XFILLER_33_235 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_327 vgnd vpwr scs8hd_decap_6
XFILLER_49_390 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_24_246 vpwr vgnd scs8hd_fill_2
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_59_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_58_68 vgnd vpwr scs8hd_decap_12
XFILLER_55_382 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_15_213 vpwr vgnd scs8hd_fill_2
XFILLER_38_327 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_61_363 vgnd vpwr scs8hd_decap_3
XFILLER_61_330 vgnd vpwr scs8hd_decap_12
XFILLER_38_349 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_205 vgnd vpwr scs8hd_decap_12
XFILLER_9_40 vpwr vgnd scs8hd_fill_2
XFILLER_9_62 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_44_319 vpwr vgnd scs8hd_fill_2
XFILLER_29_316 vpwr vgnd scs8hd_fill_2
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_44_15 vgnd vpwr scs8hd_decap_12
XFILLER_37_393 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_105 vgnd vpwr scs8hd_decap_12
XFILLER_47_135 vgnd vpwr scs8hd_decap_12
XFILLER_43_341 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_561 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_550 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_80 vgnd vpwr scs8hd_decap_12
XFILLER_7_264 vpwr vgnd scs8hd_fill_2
XFILLER_7_297 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_61_171 vgnd vpwr scs8hd_decap_12
XFILLER_46_190 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XFILLER_29_157 vpwr vgnd scs8hd_fill_2
XFILLER_29_135 vgnd vpwr scs8hd_decap_12
XFILLER_40_377 vpwr vgnd scs8hd_fill_2
XFILLER_40_333 vgnd vpwr scs8hd_decap_3
XFILLER_25_363 vgnd vpwr scs8hd_decap_3
XFILLER_4_234 vgnd vpwr scs8hd_decap_4
XFILLER_4_267 vpwr vgnd scs8hd_fill_2
XFILLER_63_403 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_43_171 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_391 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_380 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_clkbuf_1_1_0_clk_A clkbuf_0_clk/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_22_311 vgnd vpwr scs8hd_decap_6
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_49_208 vgnd vpwr scs8hd_decap_12
XFILLER_60_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_149 vpwr vgnd scs8hd_fill_2
XFILLER_17_127 vgnd vpwr scs8hd_fill_1
XFILLER_17_116 vgnd vpwr scs8hd_decap_4
XFILLER_17_105 vgnd vpwr scs8hd_decap_4
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XANTENNA__71__A bottom_width_0_height_0__pin_49_lower vgnd vpwr scs8hd_diode_2
XFILLER_9_337 vgnd vpwr scs8hd_decap_12
XFILLER_13_344 vpwr vgnd scs8hd_fill_2
XFILLER_13_399 vgnd vpwr scs8hd_decap_8
XFILLER_48_285 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_288 vgnd vpwr scs8hd_decap_6
XFILLER_52_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_406 vgnd vpwr scs8hd_fill_1
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA__66__A bottom_width_0_height_0__pin_44_lower vgnd vpwr scs8hd_diode_2
XFILLER_33_406 vgnd vpwr scs8hd_fill_1
XFILLER_26_71 vpwr vgnd scs8hd_fill_2
XFILLER_9_101 vpwr vgnd scs8hd_fill_2
XFILLER_13_141 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _56_/HI
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_37_lower vgnd vpwr scs8hd_mux2_1
XFILLER_5_351 vpwr vgnd scs8hd_fill_2
XFILLER_9_189 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_75 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XFILLER_36_244 vgnd vpwr scs8hd_decap_4
XFILLER_36_222 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_406 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0_0_clk/X ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _47_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_59_358 vpwr vgnd scs8hd_fill_2
XFILLER_59_314 vpwr vgnd scs8hd_fill_2
XFILLER_47_59 vpwr vgnd scs8hd_fill_2
XFILLER_47_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_233 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_10_122 vgnd vpwr scs8hd_fill_1
XFILLER_10_177 vgnd vpwr scs8hd_decap_4
XFILLER_2_398 vgnd vpwr scs8hd_decap_8
XFILLER_2_365 vpwr vgnd scs8hd_fill_2
XFILLER_2_332 vpwr vgnd scs8hd_fill_2
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_170 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XFILLER_24_236 vgnd vpwr scs8hd_decap_8
XFILLER_24_203 vgnd vpwr scs8hd_decap_8
X_69_ bottom_width_0_height_0__pin_47_lower bottom_width_0_height_0__pin_47_upper
+ vgnd vpwr scs8hd_buf_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _45_/HI
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_46_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_55_394 vgnd vpwr scs8hd_decap_12
XFILLER_55_350 vpwr vgnd scs8hd_fill_2
XFILLER_47_328 vgnd vpwr scs8hd_decap_8
XFILLER_47_306 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_15_203 vgnd vpwr scs8hd_decap_8
XFILLER_30_206 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _49_/HI vgnd vpwr scs8hd_diode_2
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ right_width_0_height_0__pin_13_ vgnd vpwr scs8hd_diode_2
XFILLER_38_317 vgnd vpwr scs8hd_decap_8
XFILLER_2_173 vpwr vgnd scs8hd_fill_2
XFILLER_61_342 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_217 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_0_32 vgnd vpwr scs8hd_fill_1
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_74 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_306 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_180 vgnd vpwr scs8hd_decap_6
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XFILLER_52_342 vpwr vgnd scs8hd_fill_2
XFILLER_44_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_206 vgnd vpwr scs8hd_decap_8
XFILLER_12_228 vgnd vpwr scs8hd_decap_6
XFILLER_62_117 vgnd vpwr scs8hd_decap_12
XANTENNA__74__A right_width_0_height_0__pin_35_lower vgnd vpwr scs8hd_diode_2
XFILLER_47_147 vgnd vpwr scs8hd_decap_12
XFILLER_28_372 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0_0_clk/X ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XPHY_562 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_551 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_540 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_210 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_34_375 vpwr vgnd scs8hd_fill_2
XFILLER_34_331 vpwr vgnd scs8hd_fill_2
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_55_59 vpwr vgnd scs8hd_fill_2
XFILLER_55_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_147 vgnd vpwr scs8hd_decap_8
XFILLER_25_320 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA__69__A bottom_width_0_height_0__pin_47_lower vgnd vpwr scs8hd_diode_2
XFILLER_4_246 vpwr vgnd scs8hd_fill_2
XPHY_370 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_378 vpwr vgnd scs8hd_fill_2
XFILLER_31_367 vpwr vgnd scs8hd_fill_2
XFILLER_31_345 vpwr vgnd scs8hd_fill_2
XFILLER_31_334 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XPHY_392 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_381 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_64 vpwr vgnd scs8hd_fill_2
XFILLER_6_97 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_22_389 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_249 vpwr vgnd scs8hd_fill_2
XFILLER_57_220 vgnd vpwr scs8hd_decap_12
XFILLER_45_404 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_312 vpwr vgnd scs8hd_fill_2
XFILLER_13_367 vgnd vpwr scs8hd_decap_6
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_349 vgnd vpwr scs8hd_decap_12
XFILLER_15_95 vpwr vgnd scs8hd_fill_2
XFILLER_0_271 vpwr vgnd scs8hd_fill_2
XFILLER_63_245 vgnd vpwr scs8hd_decap_12
XFILLER_56_80 vgnd vpwr scs8hd_decap_12
XFILLER_48_297 vgnd vpwr scs8hd_decap_6
XFILLER_31_175 vgnd vpwr scs8hd_decap_6
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
XFILLER_39_220 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_297 vpwr vgnd scs8hd_fill_2
XFILLER_22_142 vpwr vgnd scs8hd_fill_2
XFILLER_14_109 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_10_337 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_60_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_135 vpwr vgnd scs8hd_fill_2
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_197 vgnd vpwr scs8hd_fill_1
XFILLER_42_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_363 vgnd vpwr scs8hd_decap_3
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ right_width_0_height_0__pin_7_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_337 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XFILLER_47_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_59 vpwr vgnd scs8hd_fill_2
XFILLER_42_215 vgnd vpwr scs8hd_decap_12
XFILLER_10_134 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
XANTENNA__77__A right_width_0_height_0__pin_38_lower vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ right_width_0_height_0__pin_11_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_or2_1
XFILLER_5_193 vpwr vgnd scs8hd_fill_2
X_68_ bottom_width_0_height_0__pin_46_lower bottom_width_0_height_0__pin_46_upper
+ vgnd vpwr scs8hd_buf_2
XFILLER_64_373 vgnd vpwr scs8hd_decap_12
XFILLER_24_215 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_59_123 vgnd vpwr scs8hd_decap_12
XFILLER_58_15 vgnd vpwr scs8hd_decap_12
XFILLER_55_362 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_62 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_403 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_152 vgnd vpwr scs8hd_fill_1
XFILLER_2_141 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_11 vpwr vgnd scs8hd_fill_2
XFILLER_21_229 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_97 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_37_362 vpwr vgnd scs8hd_fill_2
XFILLER_29_329 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
XFILLER_52_398 vgnd vpwr scs8hd_decap_8
XFILLER_20_295 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ccff_tail
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_406 vgnd vpwr scs8hd_fill_1
XFILLER_47_159 vgnd vpwr scs8hd_decap_12
XPHY_552 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_541 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_129 vgnd vpwr scs8hd_decap_12
XPHY_530 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_387 vgnd vpwr scs8hd_decap_12
XFILLER_43_376 vgnd vpwr scs8hd_decap_3
XFILLER_43_354 vpwr vgnd scs8hd_fill_2
XFILLER_43_332 vgnd vpwr scs8hd_decap_3
XFILLER_43_310 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
XFILLER_18_73 vpwr vgnd scs8hd_fill_2
XPHY_563 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_222 vpwr vgnd scs8hd_fill_2
XFILLER_11_240 vgnd vpwr scs8hd_decap_4
XFILLER_34_321 vpwr vgnd scs8hd_fill_2
XFILLER_19_362 vpwr vgnd scs8hd_fill_2
XFILLER_19_351 vpwr vgnd scs8hd_fill_2
XFILLER_19_340 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_61_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_398 vgnd vpwr scs8hd_decap_8
XFILLER_34_354 vpwr vgnd scs8hd_fill_2
XFILLER_57_402 vgnd vpwr scs8hd_decap_4
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
XFILLER_55_27 vgnd vpwr scs8hd_decap_12
XFILLER_44_129 vgnd vpwr scs8hd_decap_12
XFILLER_40_313 vpwr vgnd scs8hd_fill_2
XFILLER_25_343 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_357 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_16_321 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _44_/HI vgnd vpwr scs8hd_diode_2
XFILLER_43_184 vgnd vpwr scs8hd_decap_12
XPHY_393 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_382 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_371 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_360 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_398 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_32 vpwr vgnd scs8hd_fill_2
XFILLER_19_170 vgnd vpwr scs8hd_decap_8
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_30_390 vgnd vpwr scs8hd_decap_6
XFILLER_22_346 vgnd vpwr scs8hd_decap_4
XFILLER_1_239 vpwr vgnd scs8hd_fill_2
XFILLER_57_232 vgnd vpwr scs8hd_decap_12
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_162 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_302 vgnd vpwr scs8hd_decap_3
XFILLER_15_52 vgnd vpwr scs8hd_decap_3
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_257 vgnd vpwr scs8hd_decap_12
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_361 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_54_202 vgnd vpwr scs8hd_decap_12
XFILLER_39_265 vgnd vpwr scs8hd_decap_12
XFILLER_39_232 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_22_110 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_198 vgnd vpwr scs8hd_decap_12
XFILLER_10_349 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_227 vgnd vpwr scs8hd_decap_12
XFILLER_45_268 vpwr vgnd scs8hd_fill_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_8
XFILLER_26_40 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_158 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_88 vpwr vgnd scs8hd_fill_2
XFILLER_44_290 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
XFILLER_47_39 vgnd vpwr scs8hd_decap_12
XFILLER_42_227 vgnd vpwr scs8hd_decap_12
XFILLER_27_213 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_271 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_106 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_128 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ right_width_0_height_0__pin_10_ vgnd vpwr scs8hd_diode_2
XFILLER_18_213 vgnd vpwr scs8hd_fill_1
XFILLER_33_249 vpwr vgnd scs8hd_fill_2
XFILLER_33_227 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_41_282 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_64_385 vgnd vpwr scs8hd_decap_12
X_67_ bottom_width_0_height_0__pin_45_lower bottom_width_0_height_0__pin_45_upper
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_293 vgnd vpwr scs8hd_decap_12
XFILLER_32_271 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_59_135 vgnd vpwr scs8hd_decap_12
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
XFILLER_55_330 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_23_282 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ bottom_width_0_height_0__pin_30_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_58_190 vgnd vpwr scs8hd_decap_12
XFILLER_48_93 vgnd vpwr scs8hd_decap_12
XFILLER_46_363 vgnd vpwr scs8hd_decap_4
XFILLER_46_341 vgnd vpwr scs8hd_decap_3
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_61_377 vpwr vgnd scs8hd_fill_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_260 vgnd vpwr scs8hd_decap_12
XFILLER_56_105 vgnd vpwr scs8hd_decap_12
XFILLER_37_352 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_564 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_553 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_542 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_531 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_520 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_55_171 vgnd vpwr scs8hd_decap_12
XFILLER_43_399 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_196 vgnd vpwr scs8hd_decap_12
XFILLER_55_39 vgnd vpwr scs8hd_decap_12
XFILLER_52_141 vgnd vpwr scs8hd_decap_12
XFILLER_40_325 vgnd vpwr scs8hd_decap_8
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_6
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_20_64 vpwr vgnd scs8hd_fill_2
XFILLER_29_95 vpwr vgnd scs8hd_fill_2
XFILLER_16_333 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_196 vgnd vpwr scs8hd_decap_12
XPHY_394 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_383 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_372 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_361 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_350 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_358 vpwr vgnd scs8hd_fill_2
XFILLER_31_303 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_54_406 vgnd vpwr scs8hd_fill_1
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _50_/HI
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ccff_tail
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XFILLER_22_358 vgnd vpwr scs8hd_decap_3
XFILLER_1_207 vpwr vgnd scs8hd_fill_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0_0_clk/X ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XFILLER_36_406 vgnd vpwr scs8hd_fill_1
XFILLER_0_262 vpwr vgnd scs8hd_fill_2
XFILLER_63_269 vgnd vpwr scs8hd_decap_12
XFILLER_56_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_373 vgnd vpwr scs8hd_decap_12
.ends

