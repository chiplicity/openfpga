* NGSPICE file created from cby_3__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

.subckt cby_3__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_grid_pin_1_ left_grid_pin_5_ left_grid_pin_9_ right_grid_pin_0_ right_grid_pin_10_
+ right_grid_pin_12_ right_grid_pin_14_ right_grid_pin_2_ right_grid_pin_4_ right_grid_pin_6_
+ right_grid_pin_8_ vpwr vgnd
XFILLER_26_52 vgnd vpwr scs8hd_decap_4
XFILLER_42_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_39 vgnd vpwr scs8hd_decap_12
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XFILLER_12_32 vgnd vpwr scs8hd_decap_3
XFILLER_12_76 vgnd vpwr scs8hd_decap_3
XFILLER_53_83 vgnd vpwr scs8hd_decap_3
XANTENNA__124__A _140_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_2_.latch/Q mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_ipin_6.LATCH_4_.latch/Q mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__209__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
X_200_ chany_top_in[0] chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _159_/Y vgnd vpwr
+ scs8hd_diode_2
X_131_ _139_/A _135_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__110__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_9_99 vpwr vgnd scs8hd_fill_2
XFILLER_9_77 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_4.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__119__A _137_/A vgnd vpwr scs8hd_diode_2
XFILLER_50_3 vgnd vpwr scs8hd_decap_12
XFILLER_62_109 vgnd vpwr scs8hd_fill_1
X_114_ _140_/A _116_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_59_93 vpwr vgnd scs8hd_fill_2
XANTENNA__121__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_128 vgnd vpwr scs8hd_decap_12
XFILLER_61_131 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_5.INVTX1_5_.scs8hd_inv_1 chany_top_in[5] mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_19 vpwr vgnd scs8hd_fill_2
XFILLER_29_106 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_2.LATCH_1_.latch data_in _161_/A _157_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_32 vgnd vpwr scs8hd_fill_1
XFILLER_29_41 vgnd vpwr scs8hd_fill_1
XFILLER_45_95 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_2.LATCH_1_.latch/Q mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__116__B _116_/B vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _140_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XFILLER_40_145 vgnd vpwr scs8hd_fill_1
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_31_75 vpwr vgnd scs8hd_fill_2
XFILLER_56_61 vpwr vgnd scs8hd_fill_2
XANTENNA__127__A _143_/A vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XFILLER_26_97 vgnd vpwr scs8hd_decap_4
XFILLER_42_85 vgnd vpwr scs8hd_fill_1
XFILLER_42_41 vpwr vgnd scs8hd_fill_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_7.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_6.LATCH_2_.latch/Q mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _186_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_104 vgnd vpwr scs8hd_decap_8
XFILLER_10_115 vgnd vpwr scs8hd_decap_12
XFILLER_12_55 vpwr vgnd scs8hd_fill_2
XFILLER_37_52 vpwr vgnd scs8hd_fill_2
XFILLER_53_95 vpwr vgnd scs8hd_fill_2
XFILLER_53_62 vpwr vgnd scs8hd_fill_2
XFILLER_53_51 vpwr vgnd scs8hd_fill_2
XFILLER_5_130 vgnd vpwr scs8hd_decap_12
XANTENNA__124__B _128_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _140_/A vgnd vpwr scs8hd_diode_2
XFILLER_59_126 vpwr vgnd scs8hd_fill_2
XFILLER_59_115 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_1.LATCH_5_.latch data_in mem_left_ipin_1.LATCH_5_.latch/Q _173_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_4.LATCH_0_.latch/Q mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_130_ _129_/X _135_/B vgnd vpwr scs8hd_buf_1
XFILLER_48_84 vgnd vpwr scs8hd_decap_8
XANTENNA__110__D _109_/Y vgnd vpwr scs8hd_diode_2
XFILLER_64_94 vgnd vpwr scs8hd_decap_12
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__119__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__135__A _143_/A vgnd vpwr scs8hd_diode_2
XFILLER_43_3 vgnd vpwr scs8hd_decap_12
XFILLER_56_107 vgnd vpwr scs8hd_decap_4
XFILLER_47_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_ipin_1.LATCH_3_.latch/Q mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_8
X_113_ _100_/B _140_/A vgnd vpwr scs8hd_buf_1
XFILLER_50_52 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_61_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_121 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_5.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_29_86 vpwr vgnd scs8hd_fill_2
XFILLER_43_143 vgnd vpwr scs8hd_decap_3
XFILLER_43_121 vgnd vpwr scs8hd_fill_1
XFILLER_61_95 vgnd vpwr scs8hd_decap_4
XFILLER_61_62 vgnd vpwr scs8hd_decap_3
XFILLER_61_51 vgnd vpwr scs8hd_decap_4
XANTENNA__132__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_121 vpwr vgnd scs8hd_fill_2
XFILLER_34_132 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_3.INVTX1_5_.scs8hd_inv_1 chany_top_in[7] mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_121 vgnd vpwr scs8hd_fill_1
XFILLER_40_102 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_ipin_5.LATCH_4_.latch/Q mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__127__B _128_/B vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_135 vgnd vpwr scs8hd_decap_8
XANTENNA__143__A _143_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_113 vgnd vpwr scs8hd_decap_8
XFILLER_13_135 vgnd vpwr scs8hd_decap_8
XFILLER_26_65 vgnd vpwr scs8hd_decap_4
XFILLER_42_75 vpwr vgnd scs8hd_fill_2
XFILLER_3_36 vpwr vgnd scs8hd_fill_2
XANTENNA__138__A _137_/X vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_2.LATCH_1_.latch data_in mem_left_ipin_2.LATCH_1_.latch/Q _085_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_127 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_3.LATCH_2_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_20 vpwr vgnd scs8hd_fill_2
XFILLER_37_97 vgnd vpwr scs8hd_decap_3
XFILLER_5_142 vgnd vpwr scs8hd_decap_4
Xmem_left_ipin_4.LATCH_4_.latch data_in mem_left_ipin_4.LATCH_4_.latch/Q _114_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__140__B _144_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_138 vpwr vgnd scs8hd_fill_2
XFILLER_4_90 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_1.LATCH_1_.latch/Q mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_55 vgnd vpwr scs8hd_decap_4
XFILLER_23_77 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_48_52 vpwr vgnd scs8hd_fill_2
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_35 vgnd vpwr scs8hd_fill_1
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
XANTENNA__119__C _094_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__135__B _135_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__151__A _070_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_44 vpwr vgnd scs8hd_fill_2
XFILLER_55_130 vpwr vgnd scs8hd_fill_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_4
XFILLER_50_75 vgnd vpwr scs8hd_decap_4
X_112_ _139_/A _116_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_59_73 vgnd vpwr scs8hd_decap_3
XFILLER_59_40 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[7] mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__146__A _145_/X vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XFILLER_52_133 vgnd vpwr scs8hd_decap_12
XFILLER_37_130 vgnd vpwr scs8hd_decap_4
XFILLER_37_141 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_67 vgnd vpwr scs8hd_decap_4
XFILLER_43_100 vpwr vgnd scs8hd_fill_2
XFILLER_29_65 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_5.LATCH_2_.latch/Q mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_45_53 vpwr vgnd scs8hd_fill_2
XFILLER_61_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_1.LATCH_3_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_125 vgnd vpwr scs8hd_decap_12
XFILLER_15_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_22 vgnd vpwr scs8hd_decap_4
XFILLER_31_88 vgnd vpwr scs8hd_decap_6
Xmux_left_ipin_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_144 vpwr vgnd scs8hd_fill_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _144_/B vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_3.LATCH_0_.latch/Q mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_114 vgnd vpwr scs8hd_decap_3
XFILLER_7_90 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_5.LATCH_0_.latch data_in mem_left_ipin_5.LATCH_0_.latch/Q _128_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_42_32 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_1.INVTX1_5_.scs8hd_inv_1 chany_top_in[5] mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_0.LATCH_4_.latch data_in mem_right_ipin_0.LATCH_4_.latch/Q _150_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _144_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_ipin_0.LATCH_3_.latch/Q mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmem_left_ipin_7.LATCH_3_.latch data_in mem_left_ipin_7.LATCH_3_.latch/Q _141_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_139 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_53_31 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_7.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[6] mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__149__A _139_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_7.LATCH_1_.latch/Q mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
XFILLER_48_97 vgnd vpwr scs8hd_fill_1
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_63 vgnd vpwr scs8hd_decap_12
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__151__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_ipin_4.LATCH_4_.latch/Q mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_34_88 vpwr vgnd scs8hd_fill_2
XFILLER_50_32 vgnd vpwr scs8hd_decap_4
X_111_ _110_/X _116_/B vgnd vpwr scs8hd_buf_1
XFILLER_38_109 vgnd vpwr scs8hd_decap_8
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_145 vgnd vpwr scs8hd_fill_1
XFILLER_1_92 vpwr vgnd scs8hd_fill_2
XANTENNA__072__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_46 vgnd vpwr scs8hd_decap_4
XFILLER_45_65 vgnd vpwr scs8hd_decap_3
XFILLER_43_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_55 vgnd vpwr scs8hd_fill_1
XFILLER_45_98 vgnd vpwr scs8hd_decap_3
XFILLER_45_87 vpwr vgnd scs8hd_fill_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__157__A _158_/A vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_1.LATCH_0_.latch data_in _160_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_137 vgnd vpwr scs8hd_decap_8
XFILLER_25_134 vgnd vpwr scs8hd_decap_12
XANTENNA__067__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_56_97 vgnd vpwr scs8hd_fill_1
XFILLER_56_86 vgnd vpwr scs8hd_decap_6
XFILLER_56_42 vpwr vgnd scs8hd_fill_2
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_1_.latch/Q mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_126 vgnd vpwr scs8hd_decap_12
XFILLER_26_23 vgnd vpwr scs8hd_decap_8
XFILLER_26_89 vgnd vpwr scs8hd_decap_3
XFILLER_42_88 vpwr vgnd scs8hd_fill_2
XFILLER_3_27 vgnd vpwr scs8hd_decap_6
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_6.LATCH_3_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__154__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _087_/X vgnd vpwr scs8hd_diode_2
XANTENNA__080__A _067_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_33 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_77 vpwr vgnd scs8hd_fill_2
XANTENNA__149__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _091_/X vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_4.LATCH_2_.latch/Q mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_35 vgnd vpwr scs8hd_fill_1
XANTENNA__075__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_32 vgnd vpwr scs8hd_decap_4
XFILLER_48_65 vpwr vgnd scs8hd_fill_2
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
Xmem_left_ipin_0.LATCH_4_.latch data_in mem_left_ipin_0.LATCH_4_.latch/Q _166_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_left_ipin_5.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_55_121 vgnd vpwr scs8hd_fill_1
X_110_ _137_/A address[4] address[3] _109_/Y _110_/X vgnd vpwr scs8hd_or4_4
XFILLER_34_45 vgnd vpwr scs8hd_decap_12
XFILLER_34_67 vpwr vgnd scs8hd_fill_2
XFILLER_59_97 vpwr vgnd scs8hd_fill_2
XFILLER_59_53 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_2.LATCH_0_.latch/Q mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__072__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_4.LATCH_4_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_34 vgnd vpwr scs8hd_decap_4
XFILLER_43_135 vgnd vpwr scs8hd_decap_8
XFILLER_28_121 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XFILLER_19_143 vgnd vpwr scs8hd_decap_3
XANTENNA__157__B _158_/B vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_25_113 vpwr vgnd scs8hd_fill_2
XFILLER_15_36 vgnd vpwr scs8hd_decap_3
XFILLER_15_58 vgnd vpwr scs8hd_decap_3
XANTENNA__083__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_56_65 vgnd vpwr scs8hd_decap_3
XFILLER_56_32 vgnd vpwr scs8hd_decap_6
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_102 vgnd vpwr scs8hd_decap_8
XFILLER_16_113 vgnd vpwr scs8hd_decap_8
XFILLER_16_124 vgnd vpwr scs8hd_decap_12
XFILLER_31_105 vpwr vgnd scs8hd_fill_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_6.LATCH_1_.latch/Q mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__168__A _081_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_138 vgnd vpwr scs8hd_decap_8
XFILLER_13_105 vpwr vgnd scs8hd_fill_2
XANTENNA__078__A _077_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__170__B _164_/X vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_ipin_3.LATCH_4_.latch/Q mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XFILLER_12_59 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _188_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__080__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_37_56 vpwr vgnd scs8hd_fill_2
XFILLER_53_99 vpwr vgnd scs8hd_fill_2
XFILLER_53_66 vgnd vpwr scs8hd_decap_3
XFILLER_53_55 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_2.LATCH_5_.latch_SLEEPB _179_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_112 vpwr vgnd scs8hd_fill_2
XFILLER_5_101 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_1.LATCH_0_.latch data_in mem_left_ipin_1.LATCH_0_.latch/Q _178_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__165__B _164_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__075__B _074_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_3.LATCH_3_.latch data_in mem_left_ipin_3.LATCH_3_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_38 vpwr vgnd scs8hd_fill_2
XFILLER_9_27 vgnd vpwr scs8hd_decap_8
X_186_ _186_/HI _186_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_49_141 vgnd vpwr scs8hd_decap_4
XFILLER_49_130 vpwr vgnd scs8hd_fill_2
XANTENNA__176__A _081_/X vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _188_/HI mem_left_ipin_7.LATCH_5_.latch/Q
+ mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_69 vgnd vpwr scs8hd_decap_3
XFILLER_50_23 vgnd vpwr scs8hd_decap_8
XANTENNA__086__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_34_57 vgnd vpwr scs8hd_fill_1
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
XFILLER_46_133 vgnd vpwr scs8hd_decap_12
XFILLER_46_122 vpwr vgnd scs8hd_fill_2
XFILLER_61_114 vpwr vgnd scs8hd_fill_2
XFILLER_61_103 vpwr vgnd scs8hd_fill_2
X_169_ _084_/X _164_/X _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_20_59 vpwr vgnd scs8hd_fill_2
XFILLER_43_114 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[3] mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_100 vpwr vgnd scs8hd_fill_2
XFILLER_19_111 vpwr vgnd scs8hd_fill_2
XANTENNA__157__C _068_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_125 vpwr vgnd scs8hd_fill_2
XANTENNA__173__B _172_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_106 vpwr vgnd scs8hd_fill_2
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__083__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_31_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_decap_3
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_136 vgnd vpwr scs8hd_decap_8
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__B _164_/X vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_3.LATCH_2_.latch/Q mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XANTENNA__094__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_26_36 vgnd vpwr scs8hd_fill_1
XFILLER_26_69 vgnd vpwr scs8hd_fill_1
XFILLER_42_79 vgnd vpwr scs8hd_decap_6
XFILLER_8_121 vgnd vpwr scs8hd_decap_12
XANTENNA__179__A _079_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_38 vgnd vpwr scs8hd_decap_6
Xmux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_1.LATCH_0_.latch/Q mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__080__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__089__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_53_78 vgnd vpwr scs8hd_decap_3
XFILLER_53_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_6.LATCH_2_.latch data_in mem_left_ipin_6.LATCH_2_.latch/Q _134_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XANTENNA__075__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_2_138 vgnd vpwr scs8hd_decap_8
XFILLER_64_77 vgnd vpwr scs8hd_decap_12
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_92 vgnd vpwr scs8hd_fill_1
X_185_ _185_/HI _185_/LO vgnd vpwr scs8hd_conb_1
XFILLER_64_145 vgnd vpwr scs8hd_fill_1
XANTENNA__176__B _172_/X vgnd vpwr scs8hd_diode_2
XANTENNA__192__A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XFILLER_55_134 vgnd vpwr scs8hd_decap_12
XFILLER_18_48 vgnd vpwr scs8hd_decap_4
XANTENNA__086__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_8_ vgnd vpwr scs8hd_inv_1
Xmux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_5.LATCH_1_.latch/Q mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_ipin_7.LATCH_5_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_46_145 vgnd vpwr scs8hd_fill_1
X_168_ _081_/X _164_/X _168_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
X_099_ _098_/X _100_/B vgnd vpwr scs8hd_buf_1
XFILLER_52_104 vpwr vgnd scs8hd_fill_2
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
XFILLER_1_73 vpwr vgnd scs8hd_fill_2
XFILLER_37_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB _178_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_145 vgnd vpwr scs8hd_fill_1
XFILLER_29_58 vgnd vpwr scs8hd_decap_3
XFILLER_29_69 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_5_ vgnd vpwr scs8hd_inv_1
XFILLER_45_57 vpwr vgnd scs8hd_fill_2
XFILLER_45_35 vgnd vpwr scs8hd_decap_4
XFILLER_43_104 vpwr vgnd scs8hd_fill_2
XANTENNA__097__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_61_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_ipin_2.LATCH_4_.latch/Q mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XFILLER_34_104 vpwr vgnd scs8hd_fill_2
XFILLER_15_27 vgnd vpwr scs8hd_decap_4
XFILLER_25_104 vpwr vgnd scs8hd_fill_2
XFILLER_25_126 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_4
XFILLER_31_26 vgnd vpwr scs8hd_fill_1
XANTENNA__083__C _068_/Y vgnd vpwr scs8hd_diode_2
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_92 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_1.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[1] mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_26_15 vgnd vpwr scs8hd_decap_4
XFILLER_26_48 vpwr vgnd scs8hd_fill_2
XFILLER_42_58 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_133 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _187_/HI mem_left_ipin_6.LATCH_5_.latch/Q
+ mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__179__B _091_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__195__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XFILLER_4_84 vgnd vpwr scs8hd_decap_4
XFILLER_4_73 vpwr vgnd scs8hd_fill_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_8
XFILLER_23_38 vpwr vgnd scs8hd_fill_2
XFILLER_2_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_121 vpwr vgnd scs8hd_fill_2
XFILLER_64_89 vgnd vpwr scs8hd_decap_4
XFILLER_64_56 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_71 vpwr vgnd scs8hd_fill_2
X_184_ _184_/HI _184_/LO vgnd vpwr scs8hd_conb_1
XFILLER_49_121 vgnd vpwr scs8hd_fill_1
XFILLER_55_113 vpwr vgnd scs8hd_fill_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XANTENNA__086__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_50_58 vpwr vgnd scs8hd_fill_2
XFILLER_50_36 vgnd vpwr scs8hd_fill_1
XFILLER_59_78 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_2.LATCH_2_.latch/Q mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_61_127 vpwr vgnd scs8hd_fill_2
X_167_ _070_/X _164_/X _167_/Y vgnd vpwr scs8hd_nor2_4
X_098_ address[1] _089_/Y address[0] _098_/X vgnd vpwr scs8hd_or3_4
XFILLER_37_102 vgnd vpwr scs8hd_decap_3
XFILLER_1_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_15 vgnd vpwr scs8hd_decap_3
XANTENNA__097__B _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_61_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_83 vgnd vpwr scs8hd_decap_8
XFILLER_19_135 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_0_.latch/Q mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__198__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_40_119 vgnd vpwr scs8hd_decap_4
XFILLER_56_46 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_decap_3
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_71 vgnd vpwr scs8hd_decap_3
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_30_130 vgnd vpwr scs8hd_decap_12
XFILLER_7_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_6.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_37 vpwr vgnd scs8hd_fill_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_145 vgnd vpwr scs8hd_fill_1
XFILLER_32_81 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_4.LATCH_1_.latch/Q mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_37 vpwr vgnd scs8hd_fill_2
XFILLER_53_47 vpwr vgnd scs8hd_fill_2
XFILLER_5_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_48_69 vgnd vpwr scs8hd_decap_6
XFILLER_48_36 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_ipin_1.LATCH_4_.latch/Q mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
XFILLER_64_125 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_2.LATCH_2_.latch data_in mem_left_ipin_2.LATCH_2_.latch/Q _082_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_50_48 vpwr vgnd scs8hd_fill_2
XFILLER_50_15 vgnd vpwr scs8hd_decap_4
XFILLER_59_57 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_6.INVTX1_3_.scs8hd_inv_1 chany_top_in[5] mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_4.LATCH_1_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_166_ _140_/A _164_/X _166_/Y vgnd vpwr scs8hd_nor2_4
X_097_ _139_/A _096_/X _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_70 vpwr vgnd scs8hd_fill_2
XFILLER_40_81 vpwr vgnd scs8hd_fill_2
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_37_114 vgnd vpwr scs8hd_decap_3
XFILLER_29_27 vpwr vgnd scs8hd_fill_2
XFILLER_29_38 vgnd vpwr scs8hd_fill_1
Xmem_left_ipin_4.LATCH_5_.latch data_in mem_left_ipin_4.LATCH_5_.latch/Q _112_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_45_15 vgnd vpwr scs8hd_decap_12
XFILLER_28_125 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _186_/HI mem_left_ipin_5.LATCH_5_.latch/Q
+ mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_70 vpwr vgnd scs8hd_fill_2
X_149_ _139_/A _149_/B _149_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_117 vpwr vgnd scs8hd_fill_2
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_decap_3
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_109 vgnd vpwr scs8hd_decap_12
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_22_109 vgnd vpwr scs8hd_decap_3
XFILLER_30_142 vgnd vpwr scs8hd_decap_4
XFILLER_13_109 vpwr vgnd scs8hd_fill_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_131 vgnd vpwr scs8hd_decap_12
XFILLER_32_60 vpwr vgnd scs8hd_fill_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_2.LATCH_2_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_1.LATCH_2_.latch/Q mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_16 vpwr vgnd scs8hd_fill_2
XFILLER_53_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_116 vgnd vpwr scs8hd_decap_6
XFILLER_43_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_48_48 vpwr vgnd scs8hd_fill_2
XFILLER_48_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_119 vgnd vpwr scs8hd_decap_12
XFILLER_58_145 vgnd vpwr scs8hd_fill_1
X_182_ _182_/HI _182_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_95 vgnd vpwr scs8hd_fill_1
XFILLER_49_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_5.LATCH_1_.latch data_in mem_left_ipin_5.LATCH_1_.latch/Q _127_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_64_137 vgnd vpwr scs8hd_decap_8
XANTENNA__100__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_0.LATCH_5_.latch data_in mem_right_ipin_0.LATCH_5_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_55_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_36 vpwr vgnd scs8hd_fill_2
XFILLER_61_118 vpwr vgnd scs8hd_fill_2
XFILLER_61_107 vgnd vpwr scs8hd_decap_4
XFILLER_46_126 vgnd vpwr scs8hd_decap_4
Xmem_left_ipin_7.LATCH_4_.latch data_in mem_left_ipin_7.LATCH_4_.latch/Q _140_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_165_ _091_/X _164_/X _165_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_72 vpwr vgnd scs8hd_fill_2
XFILLER_24_83 vgnd vpwr scs8hd_decap_4
X_096_ _095_/X _096_/X vgnd vpwr scs8hd_buf_1
XFILLER_1_21 vgnd vpwr scs8hd_fill_1
XFILLER_37_126 vpwr vgnd scs8hd_fill_2
XFILLER_37_137 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_104 vgnd vpwr scs8hd_decap_8
XFILLER_45_27 vgnd vpwr scs8hd_decap_6
XFILLER_43_118 vgnd vpwr scs8hd_fill_1
XFILLER_28_137 vgnd vpwr scs8hd_decap_8
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_83 vpwr vgnd scs8hd_fill_2
XFILLER_19_104 vpwr vgnd scs8hd_fill_2
XFILLER_19_115 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_81 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_3.LATCH_1_.latch/Q mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
X_148_ _147_/X _149_/B vgnd vpwr scs8hd_buf_1
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
X_079_ _141_/A _079_/B _079_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_ipin_4.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_29 vpwr vgnd scs8hd_fill_2
XFILLER_56_15 vgnd vpwr scs8hd_decap_12
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_75 vgnd vpwr scs8hd_decap_4
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_42 vgnd vpwr scs8hd_decap_6
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_ipin_0.LATCH_4_.latch/Q mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_12_143 vgnd vpwr scs8hd_decap_3
XFILLER_16_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__103__A _134_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_7.LATCH_2_.latch/Q mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_27 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_1.LATCH_1_.latch data_in _159_/A _155_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_54 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_48_27 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _185_/HI mem_left_ipin_4.LATCH_5_.latch/Q
+ mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
X_181_ _181_/HI _181_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_131 vpwr vgnd scs8hd_fill_2
XFILLER_1_142 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_14_ vgnd vpwr scs8hd_inv_1
XANTENNA__100__B _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_71 vgnd vpwr scs8hd_decap_4
XFILLER_38_93 vgnd vpwr scs8hd_decap_4
XFILLER_55_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_7.LATCH_2_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_55_105 vpwr vgnd scs8hd_fill_2
XFILLER_59_15 vgnd vpwr scs8hd_decap_12
XANTENNA__201__A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_46_105 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_095_ _137_/A _074_/Y _094_/Y _072_/X _095_/X vgnd vpwr scs8hd_or4_4
X_164_ _163_/X _164_/X vgnd vpwr scs8hd_buf_1
XFILLER_52_108 vgnd vpwr scs8hd_decap_4
XFILLER_49_92 vpwr vgnd scs8hd_fill_2
XFILLER_1_77 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _110_/X vgnd vpwr scs8hd_diode_2
XFILLER_60_130 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_39 vgnd vpwr scs8hd_fill_1
XFILLER_43_108 vgnd vpwr scs8hd_decap_3
XFILLER_61_27 vgnd vpwr scs8hd_decap_12
XFILLER_19_40 vpwr vgnd scs8hd_fill_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_4
XFILLER_34_108 vgnd vpwr scs8hd_decap_4
XFILLER_35_83 vgnd vpwr scs8hd_decap_3
XANTENNA__106__A _087_/X vgnd vpwr scs8hd_diode_2
X_078_ _077_/X _079_/B vgnd vpwr scs8hd_buf_1
X_147_ _137_/A address[4] address[3] _158_/B _147_/X vgnd vpwr scs8hd_or4_4
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_2_.latch/Q mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_130 vpwr vgnd scs8hd_fill_2
XFILLER_33_141 vgnd vpwr scs8hd_decap_4
XFILLER_31_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_38 vgnd vpwr scs8hd_fill_1
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XPHY_103 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_0.LATCH_5_.latch data_in mem_left_ipin_0.LATCH_5_.latch/Q _165_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_52 vgnd vpwr scs8hd_decap_3
XFILLER_46_93 vgnd vpwr scs8hd_decap_3
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_26_19 vgnd vpwr scs8hd_fill_1
XFILLER_21_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_5.LATCH_3_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_2.INVTX1_3_.scs8hd_inv_1 chany_top_in[2] mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_52 vpwr vgnd scs8hd_fill_2
XFILLER_8_104 vpwr vgnd scs8hd_fill_2
XFILLER_12_100 vpwr vgnd scs8hd_fill_2
XANTENNA__103__B _096_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__204__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_62 vpwr vgnd scs8hd_fill_2
XANTENNA__114__A _140_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_125 vgnd vpwr scs8hd_decap_8
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_31 vgnd vpwr scs8hd_fill_1
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XFILLER_13_75 vpwr vgnd scs8hd_fill_2
X_180_ _079_/B _100_/B _180_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_121 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_2.LATCH_1_.latch/Q mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_106 vgnd vpwr scs8hd_decap_12
XFILLER_54_71 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
XFILLER_55_117 vpwr vgnd scs8hd_fill_2
XFILLER_59_27 vgnd vpwr scs8hd_decap_6
XFILLER_24_41 vgnd vpwr scs8hd_decap_3
X_094_ address[3] _094_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_left_ipin_3.LATCH_4_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
X_163_ _137_/A address[4] address[3] _072_/X _163_/X vgnd vpwr scs8hd_or4_4
XFILLER_49_71 vgnd vpwr scs8hd_decap_4
XFILLER_60_142 vgnd vpwr scs8hd_decap_4
Xmem_left_ipin_1.LATCH_1_.latch data_in mem_left_ipin_1.LATCH_1_.latch/Q _177_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_39 vgnd vpwr scs8hd_decap_12
XFILLER_10_32 vgnd vpwr scs8hd_decap_8
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_42_131 vgnd vpwr scs8hd_decap_12
XFILLER_35_62 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_6.LATCH_2_.latch/Q mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _162_/A vgnd vpwr
+ scs8hd_diode_2
X_146_ _145_/X _158_/B vgnd vpwr scs8hd_buf_1
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
X_077_ _072_/X _158_/A _077_/X vgnd vpwr scs8hd_or2_4
Xmem_left_ipin_3.LATCH_4_.latch data_in mem_left_ipin_3.LATCH_4_.latch/Q _100_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_25_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_0_.latch/Q mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__207__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XPHY_126 vgnd vpwr scs8hd_decap_3
XPHY_115 vgnd vpwr scs8hd_decap_3
XPHY_104 vgnd vpwr scs8hd_decap_3
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_83 vpwr vgnd scs8hd_fill_2
XFILLER_46_61 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__117__A _143_/A vgnd vpwr scs8hd_diode_2
X_129_ _158_/A _109_/Y _129_/X vgnd vpwr scs8hd_or2_4
Xmux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _184_/HI mem_left_ipin_3.LATCH_5_.latch/Q
+ mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_123 vpwr vgnd scs8hd_fill_2
XFILLER_21_145 vgnd vpwr scs8hd_fill_1
XFILLER_32_85 vgnd vpwr scs8hd_decap_4
XFILLER_57_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_1.LATCH_5_.latch_SLEEPB _173_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_62 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_0.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__114__B _116_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__130__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_67 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_58_137 vgnd vpwr scs8hd_decap_8
XFILLER_58_104 vpwr vgnd scs8hd_fill_2
XFILLER_49_137 vpwr vgnd scs8hd_fill_2
XFILLER_49_126 vpwr vgnd scs8hd_fill_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_64_118 vgnd vpwr scs8hd_decap_6
XFILLER_38_84 vpwr vgnd scs8hd_fill_2
XANTENNA__109__B _145_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _141_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_6.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_50_19 vgnd vpwr scs8hd_fill_1
Xmem_left_ipin_4.LATCH_0_.latch data_in mem_left_ipin_4.LATCH_0_.latch/Q _118_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_162_ _162_/A _162_/Y vgnd vpwr scs8hd_inv_8
X_093_ _075_/A _137_/A vgnd vpwr scs8hd_buf_1
XFILLER_40_74 vgnd vpwr scs8hd_decap_4
XFILLER_40_85 vpwr vgnd scs8hd_fill_2
XFILLER_49_50 vgnd vpwr scs8hd_decap_4
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_7.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_51_143 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_6.LATCH_3_.latch data_in mem_left_ipin_6.LATCH_3_.latch/Q _133_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_66 vgnd vpwr scs8hd_decap_8
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_42_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_30 vpwr vgnd scs8hd_fill_2
X_145_ address[5] _145_/B _145_/X vgnd vpwr scs8hd_or2_4
XFILLER_51_73 vpwr vgnd scs8hd_fill_2
XFILLER_51_51 vgnd vpwr scs8hd_decap_4
XFILLER_51_40 vpwr vgnd scs8hd_fill_2
X_076_ _075_/X _158_/A vgnd vpwr scs8hd_buf_1
XFILLER_33_121 vgnd vpwr scs8hd_fill_1
XFILLER_56_29 vpwr vgnd scs8hd_fill_2
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
XFILLER_24_121 vgnd vpwr scs8hd_decap_8
XFILLER_24_132 vgnd vpwr scs8hd_decap_12
XPHY_127 vgnd vpwr scs8hd_decap_3
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_76 vgnd vpwr scs8hd_decap_3
XFILLER_46_40 vpwr vgnd scs8hd_fill_2
XFILLER_46_73 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_110 vpwr vgnd scs8hd_fill_2
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XANTENNA__133__A _141_/A vgnd vpwr scs8hd_diode_2
X_128_ _144_/A _128_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__117__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_1.LATCH_1_.latch/Q mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_6
XFILLER_16_65 vpwr vgnd scs8hd_fill_2
XFILLER_32_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_57_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_31 vpwr vgnd scs8hd_fill_2
XFILLER_27_42 vpwr vgnd scs8hd_fill_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XFILLER_43_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XFILLER_4_46 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_0.LATCH_0_.latch data_in mem_right_ipin_0.LATCH_0_.latch/Q _154_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_5.LATCH_2_.latch/Q mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_88 vgnd vpwr scs8hd_decap_4
XFILLER_38_63 vpwr vgnd scs8hd_fill_2
XFILLER_54_84 vpwr vgnd scs8hd_fill_2
XANTENNA__125__B _128_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _141_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_6.LATCH_5_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
X_161_ _161_/A _161_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_6
XFILLER_24_76 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _183_/HI mem_left_ipin_2.LATCH_5_.latch/Q
+ mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_092_ _091_/X _139_/A vgnd vpwr scs8hd_buf_1
XFILLER_40_42 vpwr vgnd scs8hd_fill_2
XFILLER_40_53 vpwr vgnd scs8hd_fill_2
XFILLER_1_25 vpwr vgnd scs8hd_fill_2
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XFILLER_37_119 vgnd vpwr scs8hd_decap_3
XANTENNA__136__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_53_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_4.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_87 vpwr vgnd scs8hd_fill_2
XFILLER_19_119 vgnd vpwr scs8hd_decap_3
X_144_ _144_/A _144_/B _144_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_51_85 vpwr vgnd scs8hd_fill_2
X_075_ _075_/A _074_/Y address[3] _075_/X vgnd vpwr scs8hd_or3_4
XFILLER_18_130 vgnd vpwr scs8hd_decap_12
XFILLER_33_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XPHY_106 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_5.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_144 vpwr vgnd scs8hd_fill_2
XFILLER_21_22 vpwr vgnd scs8hd_fill_2
XFILLER_21_33 vpwr vgnd scs8hd_fill_2
XFILLER_21_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_84 vgnd vpwr scs8hd_decap_8
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA__133__B _135_/B vgnd vpwr scs8hd_diode_2
X_127_ _143_/A _128_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_16_88 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vpwr vgnd scs8hd_fill_2
XFILLER_32_43 vpwr vgnd scs8hd_fill_2
XFILLER_32_98 vpwr vgnd scs8hd_fill_2
XANTENNA__144__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _128_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_98 vpwr vgnd scs8hd_fill_2
XFILLER_43_53 vgnd vpwr scs8hd_decap_4
XFILLER_43_42 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_34 vpwr vgnd scs8hd_fill_2
XFILLER_1_113 vpwr vgnd scs8hd_fill_2
XFILLER_38_42 vgnd vpwr scs8hd_decap_3
XFILLER_38_97 vgnd vpwr scs8hd_fill_1
XANTENNA__141__B _144_/B vgnd vpwr scs8hd_diode_2
XFILLER_55_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_109 vpwr vgnd scs8hd_fill_2
XFILLER_24_55 vgnd vpwr scs8hd_decap_6
X_091_ _091_/A _091_/X vgnd vpwr scs8hd_buf_1
X_160_ _160_/A _160_/Y vgnd vpwr scs8hd_inv_8
XFILLER_40_32 vgnd vpwr scs8hd_fill_1
XFILLER_49_96 vpwr vgnd scs8hd_fill_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_6
XANTENNA__136__B _135_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_1_.latch/Q mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__152__A _134_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _161_/A mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_46_3 vgnd vpwr scs8hd_decap_12
XFILLER_51_123 vgnd vpwr scs8hd_decap_12
X_143_ _143_/A _144_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_0.LATCH_0_.latch data_in mem_left_ipin_0.LATCH_0_.latch/Q _170_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_074_ address[4] _074_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_142 vgnd vpwr scs8hd_decap_4
XFILLER_33_145 vgnd vpwr scs8hd_fill_1
XANTENNA__147__A _137_/A vgnd vpwr scs8hd_diode_2
XPHY_129 vgnd vpwr scs8hd_decap_3
XPHY_118 vgnd vpwr scs8hd_decap_3
XPHY_107 vgnd vpwr scs8hd_decap_3
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_2.LATCH_3_.latch data_in mem_left_ipin_2.LATCH_3_.latch/Q _079_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_62_74 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_ipin_5.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_145 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_2.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_126_ _134_/A _128_/B _126_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_115 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_4.LATCH_2_.latch/Q mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_108 vgnd vpwr scs8hd_decap_4
XFILLER_32_77 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_3.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__144__B _144_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_109_ address[5] _145_/B _109_/Y vgnd vpwr scs8hd_nand2_4
XANTENNA__160__A _160_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_90 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _182_/HI mem_left_ipin_1.LATCH_5_.latch/Q
+ mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__070__A _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_22 vgnd vpwr scs8hd_decap_6
XFILLER_27_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XANTENNA__139__B _144_/B vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_54_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _161_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_63_143 vgnd vpwr scs8hd_decap_3
XFILLER_63_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_ipin_3.LATCH_1_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_80 vpwr vgnd scs8hd_fill_2
XFILLER_24_89 vgnd vpwr scs8hd_decap_3
X_090_ address[1] _089_/Y _068_/Y _091_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_45_132 vgnd vpwr scs8hd_decap_12
XFILLER_45_110 vgnd vpwr scs8hd_decap_3
XANTENNA__152__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XFILLER_51_135 vgnd vpwr scs8hd_decap_8
XFILLER_36_121 vpwr vgnd scs8hd_fill_2
XFILLER_27_132 vgnd vpwr scs8hd_decap_12
XFILLER_35_22 vgnd vpwr scs8hd_decap_6
X_142_ _134_/A _144_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_35_66 vpwr vgnd scs8hd_fill_2
XFILLER_35_88 vpwr vgnd scs8hd_fill_2
X_073_ enable _075_/A vgnd vpwr scs8hd_inv_8
XFILLER_33_113 vpwr vgnd scs8hd_fill_2
XANTENNA__147__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__163__A _137_/A vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_5.LATCH_2_.latch data_in mem_left_ipin_5.LATCH_2_.latch/Q _126_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_119 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_decap_3
XANTENNA__073__A enable vgnd vpwr scs8hd_diode_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_87 vgnd vpwr scs8hd_decap_3
XFILLER_46_65 vgnd vpwr scs8hd_decap_8
XFILLER_46_32 vgnd vpwr scs8hd_fill_1
XFILLER_62_97 vgnd vpwr scs8hd_decap_12
XFILLER_62_64 vgnd vpwr scs8hd_fill_1
X_125_ _141_/A _128_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_90 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_7.LATCH_5_.latch data_in mem_left_ipin_7.LATCH_5_.latch/Q _139_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__158__A _158_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_127 vgnd vpwr scs8hd_decap_12
XANTENNA__068__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_1.LATCH_2_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_23 vgnd vpwr scs8hd_decap_8
XFILLER_32_89 vgnd vpwr scs8hd_fill_1
XFILLER_57_75 vpwr vgnd scs8hd_fill_2
XFILLER_57_53 vpwr vgnd scs8hd_fill_2
XFILLER_57_42 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
X_108_ address[6] _145_/B vgnd vpwr scs8hd_inv_8
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_0.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _159_/A mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__155__B _158_/B vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__171__A _072_/X vgnd vpwr scs8hd_diode_2
XFILLER_58_108 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__081__A _080_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_88 vgnd vpwr scs8hd_decap_4
XFILLER_54_54 vpwr vgnd scs8hd_fill_2
XFILLER_54_43 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _140_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_7.INVTX1_1_.scs8hd_inv_1 chany_top_in[2] mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__076__A _075_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_23 vpwr vgnd scs8hd_fill_2
XFILLER_40_89 vgnd vpwr scs8hd_decap_3
XFILLER_49_54 vgnd vpwr scs8hd_fill_1
XFILLER_60_125 vgnd vpwr scs8hd_fill_1
XFILLER_60_103 vpwr vgnd scs8hd_fill_2
XFILLER_45_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_3.LATCH_2_.latch/Q mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_51_114 vpwr vgnd scs8hd_fill_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
XFILLER_19_68 vpwr vgnd scs8hd_fill_2
XFILLER_27_144 vpwr vgnd scs8hd_fill_2
XFILLER_35_34 vpwr vgnd scs8hd_fill_2
X_141_ _141_/A _144_/B _141_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_51_77 vpwr vgnd scs8hd_fill_2
XFILLER_51_55 vgnd vpwr scs8hd_fill_1
X_072_ address[5] address[6] _072_/X vgnd vpwr scs8hd_or2_4
XANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__147__C address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__163__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_51_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _181_/HI mem_left_ipin_0.LATCH_5_.latch/Q
+ mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_71 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
X_124_ _140_/A _128_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__158__B _158_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_139 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_16_69 vpwr vgnd scs8hd_fill_2
XANTENNA__084__A _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_57_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_143 vgnd vpwr scs8hd_decap_3
X_107_ _144_/A _096_/X _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XANTENNA__169__A _084_/X vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XFILLER_27_35 vpwr vgnd scs8hd_fill_2
XFILLER_27_46 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _141_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_79 vgnd vpwr scs8hd_decap_6
XFILLER_4_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__155__C _068_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_1_ vgnd vpwr scs8hd_inv_1
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_6.LATCH_2_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_49_109 vgnd vpwr scs8hd_decap_12
XFILLER_1_127 vpwr vgnd scs8hd_fill_2
XFILLER_1_138 vpwr vgnd scs8hd_fill_2
XFILLER_38_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_67 vpwr vgnd scs8hd_fill_2
XFILLER_54_88 vgnd vpwr scs8hd_decap_4
XFILLER_63_123 vgnd vpwr scs8hd_decap_12
XANTENNA__166__B _164_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_46 vpwr vgnd scs8hd_fill_2
XFILLER_40_57 vpwr vgnd scs8hd_fill_2
XFILLER_49_77 vpwr vgnd scs8hd_fill_2
XFILLER_49_33 vpwr vgnd scs8hd_fill_2
XFILLER_49_22 vgnd vpwr scs8hd_decap_8
XFILLER_1_29 vpwr vgnd scs8hd_fill_2
XFILLER_14_80 vpwr vgnd scs8hd_fill_2
XANTENNA__177__A _084_/X vgnd vpwr scs8hd_diode_2
XFILLER_51_104 vpwr vgnd scs8hd_fill_2
XFILLER_10_49 vgnd vpwr scs8hd_decap_6
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_19_36 vpwr vgnd scs8hd_fill_2
XFILLER_42_115 vpwr vgnd scs8hd_fill_2
XFILLER_42_104 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A _086_/X vgnd vpwr scs8hd_diode_2
XFILLER_51_89 vpwr vgnd scs8hd_fill_2
XFILLER_51_34 vgnd vpwr scs8hd_decap_4
X_140_ _140_/A _144_/B _140_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_071_ _070_/X _141_/A vgnd vpwr scs8hd_buf_1
Xmux_left_ipin_5.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_decap_3
XFILLER_33_126 vpwr vgnd scs8hd_fill_2
XFILLER_33_137 vpwr vgnd scs8hd_fill_2
XANTENNA__147__D _158_/B vgnd vpwr scs8hd_diode_2
XANTENNA__163__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_44_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_4
XFILLER_21_26 vgnd vpwr scs8hd_decap_4
XFILLER_21_37 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_ipin_0.LATCH_3_.latch/Q mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_46_23 vpwr vgnd scs8hd_fill_2
XFILLER_62_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_30_107 vgnd vpwr scs8hd_decap_8
XFILLER_30_118 vgnd vpwr scs8hd_decap_12
X_123_ _139_/A _128_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_39 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_ipin_4.LATCH_3_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_6.INVTX1_5_.scs8hd_inv_1 chany_top_in[6] mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__158__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__174__B _172_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_107 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_1.LATCH_2_.latch data_in mem_left_ipin_1.LATCH_2_.latch/Q _176_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_107 vgnd vpwr scs8hd_decap_12
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_48 vpwr vgnd scs8hd_fill_2
XFILLER_32_47 vgnd vpwr scs8hd_decap_4
XFILLER_22_91 vgnd vpwr scs8hd_fill_1
X_106_ _087_/X _144_/A vgnd vpwr scs8hd_buf_1
XANTENNA__169__B _164_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_3.LATCH_5_.latch data_in mem_left_ipin_3.LATCH_5_.latch/Q _097_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _162_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__079__B _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_43_35 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A _137_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_2.LATCH_2_.latch/Q mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_114 vgnd vpwr scs8hd_decap_8
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_38 vpwr vgnd scs8hd_fill_2
XFILLER_57_132 vpwr vgnd scs8hd_fill_2
XFILLER_1_117 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_35 vgnd vpwr scs8hd_decap_4
XFILLER_63_135 vgnd vpwr scs8hd_decap_8
XFILLER_63_113 vgnd vpwr scs8hd_decap_8
XFILLER_48_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_2.LATCH_4_.latch_SLEEPB _180_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_132 vgnd vpwr scs8hd_decap_12
XFILLER_39_110 vpwr vgnd scs8hd_fill_2
XFILLER_54_113 vgnd vpwr scs8hd_decap_12
XFILLER_54_102 vpwr vgnd scs8hd_fill_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__177__B _172_/X vgnd vpwr scs8hd_diode_2
XANTENNA__193__A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_1_.latch/Q mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_102 vgnd vpwr scs8hd_decap_4
XFILLER_27_113 vpwr vgnd scs8hd_fill_2
XFILLER_35_47 vpwr vgnd scs8hd_fill_2
X_070_ _069_/X _070_/X vgnd vpwr scs8hd_buf_1
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_102 vgnd vpwr scs8hd_decap_8
XPHY_91 vgnd vpwr scs8hd_decap_3
XPHY_80 vgnd vpwr scs8hd_decap_3
X_199_ chany_top_in[1] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__163__D _072_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_57 vpwr vgnd scs8hd_fill_2
XANTENNA__098__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_62_56 vgnd vpwr scs8hd_decap_8
XFILLER_15_127 vgnd vpwr scs8hd_decap_12
X_122_ _122_/A _128_/B vgnd vpwr scs8hd_buf_1
Xmem_left_ipin_4.LATCH_1_.latch data_in mem_left_ipin_4.LATCH_1_.latch/Q _117_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_119 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_3.INVTX1_1_.scs8hd_inv_1 chany_top_in[2] mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_12_119 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_38 vgnd vpwr scs8hd_fill_1
XFILLER_32_15 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XFILLER_57_23 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_6.LATCH_4_.latch data_in mem_left_ipin_6.LATCH_4_.latch/Q _132_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XFILLER_22_70 vpwr vgnd scs8hd_fill_2
X_105_ _143_/A _096_/X _105_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_83 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_4.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_15 vgnd vpwr scs8hd_decap_4
XANTENNA__095__B _074_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_126 vgnd vpwr scs8hd_decap_8
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ _162_/A mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__196__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_144 vpwr vgnd scs8hd_fill_2
XFILLER_38_58 vgnd vpwr scs8hd_decap_3
XFILLER_54_79 vpwr vgnd scs8hd_fill_2
XFILLER_54_35 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_3
XFILLER_39_144 vpwr vgnd scs8hd_fill_2
XFILLER_5_84 vpwr vgnd scs8hd_fill_2
XFILLER_54_125 vgnd vpwr scs8hd_decap_12
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_24_38 vgnd vpwr scs8hd_fill_1
XFILLER_40_15 vgnd vpwr scs8hd_decap_4
XFILLER_49_57 vpwr vgnd scs8hd_fill_2
XFILLER_60_117 vgnd vpwr scs8hd_decap_8
XFILLER_30_70 vgnd vpwr scs8hd_decap_3
XFILLER_36_125 vgnd vpwr scs8hd_decap_4
XFILLER_35_15 vgnd vpwr scs8hd_decap_4
XFILLER_51_58 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_0.LATCH_1_.latch data_in mem_right_ipin_0.LATCH_1_.latch/Q _153_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_33_117 vpwr vgnd scs8hd_fill_2
XPHY_92 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
X_198_ chany_top_in[2] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_2_63 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_7.LATCH_4_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_1.LATCH_2_.latch/Q mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_left_ipin_7.LATCH_0_.latch data_in mem_left_ipin_7.LATCH_0_.latch/Q _144_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_36 vpwr vgnd scs8hd_fill_2
XFILLER_15_106 vpwr vgnd scs8hd_fill_2
XFILLER_15_139 vgnd vpwr scs8hd_decap_6
XANTENNA__098__B _089_/Y vgnd vpwr scs8hd_diode_2
X_121_ _109_/Y _121_/B _122_/A vgnd vpwr scs8hd_or2_4
XANTENNA_mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__199__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_79 vpwr vgnd scs8hd_fill_2
XFILLER_57_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_135 vgnd vpwr scs8hd_decap_8
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
X_104_ _084_/X _143_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mem_left_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_43_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__095__C _094_/Y vgnd vpwr scs8hd_diode_2
XFILLER_43_59 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_138 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_81 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_fill_1
XFILLER_54_58 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_5.LATCH_5_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_2.INVTX1_5_.scs8hd_inv_1 chany_top_in[6] mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_63_104 vgnd vpwr scs8hd_fill_1
XFILLER_44_91 vgnd vpwr scs8hd_fill_1
XFILLER_54_137 vgnd vpwr scs8hd_decap_8
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_60_107 vgnd vpwr scs8hd_decap_6
XFILLER_45_126 vgnd vpwr scs8hd_decap_4
XFILLER_45_115 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_104 vpwr vgnd scs8hd_fill_2
XFILLER_39_91 vpwr vgnd scs8hd_fill_2
XFILLER_51_118 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_51_15 vgnd vpwr scs8hd_decap_12
XPHY_82 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_93 vgnd vpwr scs8hd_decap_3
XFILLER_41_81 vgnd vpwr scs8hd_decap_3
X_197_ chany_top_in[3] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_46_15 vgnd vpwr scs8hd_decap_8
XANTENNA__098__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_15_118 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _160_/A mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_120_ _119_/X _121_/B vgnd vpwr scs8hd_buf_1
XFILLER_11_40 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vpwr vgnd scs8hd_fill_2
XFILLER_11_73 vpwr vgnd scs8hd_fill_2
XFILLER_52_80 vpwr vgnd scs8hd_fill_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_36 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_12_ vgnd vpwr scs8hd_inv_1
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_11_143 vgnd vpwr scs8hd_decap_3
XFILLER_22_83 vpwr vgnd scs8hd_fill_2
X_103_ _134_/A _096_/X _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_47_91 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_0.LATCH_1_.latch data_in mem_left_ipin_0.LATCH_1_.latch/Q _169_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_43_38 vpwr vgnd scs8hd_fill_2
XFILLER_43_27 vgnd vpwr scs8hd_decap_8
XANTENNA__095__D _072_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_106 vgnd vpwr scs8hd_decap_4
XFILLER_17_83 vpwr vgnd scs8hd_fill_2
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_60 vgnd vpwr scs8hd_fill_1
Xmem_left_ipin_2.LATCH_4_.latch data_in mem_left_ipin_2.LATCH_4_.latch/Q _180_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_27 vpwr vgnd scs8hd_fill_2
XFILLER_57_113 vpwr vgnd scs8hd_fill_2
XFILLER_54_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_48_135 vgnd vpwr scs8hd_decap_8
XFILLER_48_124 vgnd vpwr scs8hd_decap_8
XFILLER_28_82 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _191_/HI _161_/Y mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_2_.latch/Q mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_97 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_37 vpwr vgnd scs8hd_fill_2
XFILLER_49_15 vgnd vpwr scs8hd_decap_4
XFILLER_14_40 vgnd vpwr scs8hd_decap_4
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__101__A _141_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_138 vgnd vpwr scs8hd_decap_8
XFILLER_51_108 vgnd vpwr scs8hd_decap_4
XFILLER_19_29 vpwr vgnd scs8hd_fill_2
XFILLER_42_119 vgnd vpwr scs8hd_decap_12
XFILLER_42_108 vgnd vpwr scs8hd_decap_4
XFILLER_51_27 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_7.LATCH_0_.latch/Q mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_94 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_25_83 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
X_196_ chany_top_in[4] chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_3
XFILLER_24_108 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_6.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[5] mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_4.LATCH_0_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _161_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_27 vgnd vpwr scs8hd_decap_4
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_141 vgnd vpwr scs8hd_decap_4
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
X_179_ _079_/B _091_/X _179_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_15 vgnd vpwr scs8hd_decap_8
Xmem_left_ipin_3.LATCH_0_.latch data_in mem_left_ipin_3.LATCH_0_.latch/Q _107_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_40 vpwr vgnd scs8hd_fill_2
X_102_ _081_/X _134_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_5.LATCH_3_.latch data_in mem_left_ipin_5.LATCH_3_.latch/Q _125_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_62 vgnd vpwr scs8hd_decap_4
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _084_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_39 vgnd vpwr scs8hd_fill_1
XFILLER_57_136 vgnd vpwr scs8hd_decap_8
XFILLER_54_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_2.LATCH_1_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_93 vgnd vpwr scs8hd_decap_3
XFILLER_39_114 vpwr vgnd scs8hd_fill_2
XFILLER_54_106 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_0_.latch/Q mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_63 vpwr vgnd scs8hd_fill_2
XFILLER_30_84 vgnd vpwr scs8hd_decap_8
XANTENNA__101__B _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_55_92 vpwr vgnd scs8hd_fill_2
XFILLER_27_117 vgnd vpwr scs8hd_decap_3
XANTENNA__202__A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XPHY_95 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
X_195_ chany_top_in[5] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_2_44 vpwr vgnd scs8hd_fill_2
XANTENNA__112__A _139_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XFILLER_32_120 vgnd vpwr scs8hd_decap_12
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
XFILLER_23_131 vgnd vpwr scs8hd_decap_3
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_11_86 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__107__A _144_/A vgnd vpwr scs8hd_diode_2
X_178_ _087_/X _172_/X _178_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_19 vgnd vpwr scs8hd_fill_1
XFILLER_20_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_4.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
X_101_ _141_/A _096_/X _101_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _190_/HI _159_/Y mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_70 vgnd vpwr scs8hd_decap_3
XFILLER_8_87 vgnd vpwr scs8hd_fill_1
XFILLER_8_43 vpwr vgnd scs8hd_fill_2
XFILLER_8_32 vgnd vpwr scs8hd_decap_8
XFILLER_27_19 vgnd vpwr scs8hd_fill_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_4
XANTENNA__120__A _119_/X vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_6.LATCH_0_.latch/Q mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__205__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_133 vgnd vpwr scs8hd_decap_12
XFILLER_28_62 vpwr vgnd scs8hd_fill_2
XFILLER_60_93 vgnd vpwr scs8hd_fill_1
XFILLER_60_71 vpwr vgnd scs8hd_fill_2
XANTENNA__115__A _141_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_19 vgnd vpwr scs8hd_fill_1
XFILLER_30_52 vpwr vgnd scs8hd_fill_2
XFILLER_30_96 vgnd vpwr scs8hd_decap_4
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XFILLER_35_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_140 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_ipin_7.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_26_140 vgnd vpwr scs8hd_decap_6
XPHY_96 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_143 vgnd vpwr scs8hd_decap_3
XFILLER_41_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_25_41 vpwr vgnd scs8hd_fill_2
XFILLER_25_52 vgnd vpwr scs8hd_decap_4
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
XFILLER_41_73 vpwr vgnd scs8hd_fill_2
XFILLER_41_62 vpwr vgnd scs8hd_fill_2
X_194_ chany_top_in[6] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_2_67 vpwr vgnd scs8hd_fill_2
XANTENNA__112__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_132 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_84 vpwr vgnd scs8hd_fill_2
X_177_ _084_/X _172_/X _177_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__107__B _096_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XFILLER_20_113 vgnd vpwr scs8hd_decap_12
XANTENNA__208__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_135 vgnd vpwr scs8hd_decap_8
XFILLER_22_53 vgnd vpwr scs8hd_decap_4
X_100_ _096_/X _100_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_97 vgnd vpwr scs8hd_decap_3
XFILLER_47_72 vpwr vgnd scs8hd_fill_2
XANTENNA__118__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_66 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_42 vpwr vgnd scs8hd_fill_2
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_52 vpwr vgnd scs8hd_fill_2
XFILLER_33_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_5.LATCH_2_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_142 vgnd vpwr scs8hd_decap_4
XFILLER_3_131 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_2.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[2] mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_123 vgnd vpwr scs8hd_fill_1
XFILLER_0_145 vgnd vpwr scs8hd_fill_1
XFILLER_28_52 vgnd vpwr scs8hd_decap_4
XFILLER_44_84 vgnd vpwr scs8hd_decap_4
Xmem_left_ipin_1.LATCH_3_.latch data_in mem_left_ipin_1.LATCH_3_.latch/Q _175_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_60_50 vgnd vpwr scs8hd_fill_1
XFILLER_5_67 vpwr vgnd scs8hd_fill_2
XANTENNA__115__B _116_/B vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _139_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_119 vgnd vpwr scs8hd_fill_1
XFILLER_14_32 vgnd vpwr scs8hd_decap_4
XFILLER_14_76 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_108 vpwr vgnd scs8hd_fill_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_3
XFILLER_39_95 vpwr vgnd scs8hd_fill_2
XFILLER_55_83 vgnd vpwr scs8hd_decap_6
XANTENNA__126__A _134_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_50_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_ipin_0.LATCH_4_.latch/Q mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_18_119 vgnd vpwr scs8hd_decap_8
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_decap_3
X_193_ chany_top_in[7] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XPHY_75 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_130 vpwr vgnd scs8hd_fill_2
XFILLER_32_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_3.LATCH_3_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_100 vpwr vgnd scs8hd_fill_2
XFILLER_11_33 vgnd vpwr scs8hd_fill_1
XFILLER_52_51 vgnd vpwr scs8hd_decap_4
XFILLER_52_84 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_5.LATCH_0_.latch/Q mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_176_ _081_/X _172_/X _176_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__123__B _128_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_125 vgnd vpwr scs8hd_decap_12
XFILLER_11_103 vpwr vgnd scs8hd_fill_2
XFILLER_7_118 vgnd vpwr scs8hd_decap_4
XFILLER_22_32 vgnd vpwr scs8hd_decap_8
XFILLER_22_87 vgnd vpwr scs8hd_decap_4
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_95 vpwr vgnd scs8hd_fill_2
XFILLER_47_62 vgnd vpwr scs8hd_fill_1
XANTENNA__118__B _116_/B vgnd vpwr scs8hd_diode_2
XANTENNA__134__A _134_/A vgnd vpwr scs8hd_diode_2
X_159_ _159_/A _159_/Y vgnd vpwr scs8hd_inv_8
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_0.INVTX1_3_.scs8hd_inv_1 chany_top_in[7] mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_87 vgnd vpwr scs8hd_decap_4
XFILLER_33_31 vpwr vgnd scs8hd_fill_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__129__A _158_/A vgnd vpwr scs8hd_diode_2
XFILLER_57_117 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_4.LATCH_2_.latch data_in mem_left_ipin_4.LATCH_2_.latch/Q _116_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_1.LATCH_4_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
XFILLER_63_109 vpwr vgnd scs8hd_fill_2
XFILLER_44_74 vgnd vpwr scs8hd_fill_1
XFILLER_60_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__131__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB _155_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_6.LATCH_5_.latch data_in mem_left_ipin_6.LATCH_5_.latch/Q _131_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_left_ipin_0.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_2_.latch/Q mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_88 vgnd vpwr scs8hd_decap_4
XFILLER_30_32 vgnd vpwr scs8hd_decap_4
XFILLER_30_65 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_74 vpwr vgnd scs8hd_fill_2
XFILLER_55_62 vgnd vpwr scs8hd_decap_4
XFILLER_55_40 vpwr vgnd scs8hd_fill_2
XANTENNA__126__B _128_/B vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _134_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_98 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_decap_3
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XFILLER_41_101 vpwr vgnd scs8hd_fill_2
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_decap_3
XFILLER_41_97 vpwr vgnd scs8hd_fill_2
XFILLER_41_53 vpwr vgnd scs8hd_fill_2
X_192_ chany_top_in[8] chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_25_98 vgnd vpwr scs8hd_decap_4
XANTENNA__137__A _137_/A vgnd vpwr scs8hd_diode_2
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
XFILLER_23_145 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_7.INVTX1_3_.scs8hd_inv_1 chany_top_in[6] mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_53 vgnd vpwr scs8hd_decap_3
XFILLER_52_63 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vgnd vpwr scs8hd_fill_1
X_175_ _070_/X _172_/X _175_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_20_137 vgnd vpwr scs8hd_decap_8
XFILLER_3_90 vpwr vgnd scs8hd_fill_2
XFILLER_7_108 vgnd vpwr scs8hd_decap_4
XFILLER_22_66 vpwr vgnd scs8hd_fill_2
XFILLER_63_51 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ _162_/Y mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_63_84 vgnd vpwr scs8hd_decap_12
XFILLER_63_62 vgnd vpwr scs8hd_fill_1
XANTENNA__134__B _135_/B vgnd vpwr scs8hd_diode_2
X_158_ _158_/A _158_/B address[0] _158_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_6_141 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_0.LATCH_2_.latch data_in mem_right_ipin_0.LATCH_2_.latch/Q _152_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_089_ address[2] _089_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__150__A _140_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _160_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_ipin_7.LATCH_1_.latch data_in mem_left_ipin_7.LATCH_1_.latch/Q _143_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_58_84 vgnd vpwr scs8hd_decap_6
XFILLER_58_62 vpwr vgnd scs8hd_fill_2
XANTENNA__129__B _109_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__145__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XFILLER_48_107 vgnd vpwr scs8hd_decap_8
XFILLER_28_32 vgnd vpwr scs8hd_decap_6
XFILLER_44_53 vgnd vpwr scs8hd_decap_4
XFILLER_5_47 vgnd vpwr scs8hd_fill_1
XFILLER_39_118 vpwr vgnd scs8hd_fill_2
XFILLER_53_143 vgnd vpwr scs8hd_decap_3
XFILLER_53_121 vgnd vpwr scs8hd_fill_1
XFILLER_38_140 vgnd vpwr scs8hd_decap_6
Xmux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_4.LATCH_0_.latch/Q mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_53 vpwr vgnd scs8hd_fill_2
XANTENNA__142__B _144_/B vgnd vpwr scs8hd_diode_2
XFILLER_50_124 vgnd vpwr scs8hd_decap_12
XFILLER_50_113 vgnd vpwr scs8hd_decap_8
XFILLER_50_102 vpwr vgnd scs8hd_fill_2
XFILLER_35_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_6.LATCH_4_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XPHY_99 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_decap_3
XFILLER_41_135 vgnd vpwr scs8hd_decap_8
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_25_22 vgnd vpwr scs8hd_decap_8
XFILLER_25_66 vpwr vgnd scs8hd_fill_2
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_2_48 vpwr vgnd scs8hd_fill_2
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_17_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__137__B _074_/Y vgnd vpwr scs8hd_diode_2
XFILLER_56_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _143_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_113 vpwr vgnd scs8hd_fill_2
XFILLER_11_57 vgnd vpwr scs8hd_decap_4
XFILLER_36_32 vgnd vpwr scs8hd_decap_4
XFILLER_36_65 vpwr vgnd scs8hd_fill_2
X_174_ _100_/B _172_/X _174_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__148__A _147_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _181_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_45 vpwr vgnd scs8hd_fill_2
XFILLER_47_53 vpwr vgnd scs8hd_fill_2
XFILLER_63_96 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_5.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_157_ _158_/A _158_/B _068_/Y _157_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_8_47 vpwr vgnd scs8hd_fill_2
XANTENNA__150__B _149_/B vgnd vpwr scs8hd_diode_2
X_088_ _079_/B _087_/X _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_44 vpwr vgnd scs8hd_fill_2
XFILLER_33_77 vpwr vgnd scs8hd_fill_2
XFILLER_3_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_4.LATCH_5_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
X_209_ chany_bottom_in[0] chany_top_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA__145__B _145_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_115 vpwr vgnd scs8hd_fill_2
XANTENNA__071__A _070_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_66 vgnd vpwr scs8hd_decap_3
XFILLER_44_98 vpwr vgnd scs8hd_fill_2
XFILLER_44_32 vgnd vpwr scs8hd_decap_6
XFILLER_60_75 vgnd vpwr scs8hd_decap_6
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_47_130 vpwr vgnd scs8hd_fill_2
XANTENNA__156__A _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_0.LATCH_2_.latch data_in mem_left_ipin_0.LATCH_2_.latch/Q _168_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_39_32 vpwr vgnd scs8hd_fill_2
XFILLER_55_53 vpwr vgnd scs8hd_fill_2
XFILLER_44_122 vgnd vpwr scs8hd_decap_12
XFILLER_44_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_50_136 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_6_80 vpwr vgnd scs8hd_fill_2
XPHY_12 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_2.LATCH_5_.latch data_in mem_left_ipin_2.LATCH_5_.latch/Q _179_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_111 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _160_/Y mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_ipin_7.LATCH_3_.latch/Q mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_89 vgnd vpwr scs8hd_decap_3
XFILLER_41_114 vgnd vpwr scs8hd_decap_8
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XFILLER_41_77 vpwr vgnd scs8hd_fill_2
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XANTENNA__137__C _094_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__153__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_49_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_4_ vgnd vpwr scs8hd_inv_1
Xmux_right_ipin_2.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_36 vpwr vgnd scs8hd_fill_2
XFILLER_11_69 vpwr vgnd scs8hd_fill_2
XFILLER_36_88 vgnd vpwr scs8hd_decap_4
XFILLER_52_32 vgnd vpwr scs8hd_decap_6
X_173_ _091_/X _172_/X _173_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vgnd vpwr scs8hd_decap_4
XANTENNA__164__A _163_/X vgnd vpwr scs8hd_diode_2
XANTENNA__074__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_47_76 vpwr vgnd scs8hd_fill_2
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
X_087_ _086_/X _087_/X vgnd vpwr scs8hd_buf_1
X_156_ _121_/B _158_/B address[0] _156_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__159__A _159_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_3.LATCH_0_.latch/Q mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__069__A _067_/Y vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_46 vpwr vgnd scs8hd_fill_2
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_17_68 vpwr vgnd scs8hd_fill_2
XFILLER_33_23 vgnd vpwr scs8hd_fill_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_56 vpwr vgnd scs8hd_fill_2
X_208_ chany_bottom_in[1] chany_top_out[1] vgnd vpwr scs8hd_buf_2
X_139_ _139_/A _144_/B _139_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_3.INVTX1_3_.scs8hd_inv_1 chany_top_in[3] mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_23 vgnd vpwr scs8hd_decap_8
XFILLER_28_78 vpwr vgnd scs8hd_fill_2
XFILLER_44_88 vgnd vpwr scs8hd_fill_1
XFILLER_44_66 vgnd vpwr scs8hd_decap_6
XFILLER_60_54 vgnd vpwr scs8hd_decap_6
XFILLER_60_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_3.LATCH_1_.latch data_in mem_left_ipin_3.LATCH_1_.latch/Q _105_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _171_/X vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _158_/B vgnd vpwr scs8hd_diode_2
XFILLER_53_123 vgnd vpwr scs8hd_decap_12
XFILLER_14_36 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_7.LATCH_1_.latch/Q mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__082__A _079_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_39_99 vpwr vgnd scs8hd_fill_2
XFILLER_44_134 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_5.LATCH_4_.latch data_in mem_left_ipin_5.LATCH_4_.latch/Q _124_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__167__A _070_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_70 vgnd vpwr scs8hd_fill_1
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_25_35 vgnd vpwr scs8hd_decap_4
XFILLER_26_101 vgnd vpwr scs8hd_fill_1
XANTENNA__077__A _072_/X vgnd vpwr scs8hd_diode_2
XPHY_79 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_3.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_79 vpwr vgnd scs8hd_fill_2
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XANTENNA__137__D _109_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_134 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_126 vgnd vpwr scs8hd_decap_3
XFILLER_23_137 vpwr vgnd scs8hd_fill_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_104 vgnd vpwr scs8hd_decap_8
XFILLER_14_115 vgnd vpwr scs8hd_decap_12
XFILLER_36_23 vpwr vgnd scs8hd_fill_2
XFILLER_52_88 vgnd vpwr scs8hd_decap_4
XFILLER_52_55 vgnd vpwr scs8hd_fill_1
X_172_ _171_/X _172_/X vgnd vpwr scs8hd_buf_1
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XANTENNA__180__A _079_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _182_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_71 vpwr vgnd scs8hd_fill_2
XFILLER_11_107 vgnd vpwr scs8hd_decap_12
XANTENNA__090__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_0.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_91 vgnd vpwr scs8hd_fill_1
X_086_ address[1] address[2] address[0] _086_/X vgnd vpwr scs8hd_or3_4
X_155_ _121_/B _158_/B _068_/Y _155_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _070_/X vgnd vpwr scs8hd_diode_2
XANTENNA__069__B address[2] vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__A _079_/B vgnd vpwr scs8hd_diode_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_58_43 vpwr vgnd scs8hd_fill_2
XFILLER_58_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
X_207_ chany_bottom_in[2] chany_top_out[2] vgnd vpwr scs8hd_buf_2
X_138_ _137_/X _144_/B vgnd vpwr scs8hd_buf_1
X_069_ _067_/Y address[2] _068_/Y _069_/X vgnd vpwr scs8hd_or3_4
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_ipin_6.LATCH_3_.latch/Q mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_1_.latch/Q mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_81 vgnd vpwr scs8hd_decap_4
Xmem_left_ipin_6.LATCH_0_.latch data_in mem_left_ipin_6.LATCH_0_.latch/Q _136_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_143 vgnd vpwr scs8hd_decap_3
XFILLER_5_39 vgnd vpwr scs8hd_decap_8
XFILLER_47_110 vpwr vgnd scs8hd_fill_2
XANTENNA__156__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_53_135 vgnd vpwr scs8hd_decap_8
XFILLER_53_113 vpwr vgnd scs8hd_fill_2
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__082__B _081_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_36 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_1.INVTX1_3_.scs8hd_inv_1 chany_top_in[1] mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_143 vgnd vpwr scs8hd_decap_3
XFILLER_39_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__167__B _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_25_58 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _158_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_57 vpwr vgnd scs8hd_fill_2
XANTENNA__093__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_102 vpwr vgnd scs8hd_fill_2
XFILLER_17_113 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_2.LATCH_0_.latch/Q mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_ipin_7.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _159_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__178__A _087_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_27 vgnd vpwr scs8hd_decap_6
XANTENNA__088__A _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_127 vgnd vpwr scs8hd_decap_12
XFILLER_52_67 vpwr vgnd scs8hd_fill_2
X_171_ _072_/X _121_/B _171_/X vgnd vpwr scs8hd_or2_4
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XANTENNA__180__B _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_94 vpwr vgnd scs8hd_fill_2
XFILLER_11_119 vgnd vpwr scs8hd_decap_3
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA__090__B _089_/Y vgnd vpwr scs8hd_diode_2
XFILLER_47_34 vpwr vgnd scs8hd_fill_2
XFILLER_63_66 vpwr vgnd scs8hd_fill_2
XFILLER_6_145 vgnd vpwr scs8hd_fill_1
XFILLER_12_81 vpwr vgnd scs8hd_fill_2
X_085_ _079_/B _084_/X _085_/Y vgnd vpwr scs8hd_nor2_4
X_154_ _144_/A _149_/B _154_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__175__B _172_/X vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_6.LATCH_1_.latch/Q mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_ipin_2.LATCH_0_.latch data_in _162_/A _158_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XANTENNA__069__C _068_/Y vgnd vpwr scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__B _084_/X vgnd vpwr scs8hd_diode_2
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_59_130 vpwr vgnd scs8hd_fill_2
XFILLER_58_66 vpwr vgnd scs8hd_fill_2
X_206_ chany_bottom_in[3] chany_top_out[3] vgnd vpwr scs8hd_buf_2
X_137_ _137_/A _074_/Y _094_/Y _109_/Y _137_/X vgnd vpwr scs8hd_or4_4
X_068_ address[0] _068_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_73 vpwr vgnd scs8hd_fill_2
XFILLER_56_111 vgnd vpwr scs8hd_fill_1
XFILLER_0_107 vpwr vgnd scs8hd_fill_2
XFILLER_0_129 vpwr vgnd scs8hd_fill_2
XFILLER_28_58 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _095_/X vgnd vpwr scs8hd_diode_2
XFILLER_62_114 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_103 vgnd vpwr scs8hd_fill_1
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_30_48 vpwr vgnd scs8hd_fill_2
XFILLER_39_57 vpwr vgnd scs8hd_fill_2
XFILLER_55_89 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_6.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_50_106 vgnd vpwr scs8hd_decap_4
XFILLER_35_103 vpwr vgnd scs8hd_fill_2
XFILLER_35_114 vpwr vgnd scs8hd_fill_2
XFILLER_35_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_4
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_41_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__194__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__178__B _172_/X vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_1.LATCH_4_.latch data_in mem_left_ipin_1.LATCH_4_.latch/Q _174_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__088__B _087_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_58 vpwr vgnd scs8hd_fill_2
XFILLER_36_69 vpwr vgnd scs8hd_fill_2
X_170_ _087_/X _164_/X _170_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_139 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_ipin_5.LATCH_3_.latch/Q mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_9_143 vgnd vpwr scs8hd_decap_3
XFILLER_9_110 vpwr vgnd scs8hd_fill_2
XFILLER_47_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_5.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XFILLER_22_49 vpwr vgnd scs8hd_fill_2
XANTENNA__090__C _068_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__099__A _098_/X vgnd vpwr scs8hd_diode_2
XFILLER_47_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
X_153_ _143_/A _149_/B _153_/Y vgnd vpwr scs8hd_nor2_4
X_084_ _083_/X _084_/X vgnd vpwr scs8hd_buf_1
Xmux_left_ipin_6.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_4.LATCH_2_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_15 vgnd vpwr scs8hd_decap_8
XFILLER_33_48 vpwr vgnd scs8hd_fill_2
XFILLER_3_138 vpwr vgnd scs8hd_fill_2
XFILLER_3_127 vpwr vgnd scs8hd_fill_2
XFILLER_3_116 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_205_ chany_bottom_in[4] chany_top_out[4] vgnd vpwr scs8hd_buf_2
X_136_ _144_/A _135_/B _136_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_81 vpwr vgnd scs8hd_fill_2
X_067_ address[1] _067_/Y vgnd vpwr scs8hd_inv_8
XFILLER_0_41 vpwr vgnd scs8hd_fill_2
XFILLER_0_63 vgnd vpwr scs8hd_fill_1
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_119 vgnd vpwr scs8hd_decap_4
XFILLER_28_15 vgnd vpwr scs8hd_decap_4
XFILLER_60_46 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_1.LATCH_0_.latch/Q mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_62_126 vgnd vpwr scs8hd_decap_12
XFILLER_47_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
X_119_ _137_/A address[4] _094_/Y _119_/X vgnd vpwr scs8hd_or3_4
XANTENNA__197__A chany_top_in[3] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _189_/HI mem_right_ipin_0.LATCH_5_.latch/Q
+ mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_55_57 vpwr vgnd scs8hd_fill_2
XFILLER_44_115 vgnd vpwr scs8hd_decap_4
XFILLER_29_101 vgnd vpwr scs8hd_decap_3
XFILLER_29_112 vpwr vgnd scs8hd_fill_2
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XFILLER_55_79 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_2.LATCH_0_.latch data_in mem_left_ipin_2.LATCH_0_.latch/Q _088_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vgnd vpwr scs8hd_decap_8
XFILLER_6_62 vpwr vgnd scs8hd_fill_2
XFILLER_26_115 vgnd vpwr scs8hd_decap_4
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_2.LATCH_3_.latch_SLEEPB _079_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_4.LATCH_3_.latch data_in mem_left_ipin_4.LATCH_3_.latch/Q _115_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_126 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_5.LATCH_1_.latch/Q mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XFILLER_15_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_15 vgnd vpwr scs8hd_fill_1
XFILLER_52_47 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_9_ vgnd vpwr scs8hd_inv_1
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
X_152_ _134_/A _149_/B _152_/Y vgnd vpwr scs8hd_nor2_4
X_083_ address[1] address[2] _068_/Y _083_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_27 vpwr vgnd scs8hd_fill_2
XFILLER_59_121 vgnd vpwr scs8hd_fill_1
XFILLER_59_110 vgnd vpwr scs8hd_decap_3
XFILLER_58_79 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_3.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_204_ chany_bottom_in[5] chany_top_out[5] vgnd vpwr scs8hd_buf_2
X_135_ _143_/A _135_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_73 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_7.LATCH_0_.latch/Q mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_135 vgnd vpwr scs8hd_decap_8
XFILLER_56_124 vgnd vpwr scs8hd_decap_8
XFILLER_28_38 vgnd vpwr scs8hd_fill_1
XFILLER_44_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_4.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_62_138 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_118_ _144_/A _116_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_124 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_0.LATCH_3_.latch data_in mem_right_ipin_0.LATCH_3_.latch/Q _151_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_15 vpwr vgnd scs8hd_fill_2
XFILLER_55_36 vpwr vgnd scs8hd_fill_2
XFILLER_29_135 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_ipin_4.LATCH_3_.latch/Q mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _160_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_45_91 vgnd vpwr scs8hd_decap_4
Xmem_left_ipin_7.LATCH_2_.latch data_in mem_left_ipin_7.LATCH_2_.latch/Q _142_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_52 vgnd vpwr scs8hd_fill_1
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_71 vpwr vgnd scs8hd_fill_2
XFILLER_52_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_36_38 vpwr vgnd scs8hd_fill_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_26_93 vpwr vgnd scs8hd_fill_2
XFILLER_3_75 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_0_.latch/Q mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _184_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_47_15 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_ipin_7.LATCH_3_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
X_151_ _070_/X _149_/B _151_/Y vgnd vpwr scs8hd_nor2_4
X_082_ _079_/B _081_/X _082_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_81 vgnd vpwr scs8hd_decap_3
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_107 vgnd vpwr scs8hd_decap_3
XFILLER_58_47 vpwr vgnd scs8hd_fill_2
X_203_ chany_bottom_in[6] chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_134_ _134_/A _135_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_9_85 vgnd vpwr scs8hd_fill_1
XFILLER_56_114 vgnd vpwr scs8hd_fill_1
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_49 vpwr vgnd scs8hd_fill_2
XFILLER_44_27 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_4.LATCH_1_.latch/Q mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_114 vpwr vgnd scs8hd_fill_2
XFILLER_18_61 vgnd vpwr scs8hd_decap_8
XFILLER_34_71 vpwr vgnd scs8hd_fill_2
X_117_ _143_/A _116_/B _117_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_ipin_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_53_117 vgnd vpwr scs8hd_decap_4
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_29_82 vpwr vgnd scs8hd_fill_2
XFILLER_45_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_5.LATCH_4_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_2.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_61_91 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_26_128 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_106 vpwr vgnd scs8hd_fill_2
XFILLER_17_117 vpwr vgnd scs8hd_fill_2
XFILLER_32_109 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _081_/X vgnd vpwr scs8hd_diode_2
XFILLER_52_27 vgnd vpwr scs8hd_decap_4
XFILLER_9_135 vgnd vpwr scs8hd_decap_8
Xmem_left_ipin_0.LATCH_3_.latch data_in mem_left_ipin_0.LATCH_3_.latch/Q _167_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_72 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_6.LATCH_0_.latch/Q mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XFILLER_47_38 vpwr vgnd scs8hd_fill_2
XFILLER_63_59 vpwr vgnd scs8hd_fill_2
X_150_ _140_/A _149_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_145 vgnd vpwr scs8hd_fill_1
XFILLER_12_85 vgnd vpwr scs8hd_decap_6
XFILLER_12_96 vpwr vgnd scs8hd_fill_2
X_081_ _080_/X _081_/X vgnd vpwr scs8hd_buf_1
XFILLER_37_60 vgnd vpwr scs8hd_fill_1
XFILLER_37_71 vgnd vpwr scs8hd_decap_4
XFILLER_45_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_ipin_3.LATCH_3_.latch/Q mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_left_ipin_3.LATCH_5_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_15 vgnd vpwr scs8hd_decap_12
XANTENNA__200__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
X_202_ chany_bottom_in[7] chany_top_out[7] vgnd vpwr scs8hd_buf_2
X_133_ _141_/A _135_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_51 vpwr vgnd scs8hd_fill_2
XFILLER_23_73 vpwr vgnd scs8hd_fill_2
XANTENNA__110__A _137_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_9_42 vpwr vgnd scs8hd_fill_2
XFILLER_0_77 vpwr vgnd scs8hd_fill_2
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_18_40 vgnd vpwr scs8hd_fill_1
XFILLER_18_84 vgnd vpwr scs8hd_decap_6
XFILLER_50_82 vgnd vpwr scs8hd_decap_8
XFILLER_50_71 vpwr vgnd scs8hd_fill_2
XANTENNA__105__A _143_/A vgnd vpwr scs8hd_diode_2
X_116_ _134_/A _116_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_55_27 vgnd vpwr scs8hd_decap_6
Xmux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_ipin_7.LATCH_4_.latch/Q mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_ipin_0.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_63 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_107 vpwr vgnd scs8hd_fill_2
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_25_19 vgnd vpwr scs8hd_fill_1
XFILLER_15_41 vgnd vpwr scs8hd_decap_3
XFILLER_31_40 vpwr vgnd scs8hd_fill_2
XFILLER_56_70 vgnd vpwr scs8hd_decap_3
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_121 vgnd vpwr scs8hd_fill_1
XFILLER_31_143 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_ipin_3.LATCH_2_.latch data_in mem_left_ipin_3.LATCH_2_.latch/Q _103_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_18 vpwr vgnd scs8hd_fill_2
XANTENNA__203__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_3
XFILLER_9_114 vgnd vpwr scs8hd_decap_8
XFILLER_9_103 vpwr vgnd scs8hd_fill_2
XFILLER_13_121 vgnd vpwr scs8hd_fill_1
XFILLER_13_143 vgnd vpwr scs8hd_decap_3
XANTENNA__113__A _100_/B vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_3.LATCH_1_.latch/Q mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_left_ipin_5.LATCH_5_.latch data_in mem_left_ipin_5.LATCH_5_.latch/Q _123_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _185_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XFILLER_6_106 vgnd vpwr scs8hd_decap_8
X_080_ _067_/Y address[2] address[0] _080_/X vgnd vpwr scs8hd_or3_4
Xmux_left_ipin_6.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_12_64 vgnd vpwr scs8hd_fill_1
XANTENNA__108__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
X_201_ chany_bottom_in[8] chany_top_out[8] vgnd vpwr scs8hd_buf_2
Xmux_left_ipin_7.INVTX1_5_.scs8hd_inv_1 chany_top_in[7] mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_132_ _140_/A _135_/B _132_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_96 vpwr vgnd scs8hd_fill_2
XFILLER_2_131 vgnd vpwr scs8hd_decap_3
XFILLER_48_93 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_28_19 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_7.LATCH_2_.latch/Q mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_47_138 vgnd vpwr scs8hd_decap_8
XFILLER_18_74 vgnd vpwr scs8hd_fill_1
XFILLER_34_84 vpwr vgnd scs8hd_fill_2
XANTENNA__105__B _096_/X vgnd vpwr scs8hd_diode_2
X_115_ _141_/A _116_/B _115_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__121__A _109_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_116 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__206__A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_42 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_5.LATCH_0_.latch/Q mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_86 vgnd vpwr scs8hd_decap_6
XFILLER_29_51 vgnd vpwr scs8hd_decap_4
XFILLER_45_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_2.LATCH_0_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__116__A _134_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_66 vpwr vgnd scs8hd_fill_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_8
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_130 vpwr vgnd scs8hd_fill_2
XFILLER_15_53 vgnd vpwr scs8hd_decap_3
XFILLER_15_75 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_6.LATCH_1_.latch data_in mem_left_ipin_6.LATCH_1_.latch/Q _135_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_93 vpwr vgnd scs8hd_fill_2
XFILLER_56_82 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_ipin_2.LATCH_3_.latch/Q mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

