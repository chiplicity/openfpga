* NGSPICE file created from cby_2__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

.subckt cby_2__1_ ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11]
+ chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15]
+ chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0]
+ chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12] chany_bottom_out[13]
+ chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16] chany_bottom_out[17]
+ chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in[0] chany_top_in[10]
+ chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15]
+ chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10]
+ chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15]
+ chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6]
+ chany_top_out[7] chany_top_out[8] chany_top_out[9] gfpga_pad_EMBEDDED_IO_SOC_DIR
+ gfpga_pad_EMBEDDED_IO_SOC_IN gfpga_pad_EMBEDDED_IO_SOC_OUT left_grid_pin_16_ left_grid_pin_17_
+ left_grid_pin_18_ left_grid_pin_19_ left_grid_pin_20_ left_grid_pin_21_ left_grid_pin_22_
+ left_grid_pin_23_ left_grid_pin_24_ left_grid_pin_25_ left_grid_pin_26_ left_grid_pin_27_
+ left_grid_pin_28_ left_grid_pin_29_ left_grid_pin_30_ left_grid_pin_31_ left_width_0_height_0__pin_0_
+ left_width_0_height_0__pin_1_lower left_width_0_height_0__pin_1_upper prog_clk right_grid_pin_0_
+ VPWR VGND
XANTENNA_mux_right_ipin_1.mux_l3_in_0__A1 mux_right_ipin_1.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_ipin_0.mux_l2_in_1__A1 mux_left_ipin_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_3.mux_l2_in_0__S mux_right_ipin_3.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_8.mux_l4_in_0__A0 mux_right_ipin_8.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_11.mux_l2_in_0_ mux_right_ipin_11.mux_l1_in_1_/X mux_right_ipin_11.mux_l1_in_0_/X
+ mux_right_ipin_11.mux_l2_in_0_/S mux_right_ipin_11.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0__S mux_left_ipin_0.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_66_ chany_bottom_in[7] chany_top_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_15.mux_l1_in_0_/S mux_right_ipin_15.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_23_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_ipin_0.mux_l3_in_0__A1 mux_left_ipin_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_1_0_prog_clk_A clkbuf_2_0_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_prog_clk clkbuf_3_5_0_prog_clk/A clkbuf_3_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
X_49_ chany_top_in[4] chany_bottom_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_2.mux_l3_in_0__S mux_right_ipin_2.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_11.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_11.mux_l1_in_0_/S
+ mux_right_ipin_11.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_47_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_11.mux_l1_in_1__A1 chany_bottom_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_50_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_8.mux_l2_in_1__S mux_right_ipin_8.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_11.mux_l4_in_0_/S mux_right_ipin_12.mux_l1_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_8.mux_l2_in_2__A1 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_11.mux_l1_in_0__S mux_right_ipin_11.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_3.mux_l2_in_3__S mux_right_ipin_3.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_11.mux_l2_in_0__A1 mux_right_ipin_11.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_1.mux_l4_in_0__S mux_right_ipin_1.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_ipin_0.mux_l2_in_3__S mux_left_ipin_0.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_8.mux_l3_in_1__A1 mux_right_ipin_8.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_7.mux_l3_in_1__S mux_right_ipin_7.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_10.mux_l2_in_0__S mux_right_ipin_10.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_0.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_5.mux_l2_in_0__A0 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_8.mux_l4_in_0__A1 mux_right_ipin_8.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_8.mux_l4_in_0_/X left_grid_pin_24_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_65_ chany_bottom_in[8] chany_top_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_14.mux_l4_in_0_/S mux_right_ipin_15.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_2__A0 chany_bottom_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_48_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_48_ chany_top_in[5] chany_bottom_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_ipin_11.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_11.mux_l1_in_0_/S
+ mux_right_ipin_11.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_15.mux_l2_in_1__S mux_right_ipin_15.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_14.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_3.mux_l3_in_1__A0 mux_right_ipin_3.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_10.mux_l2_in_3__S mux_right_ipin_10.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_7.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_3.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_14.mux_l3_in_1__S mux_right_ipin_14.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_3.mux_l4_in_0__A0 mux_right_ipin_3.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_15.mux_l1_in_0__A0 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0__S mux_right_ipin_0.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_5.mux_l2_in_0__A1 mux_right_ipin_5.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_64_ chany_bottom_in[9] chany_top_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_ipin_3.mux_l2_in_3_ _31_/HI chany_top_in[14] mux_right_ipin_3.mux_l2_in_3_/S
+ mux_right_ipin_3.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_59_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_15.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.mux_l2_in_2__A1 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_47_ chany_top_in[6] chany_bottom_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_6.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_13.mux_l2_in_1__A0 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_0.mux_l1_in_1__A0 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.mux_l3_in_1__A1 mux_right_ipin_3.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_1_0_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_11.mux_l2_in_3__A0 _25_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_3.mux_l4_in_0_ mux_right_ipin_3.mux_l3_in_1_/X mux_right_ipin_3.mux_l3_in_0_/X
+ mux_right_ipin_3.mux_l4_in_0_/S mux_right_ipin_3.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_13.mux_l3_in_0__A0 mux_right_ipin_13.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_4.mux_l2_in_1__S mux_right_ipin_4.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_0.mux_l2_in_0__A0 mux_right_ipin_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_8.mux_l2_in_3_ _19_/HI chany_top_in[19] mux_right_ipin_8.mux_l2_in_2_/S
+ mux_right_ipin_8.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_3.mux_l4_in_0__A1 mux_right_ipin_3.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1_0_prog_clk clkbuf_2_0_0_prog_clk/A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_3.mux_l3_in_1_ mux_right_ipin_3.mux_l2_in_3_/X mux_right_ipin_3.mux_l2_in_2_/X
+ mux_right_ipin_3.mux_l3_in_1_/S mux_right_ipin_3.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_15.mux_l1_in_0__A1 chany_bottom_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D mux_left_ipin_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.mux_l3_in_1__S mux_right_ipin_3.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_9.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_ipin_0.mux_l3_in_1__S mux_left_ipin_0.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_63_ chany_bottom_in[10] chany_top_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_ipin_3.mux_l2_in_2_ chany_bottom_in[14] chany_top_in[8] mux_right_ipin_3.mux_l2_in_3_/S
+ mux_right_ipin_3.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_9.mux_l2_in_2__S mux_right_ipin_9.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_8.mux_l4_in_0_ mux_right_ipin_8.mux_l3_in_1_/X mux_right_ipin_8.mux_l3_in_0_/X
+ mux_right_ipin_8.mux_l4_in_0_/S mux_right_ipin_8.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_9.mux_l1_in_0__A0 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l1_in_1__S mux_right_ipin_12.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_46_ chany_top_in[7] chany_bottom_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_13.mux_l2_in_1__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_7.mux_l1_in_2__A0 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_8.mux_l3_in_1_ mux_right_ipin_8.mux_l2_in_3_/X mux_right_ipin_8.mux_l2_in_2_/X
+ mux_right_ipin_8.mux_l3_in_1_/S mux_right_ipin_8.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_0.mux_l1_in_1__A1 chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_1.mux_l4_in_0_/X left_grid_pin_17_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29_ _29_/HI _29_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_ipin_11.mux_l2_in_3__A1 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_11.mux_l2_in_1__S mux_right_ipin_11.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_ipin_13.mux_l3_in_0__A1 mux_right_ipin_13.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_10.mux_l1_in_0__A0 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_7.mux_l2_in_1__A0 chany_bottom_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_0.mux_l2_in_0__A1 mux_right_ipin_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_8.mux_l2_in_2_ chany_bottom_in[19] chany_top_in[13] mux_right_ipin_8.mux_l2_in_2_/S
+ mux_right_ipin_8.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_3.mux_l3_in_0_ mux_right_ipin_3.mux_l2_in_1_/X mux_right_ipin_3.mux_l2_in_0_/X
+ mux_right_ipin_3.mux_l3_in_1_/S mux_right_ipin_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_5.mux_l2_in_3__A0 _33_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_10.mux_l3_in_1__S mux_right_ipin_10.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_7.mux_l3_in_0__A0 mux_right_ipin_7.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_62_ chany_bottom_in[11] chany_top_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_ipin_3.mux_l2_in_1_ chany_bottom_in[8] mux_right_ipin_3.mux_l1_in_2_/X
+ mux_right_ipin_3.mux_l2_in_3_/S mux_right_ipin_3.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_9.mux_l1_in_0__A1 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_45_ chany_top_in[8] chany_bottom_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_3.mux_l1_in_2_ chany_top_in[4] chany_bottom_in[4] mux_right_ipin_3.mux_l1_in_2_/S
+ mux_right_ipin_3.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_7.mux_l1_in_2__A1 chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_12.mux_l2_in_3_ _26_/HI chany_top_in[17] mux_right_ipin_12.mux_l2_in_0_/S
+ mux_right_ipin_12.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_59_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_8.mux_l3_in_0_ mux_right_ipin_8.mux_l2_in_1_/X mux_right_ipin_8.mux_l2_in_0_/X
+ mux_right_ipin_8.mux_l3_in_1_/S mux_right_ipin_8.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_28_ _28_/HI _28_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_10.mux_l1_in_0__A1 chany_bottom_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_7.mux_l2_in_1__A1 mux_right_ipin_7.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_8.mux_l2_in_1_ chany_bottom_in[13] mux_right_ipin_8.mux_l1_in_2_/X
+ mux_right_ipin_8.mux_l2_in_2_/S mux_right_ipin_8.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_12.mux_l4_in_0_ mux_right_ipin_12.mux_l3_in_1_/X mux_right_ipin_12.mux_l3_in_0_/X
+ mux_right_ipin_12.mux_l4_in_0_/S mux_right_ipin_12.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_ipin_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_5.mux_l2_in_3__A1 chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_1__S mux_right_ipin_0.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_4.mux_l1_in_0__A0 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_7.mux_l3_in_0__A1 mux_right_ipin_7.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_15.mux_l2_in_2__A0 chany_bottom_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_ipin_8.mux_l1_in_2_ chany_top_in[9] chany_bottom_in[9] mux_right_ipin_8.mux_l1_in_2_/S
+ mux_right_ipin_8.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_61_ chany_bottom_in[12] chany_top_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_ipin_3.mux_l2_in_0_ mux_right_ipin_3.mux_l1_in_1_/X mux_right_ipin_3.mux_l1_in_0_/X
+ mux_right_ipin_3.mux_l2_in_3_/S mux_right_ipin_3.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_12.mux_l3_in_1_ mux_right_ipin_12.mux_l2_in_3_/X mux_right_ipin_12.mux_l2_in_2_/X
+ mux_right_ipin_12.mux_l3_in_0_/S mux_right_ipin_12.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_15.mux_l3_in_1__A0 mux_right_ipin_15.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_44_ chany_top_in[9] chany_bottom_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_5.mux_l2_in_2__S mux_right_ipin_5.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_3_0_prog_clk_A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_3.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_3.mux_l1_in_2_/S
+ mux_right_ipin_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_12.mux_l2_in_2_ chany_bottom_in[17] chany_top_in[13] mux_right_ipin_12.mux_l2_in_0_/S
+ mux_right_ipin_12.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_2.mux_l2_in_1__A0 chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_9.mux_l3_in_0__S mux_right_ipin_9.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_27_ _27_/HI _27_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_15.mux_l4_in_0__A0 mux_right_ipin_15.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__34__A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_3__A0 _22_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_2.mux_l3_in_0__A0 mux_right_ipin_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_8.mux_l2_in_0_ mux_right_ipin_8.mux_l1_in_1_/X mux_right_ipin_8.mux_l1_in_0_/X
+ mux_right_ipin_8.mux_l2_in_2_/S mux_right_ipin_8.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_8.mux_l4_in_0__S mux_right_ipin_8.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_0__A1 chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_15.mux_l2_in_2__A1 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_8.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_8.mux_l1_in_2_/S
+ mux_right_ipin_8.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_53_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__42__A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_prog_clk clkbuf_2_0_0_prog_clk/A clkbuf_3_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
X_60_ chany_bottom_in[13] chany_top_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l3_in_0_ mux_right_ipin_12.mux_l2_in_1_/X mux_right_ipin_12.mux_l2_in_0_/X
+ mux_right_ipin_12.mux_l3_in_0_/S mux_right_ipin_12.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_13.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_12.mux_l2_in_2__S mux_right_ipin_12.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__37__A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_6.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l1_in_1__A0 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_15.mux_l3_in_1__A1 mux_right_ipin_15.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_43_ chany_top_in[10] chany_bottom_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_9.mux_l2_in_2__A0 chany_bottom_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_12.mux_l2_in_1_ chany_bottom_in[13] mux_right_ipin_12.mux_l1_in_2_/X
+ mux_right_ipin_12.mux_l2_in_0_/S mux_right_ipin_12.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_59_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_1__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_3.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_3.mux_l1_in_2_/S
+ mux_right_ipin_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_46_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26_ _26_/HI _26_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_15.mux_l4_in_0__A1 mux_right_ipin_15.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l2_in_0__A0 mux_right_ipin_12.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__50__A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_9.mux_l3_in_1__A0 mux_right_ipin_9.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_3__A1 chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_2.mux_l3_in_0__A1 mux_right_ipin_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_12.mux_l1_in_2_ chany_top_in[7] chany_bottom_in[7] mux_right_ipin_12.mux_l1_in_0_/S
+ mux_right_ipin_12.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_15.mux_l4_in_0__S mux_right_ipin_15.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_10.mux_l2_in_2__A0 chany_bottom_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__45__A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_14.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_9.mux_l4_in_0__A0 mux_right_ipin_9.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_0.mux_l3_in_1_/S mux_right_ipin_0.mux_l4_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_7.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_7.mux_l1_in_0__S mux_right_ipin_7.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_10.mux_l3_in_1__A0 mux_right_ipin_10.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_8.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_8.mux_l1_in_2_/S
+ mux_right_ipin_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_10.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__53__A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l1_in_1__A1 chany_bottom_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_43_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_10.mux_l4_in_0__A0 mux_right_ipin_10.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_42_ chany_top_in[11] chany_bottom_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_9.mux_l2_in_2__A1 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_6.mux_l2_in_0__S mux_right_ipin_6.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_12.mux_l2_in_0_ mux_right_ipin_12.mux_l1_in_1_/X mux_right_ipin_12.mux_l1_in_0_/X
+ mux_right_ipin_12.mux_l2_in_0_/S mux_right_ipin_12.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_59_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__48__A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25_ _25_/HI _25_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_12.mux_l4_in_0_/X left_grid_pin_28_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_ipin_12.mux_l2_in_0__A1 mux_right_ipin_12.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_1.mux_l2_in_2__S mux_right_ipin_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_9.mux_l3_in_1__A1 mux_right_ipin_9.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_4.mux_l4_in_0_/X left_grid_pin_20_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_2_0_prog_clk_A clkbuf_1_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_3.mux_l3_in_1_/S mux_right_ipin_3.mux_l4_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_35_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_12.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_12.mux_l1_in_0_/S
+ mux_right_ipin_12.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_5.mux_l3_in_0__S mux_right_ipin_5.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_10.mux_l2_in_2__A1 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__61__A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_13.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_6.mux_l2_in_0__A0 chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_9.mux_l4_in_0__A1 mux_right_ipin_9.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_14.mux_l1_in_0__S mux_right_ipin_14.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__56__A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_0.mux_l2_in_1_/S mux_right_ipin_0.mux_l3_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_6.mux_l2_in_3__S mux_right_ipin_6.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_10.mux_l3_in_1__A1 mux_right_ipin_10.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_4.mux_l4_in_0__S mux_right_ipin_4.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_4.mux_l2_in_2__A0 chany_bottom_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_13.mux_l2_in_0__S mux_right_ipin_13.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_10.mux_l4_in_0__A1 mux_right_ipin_10.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_41_ chany_top_in[12] chany_bottom_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_6.mux_l3_in_0_/S mux_right_ipin_6.mux_l4_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_4.mux_l3_in_1__A0 mux_right_ipin_4.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__64__A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24_ _24_/HI _24_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_11.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l3_in_0__S mux_right_ipin_12.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__59__A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_4.mux_l4_in_0__A0 mux_right_ipin_4.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_3.mux_l2_in_3_/S mux_right_ipin_3.mux_l3_in_1_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_ipin_12.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_12.mux_l1_in_0_/S
+ mux_right_ipin_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0__A mux_left_ipin_0.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_6.mux_l2_in_0__A1 mux_right_ipin_6.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_13.mux_l2_in_3__S mux_right_ipin_13.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_11.mux_l4_in_0__S mux_right_ipin_11.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_0.mux_l1_in_0_/S mux_right_ipin_0.mux_l2_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__72__A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_9.mux_l3_in_0_/S mux_right_ipin_9.mux_l4_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_4.mux_l2_in_2__A1 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__67__A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_14.mux_l2_in_1__A0 chany_bottom_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0__S mux_right_ipin_3.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_11.mux_l3_in_0_/S mux_right_ipin_11.mux_l4_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_40_ chany_top_in[13] chany_bottom_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0__S mux_left_ipin_0.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_6.mux_l2_in_0_/S mux_right_ipin_6.mux_l3_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_4.mux_l3_in_1__A1 mux_right_ipin_4.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_12.mux_l2_in_3__A0 _26_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_4.mux_l2_in_3_ _32_/HI chany_top_in[15] mux_right_ipin_4.mux_l2_in_0_/S
+ mux_right_ipin_4.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_14.mux_l3_in_0__A0 mux_right_ipin_14.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23_ _23_/HI _23_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0__S mux_right_ipin_2.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__75__A left_width_0_height_0__pin_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0__A0 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_4.mux_l4_in_0__A1 mux_right_ipin_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_3.mux_l1_in_2_/S mux_right_ipin_3.mux_l2_in_3_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_8.mux_l1_in_1__S mux_right_ipin_8.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_ipin_0.mux_l1_in_1__A0 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_1_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_4.mux_l4_in_0_ mux_right_ipin_4.mux_l3_in_1_/X mux_right_ipin_4.mux_l3_in_0_/X
+ mux_right_ipin_4.mux_l4_in_0_/S mux_right_ipin_4.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_1.mux_l3_in_0__S mux_right_ipin_1.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_ipin_0.mux_l4_in_0_/S mux_right_ipin_0.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_14.mux_l3_in_0_/S mux_right_ipin_14.mux_l4_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0__A0 mux_left_ipin_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_1__S mux_right_ipin_7.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_9.mux_l2_in_3_/S mux_right_ipin_9.mux_l3_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_9.mux_l2_in_3_ _20_/HI chany_top_in[14] mux_right_ipin_9.mux_l2_in_3_/S
+ mux_right_ipin_9.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_10.mux_l1_in_0__S mux_right_ipin_10.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1_0_prog_clk clkbuf_3_1_0_prog_clk/A clkbuf_3_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_4.mux_l3_in_1_ mux_right_ipin_4.mux_l2_in_3_/X mux_right_ipin_4.mux_l2_in_2_/X
+ mux_right_ipin_4.mux_l3_in_0_/S mux_right_ipin_4.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_14.mux_l2_in_1__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_2.mux_l2_in_3__S mux_right_ipin_2.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_11.mux_l2_in_0_/S mux_right_ipin_11.mux_l3_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_0.mux_l4_in_0__S mux_right_ipin_0.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_8.mux_l1_in_2__A0 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_6.mux_l1_in_0_/S mux_right_ipin_6.mux_l2_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_6.mux_l3_in_1__S mux_right_ipin_6.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_12.mux_l2_in_3__A1 chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_4.mux_l2_in_2_ chany_bottom_in[15] chany_top_in[9] mux_right_ipin_4.mux_l2_in_0_/S
+ mux_right_ipin_4.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_14.mux_l3_in_0__A1 mux_right_ipin_14.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_11.mux_l1_in_0__A0 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22_ _22_/HI _22_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_8.mux_l2_in_1__A0 chany_bottom_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_ipin_9.mux_l4_in_0_ mux_right_ipin_9.mux_l3_in_1_/X mux_right_ipin_9.mux_l3_in_0_/X
+ mux_right_ipin_9.mux_l4_in_0_/S mux_right_ipin_9.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_15.mux_l1_in_1__S mux_right_ipin_15.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0__A1 mux_right_ipin_1.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_2.mux_l4_in_0_/S mux_right_ipin_3.mux_l1_in_2_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_6.mux_l2_in_3__A0 _17_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_ipin_0.mux_l1_in_1__A1 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_12.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_8.mux_l3_in_0__A0 mux_right_ipin_8.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_9.mux_l3_in_1_ mux_right_ipin_9.mux_l2_in_3_/X mux_right_ipin_9.mux_l2_in_2_/X
+ mux_right_ipin_9.mux_l3_in_0_/S mux_right_ipin_9.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_14.mux_l2_in_1__S mux_right_ipin_14.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_14.mux_l2_in_3_/S mux_right_ipin_14.mux_l3_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0__A1 mux_left_ipin_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_9.mux_l1_in_0_/S mux_right_ipin_9.mux_l2_in_3_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_9.mux_l2_in_2_ chany_bottom_in[14] chany_top_in[6] mux_right_ipin_9.mux_l2_in_3_/S
+ mux_right_ipin_9.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_4.mux_l3_in_0_ mux_right_ipin_4.mux_l2_in_1_/X mux_right_ipin_4.mux_l2_in_0_/X
+ mux_right_ipin_4.mux_l3_in_0_/S mux_right_ipin_4.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_11.mux_l1_in_0_/S mux_right_ipin_11.mux_l2_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_8.mux_l1_in_2__A1 chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_13.mux_l3_in_1__S mux_right_ipin_13.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_5.mux_l4_in_0_/S mux_right_ipin_6.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_11.mux_l1_in_0__A1 chany_bottom_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_40_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_4.mux_l2_in_1_ chany_bottom_in[9] mux_right_ipin_4.mux_l1_in_2_/X
+ mux_right_ipin_4.mux_l2_in_0_/S mux_right_ipin_4.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_21_ _21_/HI _21_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_27_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_13.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_8.mux_l2_in_1__A1 mux_right_ipin_8.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_6.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_15.mux_l4_in_0_/X left_grid_pin_31_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_ipin_13.mux_l2_in_3_ _27_/HI chany_top_in[18] mux_right_ipin_13.mux_l2_in_2_/S
+ mux_right_ipin_13.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_6.mux_l2_in_3__A1 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_4.mux_l1_in_2_ chany_top_in[5] chany_bottom_in[5] mux_right_ipin_4.mux_l1_in_1_/S
+ mux_right_ipin_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_7.mux_l4_in_0_/X left_grid_pin_23_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_5.mux_l1_in_0__A0 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_8.mux_l3_in_0__A1 mux_right_ipin_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_9.mux_l3_in_0_ mux_right_ipin_9.mux_l2_in_1_/X mux_right_ipin_9.mux_l2_in_0_/X
+ mux_right_ipin_9.mux_l3_in_0_/S mux_right_ipin_9.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_4.mux_l1_in_1__S mux_right_ipin_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_14.mux_l1_in_0_/S mux_right_ipin_14.mux_l2_in_3_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_2__A0 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_8.mux_l4_in_0_/S mux_right_ipin_9.mux_l1_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_9.mux_l2_in_1_ chany_bottom_in[6] chany_top_in[2] mux_right_ipin_9.mux_l2_in_3_/S
+ mux_right_ipin_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_13.mux_l4_in_0_ mux_right_ipin_13.mux_l3_in_1_/X mux_right_ipin_13.mux_l3_in_0_/X
+ mux_right_ipin_13.mux_l4_in_0_/S mux_right_ipin_13.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_10.mux_l4_in_0_/S mux_right_ipin_11.mux_l1_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_3.mux_l2_in_1__S mux_right_ipin_3.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.mux_l2_in_1__A0 chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_ipin_0.mux_l2_in_1__S mux_left_ipin_0.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_13.mux_l3_in_1_ mux_right_ipin_13.mux_l2_in_3_/X mux_right_ipin_13.mux_l2_in_2_/X
+ mux_right_ipin_13.mux_l3_in_1_/S mux_right_ipin_13.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_4.mux_l2_in_0_ mux_right_ipin_4.mux_l1_in_1_/X mux_right_ipin_4.mux_l1_in_0_/X
+ mux_right_ipin_4.mux_l2_in_0_/S mux_right_ipin_4.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_20_ _20_/HI _20_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_ipin_1.mux_l2_in_3__A0 _23_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_3.mux_l3_in_0__A0 mux_right_ipin_3.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_2.mux_l3_in_1__S mux_right_ipin_2.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_8.mux_l2_in_2__S mux_right_ipin_8.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_13.mux_l2_in_2_ chany_bottom_in[18] chany_top_in[10] mux_right_ipin_13.mux_l2_in_2_/S
+ mux_right_ipin_13.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_4_0_prog_clk_A clkbuf_3_5_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_4.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_4.mux_l1_in_1_/S
+ mux_right_ipin_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_11.mux_l1_in_1__S mux_right_ipin_11.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_5.mux_l1_in_0__A1 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_ipin_0.mux_l2_in_3__A0 _21_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_13.mux_l4_in_0_/S mux_right_ipin_14.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_3.mux_l1_in_2__A1 chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_ipin_9.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_9.mux_l1_in_0_/X
+ mux_right_ipin_9.mux_l2_in_3_/S mux_right_ipin_9.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_ipin_10.mux_l2_in_1__S mux_right_ipin_10.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_10.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_3.mux_l2_in_1__A1 mux_right_ipin_3.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_13.mux_l2_in_0__A0 chany_bottom_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_2.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_prog_clk clkbuf_3_1_0_prog_clk/A clkbuf_3_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_13.mux_l3_in_0_ mux_right_ipin_13.mux_l2_in_1_/X mux_right_ipin_13.mux_l2_in_0_/X
+ mux_right_ipin_13.mux_l3_in_1_/S mux_right_ipin_13.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_3__A1 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0__A0 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_3.mux_l3_in_0__A1 mux_right_ipin_3.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_15.mux_l2_in_2__S mux_right_ipin_15.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_11.mux_l2_in_2__A0 chany_bottom_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_13.mux_l2_in_1_ chany_bottom_in[10] chany_top_in[2] mux_right_ipin_13.mux_l2_in_2_/S
+ mux_right_ipin_13.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_4.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_4.mux_l1_in_1_/S
+ mux_right_ipin_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_11.mux_l3_in_1__A0 mux_right_ipin_11.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_3__A1 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_5.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1__S mux_right_ipin_0.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_0.mux_l4_in_0_/X left_grid_pin_16_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_11.mux_l4_in_0__A0 mux_right_ipin_11.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_ipin_9.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_9.mux_l1_in_0_/S
+ mux_right_ipin_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_13.mux_l2_in_0__A1 mux_right_ipin_13.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_7.mux_l1_in_1__A0 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_0__A1 chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_11.mux_l2_in_2__A1 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_9.mux_l2_in_0__S mux_right_ipin_9.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_13.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_13.mux_l1_in_0_/X
+ mux_right_ipin_13.mux_l2_in_2_/S mux_right_ipin_13.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_7.mux_l2_in_0__A0 mux_right_ipin_7.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_8.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_11.mux_l3_in_1__A1 mux_right_ipin_11.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_4.mux_l2_in_2__S mux_right_ipin_4.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_5.mux_l2_in_2__A0 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_3_0_prog_clk_A clkbuf_1_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_8.mux_l3_in_0__S mux_right_ipin_8.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_11.mux_l4_in_0__A1 mux_right_ipin_11.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_5.mux_l3_in_1__A0 mux_right_ipin_5.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_9.mux_l2_in_3__S mux_right_ipin_9.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_7.mux_l4_in_0__S mux_right_ipin_7.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_7.mux_l1_in_1__A1 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l1_in_2__S mux_right_ipin_12.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_11.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_5.mux_l4_in_0__A0 mux_right_ipin_5.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_77_ gfpga_pad_EMBEDDED_IO_SOC_IN left_width_0_height_0__pin_1_upper VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_7.mux_l2_in_0__A1 mux_right_ipin_7.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_15.mux_l1_in_2__A0 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_11.mux_l2_in_2__S mux_right_ipin_11.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_15.mux_l3_in_0__S mux_right_ipin_15.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_5.mux_l2_in_2__A1 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_13.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_13.mux_l1_in_0_/S
+ mux_right_ipin_13.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_15.mux_l2_in_1__A0 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_27_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_12.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_0.mux_l2_in_3_ _22_/HI chany_top_in[17] mux_right_ipin_0.mux_l2_in_1_/S
+ mux_right_ipin_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_5.mux_l3_in_1__A1 mux_right_ipin_5.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_13.mux_l2_in_3__A0 _27_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_14.mux_l4_in_0__S mux_right_ipin_14.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_5.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_ipin_15.mux_l3_in_0__A0 mux_right_ipin_15.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D ccff_head VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_2.mux_l2_in_0__A0 chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_5.mux_l4_in_0__A1 mux_right_ipin_5.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_76_ gfpga_pad_EMBEDDED_IO_SOC_IN left_width_0_height_0__pin_1_lower VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0__S mux_right_ipin_6.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_0.mux_l4_in_0_ mux_right_ipin_0.mux_l3_in_1_/X mux_right_ipin_0.mux_l3_in_0_/X
+ mux_right_ipin_0.mux_l4_in_0_/S mux_right_ipin_0.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_2__A0 chany_bottom_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_59_ chany_bottom_in[14] chany_top_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_15.mux_l1_in_2__A1 chany_bottom_in[4] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_ipin_5.mux_l2_in_3_ _33_/HI chany_top_in[18] mux_right_ipin_5.mux_l2_in_3_/S
+ mux_right_ipin_5.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_ipin_0.mux_l3_in_1_ mux_right_ipin_0.mux_l2_in_3_/X mux_right_ipin_0.mux_l2_in_2_/X
+ mux_right_ipin_0.mux_l3_in_1_/S mux_right_ipin_0.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_5.mux_l2_in_0__S mux_right_ipin_5.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_ipin_0.mux_l3_in_1__A0 mux_right_ipin_0.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_15.mux_l2_in_1__A1 mux_right_ipin_15.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D mux_left_ipin_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_2__S mux_right_ipin_0.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_0.mux_l2_in_2_ chany_bottom_in[17] chany_top_in[11] mux_right_ipin_0.mux_l2_in_1_/S
+ mux_right_ipin_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_0.mux_l4_in_0__A0 mux_right_ipin_0.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_5.mux_l4_in_0_ mux_right_ipin_5.mux_l3_in_1_/X mux_right_ipin_5.mux_l3_in_0_/X
+ mux_right_ipin_5.mux_l4_in_0_/S mux_right_ipin_5.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_4.mux_l3_in_0__S mux_right_ipin_4.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mux_right_ipin_15.mux_l4_in_0_/S ccff_tail clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_13.mux_l2_in_3__A1 chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_12.mux_l1_in_0__A0 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_15.mux_l3_in_0__A1 mux_right_ipin_15.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_9.mux_l2_in_1__A0 chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_13.mux_l1_in_0__S mux_right_ipin_13.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_2.mux_l2_in_0__A1 mux_right_ipin_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_5.mux_l3_in_1_ mux_right_ipin_5.mux_l2_in_3_/X mux_right_ipin_5.mux_l2_in_2_/X
+ mux_right_ipin_5.mux_l3_in_1_/S mux_right_ipin_5.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_75_ left_width_0_height_0__pin_0_ gfpga_pad_EMBEDDED_IO_SOC_OUT VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__buf_2
XFILLER_51_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_5.mux_l2_in_3__S mux_right_ipin_5.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_3.mux_l4_in_0__S mux_right_ipin_3.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_7.mux_l2_in_3__A0 _18_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__40__A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_ipin_0.mux_l4_in_0__S mux_left_ipin_0.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_9.mux_l3_in_0__A0 mux_right_ipin_9.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_2__A1 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_9.mux_l3_in_1__S mux_right_ipin_9.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_58_ chany_bottom_in[15] chany_top_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_5.mux_l2_in_2_ chany_bottom_in[18] chany_top_in[10] mux_right_ipin_5.mux_l2_in_3_/S
+ mux_right_ipin_5.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_10.mux_l2_in_1__A0 chany_bottom_in[7] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l2_in_0__S mux_right_ipin_12.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__35__A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_ipin_0.mux_l3_in_0_ mux_right_ipin_0.mux_l2_in_1_/X mux_right_ipin_0.mux_l2_in_0_/X
+ mux_right_ipin_0.mux_l3_in_1_/S mux_right_ipin_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_0.mux_l3_in_1__A1 mux_right_ipin_0.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_10.mux_l3_in_0__A0 mux_right_ipin_10.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_11.mux_l4_in_0_/X left_grid_pin_27_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_11.mux_l3_in_0__S mux_right_ipin_11.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_0.mux_l2_in_1_ chany_bottom_in[11] mux_right_ipin_0.mux_l1_in_2_/X
+ mux_right_ipin_0.mux_l2_in_1_/S mux_right_ipin_0.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_0.mux_l4_in_0__A1 mux_right_ipin_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_3.mux_l4_in_0_/X left_grid_pin_19_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_57_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__43__A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l1_in_0__A1 chany_bottom_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_9.mux_l2_in_1__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_ipin_0.mux_l1_in_2_ chany_top_in[5] chany_bottom_in[5] mux_right_ipin_0.mux_l1_in_0_/S
+ mux_right_ipin_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__38__A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l2_in_3__S mux_right_ipin_12.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_10.mux_l4_in_0__S mux_right_ipin_10.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_5.mux_l3_in_0_ mux_right_ipin_5.mux_l2_in_1_/X mux_right_ipin_5.mux_l2_in_0_/X
+ mux_right_ipin_5.mux_l3_in_1_/S mux_right_ipin_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_74_ ccff_tail gfpga_pad_EMBEDDED_IO_SOC_DIR VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_7.mux_l2_in_3__A1 chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_6.mux_l1_in_0__A0 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_9.mux_l3_in_0__A1 mux_right_ipin_9.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_57_ chany_bottom_in[16] chany_top_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0__S mux_right_ipin_2.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_5.mux_l2_in_1_ chany_bottom_in[10] chany_top_in[2] mux_right_ipin_5.mux_l2_in_3_/S
+ mux_right_ipin_5.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_62_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_10.mux_l2_in_1__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__51__A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_4.mux_l1_in_2__A0 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__46__A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_14.mux_l2_in_3_ _28_/HI chany_top_in[19] mux_right_ipin_14.mux_l2_in_3_/S
+ mux_right_ipin_14.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_10.mux_l3_in_0__A1 mux_right_ipin_10.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0__S mux_right_ipin_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_4.mux_l2_in_1__A0 chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_0.mux_l2_in_0_ mux_right_ipin_0.mux_l1_in_1_/X mux_right_ipin_0.mux_l1_in_0_/X
+ mux_right_ipin_0.mux_l2_in_1_/S mux_right_ipin_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_7.mux_l1_in_1__S mux_right_ipin_7.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_2.mux_l2_in_3__A0 _30_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_2.mux_l3_in_1_/S mux_right_ipin_2.mux_l4_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_4.mux_l3_in_0__A0 mux_right_ipin_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_ipin_0.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_0.mux_l1_in_0_/S
+ mux_right_ipin_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_0_0_prog_clk_A clkbuf_3_1_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_0.mux_l3_in_0__S mux_right_ipin_0.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__54__A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_14.mux_l4_in_0_ mux_right_ipin_14.mux_l3_in_1_/X mux_right_ipin_14.mux_l3_in_0_/X
+ mux_right_ipin_14.mux_l4_in_0_/S mux_right_ipin_14.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_73_ chany_bottom_in[0] chany_top_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_6.mux_l2_in_1__S mux_right_ipin_6.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_12.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__49__A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0__A1 chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_56_ chany_bottom_in[17] chany_top_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_ipin_14.mux_l3_in_1_ mux_right_ipin_14.mux_l2_in_3_/X mux_right_ipin_14.mux_l2_in_2_/X
+ mux_right_ipin_14.mux_l3_in_0_/S mux_right_ipin_14.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_5.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_5.mux_l1_in_0_/X
+ mux_right_ipin_5.mux_l2_in_3_/S mux_right_ipin_5.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_3__S mux_right_ipin_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_4.mux_l1_in_2__A1 chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_39_ chany_top_in[14] chany_bottom_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_5.mux_l3_in_1__S mux_right_ipin_5.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__62__A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_14.mux_l2_in_2_ chany_bottom_in[19] chany_top_in[11] mux_right_ipin_14.mux_l2_in_3_/S
+ mux_right_ipin_14.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_5_0_prog_clk_A clkbuf_3_5_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_5.mux_l3_in_1_/S mux_right_ipin_5.mux_l4_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_4.mux_l2_in_1__A1 mux_right_ipin_4.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_10.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__57__A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_14.mux_l2_in_0__A0 chany_bottom_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_15.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_3__A1 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0__A0 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_2.mux_l2_in_3_/S mux_right_ipin_2.mux_l3_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_4.mux_l3_in_0__A1 mux_right_ipin_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_0.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_0.mux_l1_in_0_/S
+ mux_right_ipin_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_12.mux_l2_in_2__A0 chany_bottom_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_60_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_13.mux_l2_in_1__S mux_right_ipin_13.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__70__A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_72_ chany_bottom_in[1] chany_top_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__65__A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_55_ chany_bottom_in[18] chany_top_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_12.mux_l3_in_1__A0 mux_right_ipin_12.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_14.mux_l3_in_0_ mux_right_ipin_14.mux_l2_in_1_/X mux_right_ipin_14.mux_l2_in_0_/X
+ mux_right_ipin_14.mux_l3_in_0_/S mux_right_ipin_14.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_0__A0 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_8.mux_l3_in_1_/S mux_right_ipin_8.mux_l4_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_62_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_11.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l3_in_1__S mux_right_ipin_12.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_38_ chany_top_in[15] chany_bottom_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_12.mux_l4_in_0__A0 mux_right_ipin_12.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_10.mux_l3_in_1_/S mux_right_ipin_10.mux_l4_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_14.mux_l2_in_1_ chany_bottom_in[11] chany_top_in[3] mux_right_ipin_14.mux_l2_in_3_/S
+ mux_right_ipin_14.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_5.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_5.mux_l1_in_0_/S
+ mux_right_ipin_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_5.mux_l2_in_3_/S mux_right_ipin_5.mux_l3_in_1_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__73__A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_ipin_14.mux_l2_in_0__A1 mux_right_ipin_14.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_8.mux_l1_in_1__A0 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__68__A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_1.mux_l1_in_0__A1 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_2.mux_l1_in_0_/S mux_right_ipin_2.mux_l2_in_3_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_1__S mux_right_ipin_3.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l2_in_2__A1 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1__S mux_left_ipin_0.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_71_ chany_bottom_in[2] chany_top_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_8.mux_l2_in_0__A0 mux_right_ipin_8.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_13.mux_l3_in_1_/S mux_right_ipin_13.mux_l4_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_54_ chany_bottom_in[19] chany_top_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_12.mux_l3_in_1__A1 mux_right_ipin_12.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_6.mux_l2_in_2__A0 chany_bottom_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_0__A1 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_1__S mux_right_ipin_2.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_8.mux_l2_in_2_/S mux_right_ipin_8.mux_l3_in_1_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__76__A gfpga_pad_EMBEDDED_IO_SOC_IN VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_8.mux_l1_in_2__S mux_right_ipin_8.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_37_ chany_top_in[16] chany_bottom_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_10.mux_l2_in_2_/S mux_right_ipin_10.mux_l3_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_12.mux_l4_in_0__A1 mux_right_ipin_12.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_14.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_14.mux_l1_in_0_/X
+ mux_right_ipin_14.mux_l2_in_3_/S mux_right_ipin_14.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_6.mux_l3_in_1__A0 mux_right_ipin_6.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_5.mux_l1_in_0_/S mux_right_ipin_5.mux_l2_in_3_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_43_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_1.mux_l3_in_1__S mux_right_ipin_1.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_7.mux_l2_in_2__S mux_right_ipin_7.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_14.mux_l4_in_0_/X left_grid_pin_30_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_57_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_8.mux_l1_in_1__A1 chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_6.mux_l4_in_0__A0 mux_right_ipin_6.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_6.mux_l4_in_0_/X left_grid_pin_22_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_39_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_1.mux_l4_in_0_/S mux_right_ipin_2.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_70_ chany_bottom_in[3] chany_top_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_8.mux_l2_in_0__A1 mux_right_ipin_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_13.mux_l2_in_2_/S mux_right_ipin_13.mux_l3_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_53_ chany_top_in[0] chany_bottom_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_6.mux_l2_in_2__A1 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_15.mux_l1_in_2__S mux_right_ipin_15.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_8.mux_l1_in_2_/S mux_right_ipin_8.mux_l2_in_2_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_36_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36_ chany_top_in[17] chany_bottom_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_10.mux_l1_in_0_/S mux_right_ipin_10.mux_l2_in_2_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_1__A0 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_6.mux_l3_in_1__A1 mux_right_ipin_6.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_4.mux_l4_in_0_/S mux_right_ipin_5.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_19_ _19_/HI _19_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_ipin_14.mux_l2_in_3__A0 _28_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_14.mux_l2_in_2__S mux_right_ipin_14.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_6.mux_l4_in_0__A1 mux_right_ipin_6.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.mux_l2_in_0__A0 mux_right_ipin_3.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_14.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_14.mux_l1_in_0_/S
+ mux_right_ipin_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_1.mux_l2_in_3_ _23_/HI chany_top_in[14] mux_right_ipin_1.mux_l2_in_0_/S
+ mux_right_ipin_1.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_2__A0 chany_bottom_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_13.mux_l1_in_0_/S mux_right_ipin_13.mux_l2_in_2_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_52_ chany_top_in[1] chany_bottom_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_7.mux_l4_in_0_/S mux_right_ipin_8.mux_l1_in_2_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_1.mux_l3_in_1__A0 mux_right_ipin_1.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_9.mux_l1_in_0__S mux_right_ipin_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_35_ chany_top_in[18] chany_bottom_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_ipin_1.mux_l4_in_0_ mux_right_ipin_1.mux_l3_in_1_/X mux_right_ipin_1.mux_l3_in_0_/X
+ mux_right_ipin_1.mux_l4_in_0_/S mux_right_ipin_1.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_ipin_0.mux_l2_in_2__A0 chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_9.mux_l4_in_0_/S mux_right_ipin_10.mux_l1_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_3.mux_l1_in_1__A1 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_1.mux_l4_in_0__A0 mux_right_ipin_1.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_18_ _18_/HI _18_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_ipin_14.mux_l2_in_3__A1 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_6.mux_l2_in_3_ _17_/HI chany_top_in[19] mux_right_ipin_6.mux_l2_in_0_/S
+ mux_right_ipin_6.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_4.mux_l1_in_2__S mux_right_ipin_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_13.mux_l1_in_0__A0 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_ipin_0.mux_l3_in_1__A0 mux_left_ipin_0.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_1.mux_l3_in_1_ mux_right_ipin_1.mux_l2_in_3_/X mux_right_ipin_1.mux_l2_in_2_/X
+ mux_right_ipin_1.mux_l3_in_0_/S mux_right_ipin_1.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_8.mux_l2_in_0__S mux_right_ipin_8.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_0__A1 mux_right_ipin_3.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_11.mux_l1_in_2__A0 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_left_ipin_0.mux_l3_in_1_/S mux_left_ipin_0.mux_l4_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_8.mux_l2_in_3__A0 _19_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.mux_l2_in_2__S mux_right_ipin_3.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_ipin_0.mux_l4_in_0__A0 mux_left_ipin_0.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_1.mux_l2_in_2_ chany_bottom_in[14] chany_top_in[6] mux_right_ipin_1.mux_l2_in_0_/S
+ mux_right_ipin_1.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_2__A1 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_2__S mux_left_ipin_0.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_6.mux_l4_in_0_ mux_right_ipin_6.mux_l3_in_1_/X mux_right_ipin_6.mux_l3_in_0_/X
+ mux_right_ipin_6.mux_l4_in_0_/S mux_right_ipin_6.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_7.mux_l3_in_0__S mux_right_ipin_7.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_11.mux_l2_in_1__A0 chany_bottom_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_12.mux_l4_in_0_/S mux_right_ipin_13.mux_l1_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_51_ chany_top_in[2] chany_bottom_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_1.mux_l3_in_1__A1 mux_right_ipin_1.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_6.mux_l3_in_1_ mux_right_ipin_6.mux_l2_in_3_/X mux_right_ipin_6.mux_l2_in_2_/X
+ mux_right_ipin_6.mux_l3_in_0_/S mux_right_ipin_6.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34_ chany_top_in[19] chany_bottom_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_8.mux_l2_in_3__S mux_right_ipin_8.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_11.mux_l3_in_0__A0 mux_right_ipin_11.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_2__A1 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_6.mux_l4_in_0__S mux_right_ipin_6.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_11.mux_l1_in_2__S mux_right_ipin_11.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_1.mux_l4_in_0__A1 mux_right_ipin_1.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17_ _17_/HI _17_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_right_ipin_6.mux_l2_in_2_ chany_bottom_in[19] chany_top_in[11] mux_right_ipin_6.mux_l2_in_0_/S
+ mux_right_ipin_6.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_15.mux_l2_in_0__S mux_right_ipin_15.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_13.mux_l1_in_0__A1 chany_bottom_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_1.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_1.mux_l3_in_0_ mux_right_ipin_1.mux_l2_in_1_/X mux_right_ipin_1.mux_l2_in_0_/X
+ mux_right_ipin_1.mux_l3_in_0_/S mux_right_ipin_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_ipin_0.mux_l3_in_1__A1 mux_left_ipin_0.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_10.mux_l2_in_2__S mux_right_ipin_10.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_11.mux_l1_in_2__A1 chany_bottom_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_ipin_0.mux_l2_in_0_/S mux_left_ipin_0.mux_l3_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_8.mux_l2_in_3__A1 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_10.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_1.mux_l2_in_1_ chany_bottom_in[6] chany_top_in[2] mux_right_ipin_1.mux_l2_in_0_/S
+ mux_right_ipin_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_14.mux_l3_in_0__S mux_right_ipin_14.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_ipin_0.mux_l4_in_0__A1 mux_left_ipin_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_7.mux_l1_in_0__A0 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_11.mux_l2_in_1__A1 mux_right_ipin_11.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_50_ chany_top_in[3] chany_bottom_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_ipin_10.mux_l2_in_3_ _24_/HI chany_top_in[15] mux_right_ipin_10.mux_l2_in_2_/S
+ mux_right_ipin_10.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_15.mux_l2_in_3__S mux_right_ipin_15.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_13.mux_l4_in_0__S mux_right_ipin_13.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_6.mux_l3_in_0_ mux_right_ipin_6.mux_l2_in_1_/X mux_right_ipin_6.mux_l2_in_0_/X
+ mux_right_ipin_6.mux_l3_in_0_/S mux_right_ipin_6.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_4.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33_ _33_/HI _33_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_ipin_11.mux_l3_in_0__A1 mux_right_ipin_11.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_15.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_ipin_5.mux_l2_in_1__A0 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_8.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_ipin_6.mux_l2_in_1_ chany_bottom_in[11] chany_top_in[3] mux_right_ipin_6.mux_l2_in_0_/S
+ mux_right_ipin_6.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_5.mux_l1_in_0__S mux_right_ipin_5.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_10.mux_l4_in_0_ mux_right_ipin_10.mux_l3_in_1_/X mux_right_ipin_10.mux_l3_in_0_/X
+ mux_right_ipin_10.mux_l4_in_0_/S mux_right_ipin_10.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.mux_l2_in_3__A0 _31_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_5.mux_l3_in_0__A0 mux_right_ipin_5.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_0.mux_l1_in_2__S mux_right_ipin_0.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l2_in_3_ _29_/HI chany_top_in[16] mux_right_ipin_15.mux_l2_in_0_/S
+ mux_right_ipin_15.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_ipin_0.mux_l1_in_2_/S mux_left_ipin_0.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_4.mux_l2_in_0__S mux_right_ipin_4.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_10.mux_l3_in_1_ mux_right_ipin_10.mux_l2_in_3_/X mux_right_ipin_10.mux_l2_in_2_/X
+ mux_right_ipin_10.mux_l3_in_1_/S mux_right_ipin_10.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_1.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_1.mux_l1_in_0_/X
+ mux_right_ipin_1.mux_l2_in_0_/S mux_right_ipin_1.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_7.mux_l1_in_0__A1 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_9.mux_l4_in_0_/X left_grid_pin_25_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xclkbuf_3_7_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_7.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_10.mux_l2_in_2_ chany_bottom_in[15] chany_top_in[7] mux_right_ipin_10.mux_l2_in_2_/S
+ mux_right_ipin_10.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_1_0_prog_clk_A clkbuf_3_1_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_3.mux_l3_in_0__S mux_right_ipin_3.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_15.mux_l1_in_1__A0 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_15.mux_l4_in_0_ mux_right_ipin_15.mux_l3_in_1_/X mux_right_ipin_15.mux_l3_in_0_/X
+ mux_right_ipin_15.mux_l4_in_0_/S mux_right_ipin_15.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_ipin_0.mux_l3_in_0__S mux_left_ipin_0.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_32_ _32_/HI _32_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_ipin_9.mux_l2_in_1__S mux_right_ipin_9.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_5.mux_l2_in_1__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_12.mux_l1_in_0__S mux_right_ipin_12.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_15.mux_l2_in_0__A0 mux_right_ipin_15.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_15.mux_l3_in_1_ mux_right_ipin_15.mux_l2_in_3_/X mux_right_ipin_15.mux_l2_in_2_/X
+ mux_right_ipin_15.mux_l3_in_0_/S mux_right_ipin_15.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_6.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_6.mux_l1_in_0_/X
+ mux_right_ipin_6.mux_l2_in_0_/S mux_right_ipin_6.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_4.mux_l2_in_3__S mux_right_ipin_4.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_2.mux_l4_in_0__S mux_right_ipin_2.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_3.mux_l2_in_3__A1 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_2.mux_l1_in_0__A0 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_5.mux_l3_in_0__A1 mux_right_ipin_5.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_8.mux_l3_in_1__S mux_right_ipin_8.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_13.mux_l2_in_2__A0 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_11.mux_l2_in_0__S mux_right_ipin_11.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_ipin_15.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[10] mux_right_ipin_15.mux_l2_in_0_/S
+ mux_right_ipin_15.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_6_0_prog_clk_A clkbuf_3_7_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_left_ipin_0.mux_l1_in_2_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_0.mux_l1_in_2__A0 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_10.mux_l3_in_0_ mux_right_ipin_10.mux_l2_in_1_/X mux_right_ipin_10.mux_l2_in_0_/X
+ mux_right_ipin_10.mux_l3_in_1_/S mux_right_ipin_10.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_13.mux_l3_in_1__A0 mux_right_ipin_13.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_10.mux_l3_in_0__S mux_right_ipin_10.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_1__A0 chany_bottom_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_10.mux_l2_in_1_ chany_bottom_in[7] chany_top_in[3] mux_right_ipin_10.mux_l2_in_2_/S
+ mux_right_ipin_10.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_1.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_1.mux_l1_in_0_/S
+ mux_right_ipin_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_15.mux_l1_in_1__A1 chany_bottom_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_13.mux_l4_in_0__A0 mux_right_ipin_13.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31_ _31_/HI _31_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_0.mux_l3_in_0__A0 mux_right_ipin_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_11.mux_l2_in_3__S mux_right_ipin_11.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_15.mux_l2_in_0__A1 mux_right_ipin_15.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_15.mux_l3_in_0_ mux_right_ipin_15.mux_l2_in_1_/X mux_right_ipin_15.mux_l2_in_0_/X
+ mux_right_ipin_15.mux_l3_in_0_/S mux_right_ipin_15.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_15.mux_l3_in_1__S mux_right_ipin_15.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_ipin_2.mux_l1_in_0__A1 chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_13.mux_l2_in_2__A1 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_1.mux_l1_in_0__S mux_right_ipin_1.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_15.mux_l2_in_1_ chany_bottom_in[10] mux_right_ipin_15.mux_l1_in_2_/X
+ mux_right_ipin_15.mux_l2_in_0_/S mux_right_ipin_15.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_6.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_6.mux_l1_in_0_/S
+ mux_right_ipin_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_62_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_9.mux_l2_in_0__A0 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_ipin_0.mux_l2_in_3_ _21_/HI chany_top_in[16] mux_left_ipin_0.mux_l2_in_0_/S
+ mux_left_ipin_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_0.mux_l1_in_2__A1 chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_13.mux_l3_in_1__A1 mux_right_ipin_13.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_2__A0 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_15.mux_l1_in_2_ chany_top_in[4] chany_bottom_in[4] mux_right_ipin_15.mux_l1_in_0_/S
+ mux_right_ipin_15.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_0__S mux_right_ipin_0.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_0.mux_l2_in_1__A1 mux_right_ipin_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_10.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_10.mux_l1_in_0_/X
+ mux_right_ipin_10.mux_l2_in_2_/S mux_right_ipin_10.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_10.mux_l4_in_0_/X left_grid_pin_26_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_10.mux_l2_in_0__A0 chany_bottom_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_13.mux_l4_in_0__A1 mux_right_ipin_13.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_ipin_0.mux_l4_in_0_ mux_left_ipin_0.mux_l3_in_1_/X mux_left_ipin_0.mux_l3_in_0_/X
+ mux_left_ipin_0.mux_l4_in_0_/S mux_left_ipin_0.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_2.mux_l4_in_0_/X left_grid_pin_18_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_30_ _30_/HI _30_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_ipin_7.mux_l3_in_1__A0 mux_right_ipin_7.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0_0_prog_clk_A clkbuf_2_0_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_0.mux_l3_in_0__A1 mux_right_ipin_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_5.mux_l2_in_1__S mux_right_ipin_5.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_ipin_0.mux_l3_in_1_ mux_left_ipin_0.mux_l2_in_3_/X mux_left_ipin_0.mux_l2_in_2_/X
+ mux_left_ipin_0.mux_l3_in_1_/S mux_left_ipin_0.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_7.mux_l4_in_0__A0 mux_right_ipin_7.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_3__S mux_right_ipin_0.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_15.mux_l2_in_0_ mux_right_ipin_15.mux_l1_in_1_/X mux_right_ipin_15.mux_l1_in_0_/X
+ mux_right_ipin_15.mux_l2_in_0_/S mux_right_ipin_15.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_9.mux_l2_in_0__A1 mux_right_ipin_9.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_ipin_0.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[10] mux_left_ipin_0.mux_l2_in_0_/S
+ mux_left_ipin_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_4.mux_l3_in_1__S mux_right_ipin_4.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_7.mux_l2_in_2__A1 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_15.mux_l1_in_0_/S
+ mux_right_ipin_15.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_10.mux_l2_in_0__A1 mux_right_ipin_10.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__41__A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1__A0 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_7.mux_l3_in_1__A1 mux_right_ipin_7.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_15.mux_l2_in_3__A0 _29_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__36__A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l2_in_1__S mux_right_ipin_12.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_10.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_10.mux_l1_in_0_/S
+ mux_right_ipin_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_ipin_0.mux_l3_in_0_ mux_left_ipin_0.mux_l2_in_1_/X mux_left_ipin_0.mux_l2_in_0_/X
+ mux_left_ipin_0.mux_l3_in_1_/S mux_left_ipin_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_4.mux_l2_in_0__A0 mux_right_ipin_4.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_7.mux_l4_in_0__A1 mux_right_ipin_7.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_2.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_11.mux_l3_in_1__S mux_right_ipin_11.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_2__A0 chany_bottom_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_ipin_0.mux_l2_in_1_ chany_bottom_in[10] mux_left_ipin_0.mux_l1_in_2_/X mux_left_ipin_0.mux_l2_in_0_/S
+ mux_left_ipin_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__44__A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_15.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_15.mux_l1_in_0_/S
+ mux_right_ipin_15.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_2.mux_l3_in_1__A0 mux_right_ipin_2.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__39__A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_ipin_0.mux_l1_in_2_ chany_top_in[4] chany_bottom_in[4] mux_left_ipin_0.mux_l1_in_2_/S
+ mux_left_ipin_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_7.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_2.mux_l2_in_3_ _30_/HI chany_top_in[15] mux_right_ipin_2.mux_l2_in_3_/S
+ mux_right_ipin_2.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_4.mux_l1_in_1__A1 chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_2.mux_l4_in_0__A0 mux_right_ipin_2.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_15.mux_l2_in_3__A1 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_14.mux_l1_in_0__A0 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__52__A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_1.mux_l3_in_0_/S mux_right_ipin_1.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_4.mux_l2_in_0__A1 mux_right_ipin_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__47__A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_2.mux_l4_in_0_ mux_right_ipin_2.mux_l3_in_1_/X mux_right_ipin_2.mux_l3_in_0_/X
+ mux_right_ipin_2.mux_l4_in_0_/S mux_right_ipin_2.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_12.mux_l1_in_2__A0 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_9.mux_l2_in_3__A0 _20_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_1.mux_l2_in_1__S mux_right_ipin_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_11.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_2__A1 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_ipin_0.mux_l2_in_0_ mux_left_ipin_0.mux_l1_in_1_/X mux_left_ipin_0.mux_l1_in_0_/X
+ mux_left_ipin_0.mux_l2_in_0_/S mux_left_ipin_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_7.mux_l1_in_2__S mux_right_ipin_7.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_7.mux_l2_in_3_ _18_/HI chany_top_in[18] mux_right_ipin_7.mux_l2_in_2_/S
+ mux_right_ipin_7.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_53_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_1_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l2_in_1__A0 chany_bottom_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_2.mux_l3_in_1_ mux_right_ipin_2.mux_l2_in_3_/X mux_right_ipin_2.mux_l2_in_2_/X
+ mux_right_ipin_2.mux_l3_in_1_/S mux_right_ipin_2.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__60__A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_2.mux_l3_in_1__A1 mux_right_ipin_2.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_0.mux_l3_in_1__S mux_right_ipin_0.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__55__A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_10.mux_l2_in_3__A0 _24_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_ipin_0.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_left_ipin_0.mux_l1_in_2_/S
+ mux_left_ipin_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l3_in_0__A0 mux_right_ipin_12.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_6.mux_l2_in_2__S mux_right_ipin_6.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_2.mux_l2_in_2_ chany_bottom_in[15] chany_top_in[7] mux_right_ipin_2.mux_l2_in_3_/S
+ mux_right_ipin_2.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_4.mux_l3_in_0_/S mux_right_ipin_4.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_7.mux_l4_in_0_ mux_right_ipin_7.mux_l3_in_1_/X mux_right_ipin_7.mux_l3_in_0_/X
+ mux_right_ipin_7.mux_l4_in_0_/S mux_right_ipin_7.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_2.mux_l4_in_0__A1 mux_right_ipin_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_14.mux_l1_in_0__A1 chany_bottom_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_14.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_7.mux_l3_in_1_ mux_right_ipin_7.mux_l2_in_3_/X mux_right_ipin_7.mux_l2_in_2_/X
+ mux_right_ipin_7.mux_l3_in_1_/S mux_right_ipin_7.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_1.mux_l2_in_0_/S mux_right_ipin_1.mux_l3_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__63__A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l1_in_2__A1 chany_bottom_in[7] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_9.mux_l4_in_0__S mux_right_ipin_9.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_prog_clk clkbuf_1_1_0_prog_clk/X clkbuf_3_7_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_9.mux_l2_in_3__A1 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_8.mux_l1_in_0__A0 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__58__A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_7.mux_l2_in_2_ chany_bottom_in[18] chany_top_in[12] mux_right_ipin_7.mux_l2_in_2_/S
+ mux_right_ipin_7.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_12.mux_l2_in_1__A1 mux_right_ipin_12.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_2.mux_l3_in_0_ mux_right_ipin_2.mux_l2_in_1_/X mux_right_ipin_2.mux_l2_in_0_/X
+ mux_right_ipin_2.mux_l3_in_1_/S mux_right_ipin_2.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_7.mux_l3_in_1_/S mux_right_ipin_7.mux_l4_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_13.mux_l2_in_2__S mux_right_ipin_13.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_ipin_0.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_left_ipin_0.mux_l1_in_2_/S
+ mux_left_ipin_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_10.mux_l2_in_3__A1 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__71__A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_12.mux_l3_in_0__A1 mux_right_ipin_12.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_2.mux_l2_in_1_ chany_bottom_in[7] chany_top_in[3] mux_right_ipin_2.mux_l2_in_3_/S
+ mux_right_ipin_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_6.mux_l2_in_1__A0 chany_bottom_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_36_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_13.mux_l4_in_0_/X left_grid_pin_29_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_4.mux_l2_in_0_/S mux_right_ipin_4.mux_l3_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__66__A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_5.mux_l4_in_0_/X left_grid_pin_21_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_ipin_4.mux_l2_in_3__A0 _32_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_prog_clk clkbuf_3_5_0_prog_clk/A clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_11.mux_l2_in_3_ _25_/HI chany_top_in[16] mux_right_ipin_11.mux_l2_in_0_/S
+ mux_right_ipin_11.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_53_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_6.mux_l3_in_0__A0 mux_right_ipin_6.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_69_ chany_bottom_in[4] chany_top_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_ipin_7.mux_l3_in_0_ mux_right_ipin_7.mux_l2_in_1_/X mux_right_ipin_7.mux_l2_in_0_/X
+ mux_right_ipin_7.mux_l3_in_1_/S mux_right_ipin_7.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_1.mux_l1_in_0_/S mux_right_ipin_1.mux_l2_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_8.mux_l1_in_0__A1 chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__74__A ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_7.mux_l2_in_1_ chany_bottom_in[12] mux_right_ipin_7.mux_l1_in_2_/X
+ mux_right_ipin_7.mux_l2_in_2_/S mux_right_ipin_7.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_8.mux_l1_in_0__S mux_right_ipin_8.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_12.mux_l3_in_0_/S mux_right_ipin_12.mux_l4_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_11.mux_l4_in_0_ mux_right_ipin_11.mux_l3_in_1_/X mux_right_ipin_11.mux_l3_in_0_/X
+ mux_right_ipin_11.mux_l4_in_0_/S mux_right_ipin_11.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__69__A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_7.mux_l2_in_2_/S mux_right_ipin_7.mux_l3_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_9.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_3.mux_l1_in_2__S mux_right_ipin_3.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_7.mux_l1_in_2_ chany_top_in[8] chany_bottom_in[8] mux_right_ipin_7.mux_l1_in_2_/S
+ mux_right_ipin_7.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_ipin_0.mux_l1_in_2__S mux_left_ipin_0.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
+ mux_right_ipin_15.mux_l4_in_0_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_0__S mux_right_ipin_7.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_11.mux_l3_in_1_ mux_right_ipin_11.mux_l2_in_3_/X mux_right_ipin_11.mux_l2_in_2_/X
+ mux_right_ipin_11.mux_l3_in_0_/S mux_right_ipin_11.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_2.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_2.mux_l1_in_0_/X
+ mux_right_ipin_2.mux_l2_in_3_/S mux_right_ipin_2.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_6.mux_l2_in_1__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_4.mux_l1_in_1_/S mux_right_ipin_4.mux_l2_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_left_ipin_0.mux_l4_in_0_/X right_grid_pin_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_2.mux_l2_in_2__S mux_right_ipin_2.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_4.mux_l2_in_3__A1 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__77__A gfpga_pad_EMBEDDED_IO_SOC_IN VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_11.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[12] mux_right_ipin_11.mux_l2_in_0_/S
+ mux_right_ipin_11.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_2_0_prog_clk_A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_6.mux_l3_in_0__A1 mux_right_ipin_6.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0__A0 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_68_ chany_bottom_in[5] chany_top_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_6.mux_l3_in_0__S mux_right_ipin_6.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_14.mux_l2_in_2__A0 chany_bottom_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_15.mux_l3_in_0_/S mux_right_ipin_15.mux_l4_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_0.mux_l4_in_0_/S mux_right_ipin_1.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_ipin_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_15.mux_l1_in_0__S mux_right_ipin_15.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_ipin_14.mux_l3_in_1__A0 mux_right_ipin_14.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_7.mux_l2_in_0_ mux_right_ipin_7.mux_l1_in_1_/X mux_right_ipin_7.mux_l1_in_0_/X
+ mux_right_ipin_7.mux_l2_in_2_/S mux_right_ipin_7.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_7.mux_l2_in_3__S mux_right_ipin_7.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_12.mux_l2_in_0_/S mux_right_ipin_12.mux_l3_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_5.mux_l4_in_0__S mux_right_ipin_5.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_7.mux_l1_in_2_/S mux_right_ipin_7.mux_l2_in_2_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_1.mux_l2_in_1__A0 chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_14.mux_l2_in_0__S mux_right_ipin_14.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_2__A0 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_14.mux_l4_in_0__A0 mux_right_ipin_14.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_prog_clk_A clkbuf_3_7_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_7.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_7.mux_l1_in_2_/S
+ mux_right_ipin_7.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_0_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_ipin_11.mux_l3_in_0_ mux_right_ipin_11.mux_l2_in_1_/X mux_right_ipin_11.mux_l2_in_0_/X
+ mux_right_ipin_11.mux_l3_in_0_/S mux_right_ipin_11.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_1.mux_l3_in_0__A0 mux_right_ipin_1.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_3.mux_l4_in_0_/S mux_right_ipin_4.mux_l1_in_1_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_1.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_ipin_0.mux_l2_in_1__A0 chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_13.mux_l3_in_0__S mux_right_ipin_13.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_11.mux_l2_in_1_ chany_bottom_in[12] mux_right_ipin_11.mux_l1_in_2_/X
+ mux_right_ipin_11.mux_l2_in_0_/S mux_right_ipin_11.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_2.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_2.mux_l1_in_0_/S
+ mux_right_ipin_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_3.mux_l1_in_0__A1 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_67_ chany_bottom_in[6] chany_top_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_14.mux_l2_in_2__A1 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_15.mux_l2_in_0_/S mux_right_ipin_15.mux_l3_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_13.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_ipin_0.mux_l3_in_0__A0 mux_left_ipin_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_14.mux_l2_in_3__S mux_right_ipin_14.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_11.mux_l1_in_2_ chany_top_in[6] chany_bottom_in[6] mux_right_ipin_11.mux_l1_in_0_/S
+ mux_right_ipin_11.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_12.mux_l4_in_0__S mux_right_ipin_12.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_6.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_11.mux_l1_in_1__A0 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_14.mux_l3_in_1__A1 mux_right_ipin_14.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_12.mux_l1_in_0_/S mux_right_ipin_12.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_8.mux_l2_in_2__A0 chany_bottom_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_prog_clk clkbuf_1_1_0_prog_clk/X clkbuf_3_5_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_ipin_6.mux_l4_in_0_/S mux_right_ipin_7.mux_l1_in_2_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_45_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_1__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_4.mux_l1_in_0__S mux_right_ipin_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_11.mux_l2_in_0__A0 mux_right_ipin_11.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_14.mux_l4_in_0__A1 mux_right_ipin_14.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_2__A1 chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_7.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_7.mux_l1_in_2_/S
+ mux_right_ipin_7.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_8.mux_l3_in_1__A0 mux_right_ipin_8.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

