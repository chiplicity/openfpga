magic
tech sky130A
magscale 1 2
timestamp 1606426458
<< locali >>
rect 9815 17901 10057 17935
rect 11195 17765 11529 17799
rect 9505 13175 9539 13277
rect 12265 10455 12299 10693
rect 12265 9503 12299 9605
rect 4169 9027 4203 9129
rect 949 2023 983 8925
<< viali >>
rect 9781 17901 9815 17935
rect 10057 17901 10091 17935
rect 11161 17765 11195 17799
rect 11529 17765 11563 17799
rect 12817 17289 12851 17323
rect 13553 17289 13587 17323
rect 10701 17221 10735 17255
rect 1777 17153 1811 17187
rect 2605 17153 2639 17187
rect 4261 17153 4295 17187
rect 6285 17153 6319 17187
rect 7481 17153 7515 17187
rect 8677 17153 8711 17187
rect 1501 17085 1535 17119
rect 2421 17085 2455 17119
rect 4077 17085 4111 17119
rect 8493 17085 8527 17119
rect 9505 17085 9539 17119
rect 9781 17085 9815 17119
rect 10517 17085 10551 17119
rect 11253 17085 11287 17119
rect 12633 17085 12667 17119
rect 13369 17085 13403 17119
rect 7389 17017 7423 17051
rect 3249 16949 3283 16983
rect 3341 16949 3375 16983
rect 4905 16949 4939 16983
rect 4997 16949 5031 16983
rect 5641 16949 5675 16983
rect 6009 16949 6043 16983
rect 6101 16949 6135 16983
rect 6929 16949 6963 16983
rect 7297 16949 7331 16983
rect 8125 16949 8159 16983
rect 8585 16949 8619 16983
rect 9321 16949 9355 16983
rect 9965 16949 9999 16983
rect 11437 16949 11471 16983
rect 2513 16745 2547 16779
rect 3709 16745 3743 16779
rect 4997 16745 5031 16779
rect 5457 16745 5491 16779
rect 6285 16745 6319 16779
rect 6653 16745 6687 16779
rect 7481 16745 7515 16779
rect 7849 16745 7883 16779
rect 7941 16745 7975 16779
rect 9873 16745 9907 16779
rect 10609 16745 10643 16779
rect 13553 16745 13587 16779
rect 14289 16745 14323 16779
rect 1685 16677 1719 16711
rect 3065 16677 3099 16711
rect 6745 16677 6779 16711
rect 1409 16609 1443 16643
rect 2697 16609 2731 16643
rect 2789 16609 2823 16643
rect 3893 16609 3927 16643
rect 4077 16609 4111 16643
rect 4353 16609 4387 16643
rect 5365 16609 5399 16643
rect 8677 16609 8711 16643
rect 8953 16609 8987 16643
rect 9689 16609 9723 16643
rect 10425 16609 10459 16643
rect 11161 16609 11195 16643
rect 11897 16609 11931 16643
rect 12633 16609 12667 16643
rect 13369 16609 13403 16643
rect 14105 16609 14139 16643
rect 5549 16541 5583 16575
rect 6837 16541 6871 16575
rect 8033 16541 8067 16575
rect 11345 16473 11379 16507
rect 12081 16473 12115 16507
rect 12817 16473 12851 16507
rect 5549 16201 5583 16235
rect 8033 16201 8067 16235
rect 10609 16201 10643 16235
rect 13369 16201 13403 16235
rect 12633 16133 12667 16167
rect 1685 16065 1719 16099
rect 2605 16065 2639 16099
rect 4997 16065 5031 16099
rect 6009 16065 6043 16099
rect 6101 16065 6135 16099
rect 7389 16065 7423 16099
rect 8585 16065 8619 16099
rect 9781 16065 9815 16099
rect 1501 15997 1535 16031
rect 2421 15997 2455 16031
rect 3341 15997 3375 16031
rect 4813 15997 4847 16031
rect 5917 15997 5951 16031
rect 7297 15997 7331 16031
rect 8493 15997 8527 16031
rect 9597 15997 9631 16031
rect 9689 15997 9723 16031
rect 10425 15997 10459 16031
rect 11161 15997 11195 16031
rect 12449 15997 12483 16031
rect 13185 15997 13219 16031
rect 3617 15929 3651 15963
rect 7205 15929 7239 15963
rect 8401 15929 8435 15963
rect 4353 15861 4387 15895
rect 4721 15861 4755 15895
rect 6837 15861 6871 15895
rect 9229 15861 9263 15895
rect 11345 15861 11379 15895
rect 3433 15657 3467 15691
rect 7205 15657 7239 15691
rect 8125 15657 8159 15691
rect 9045 15657 9079 15691
rect 11069 15657 11103 15691
rect 11805 15657 11839 15691
rect 12541 15657 12575 15691
rect 4997 15589 5031 15623
rect 1409 15521 1443 15555
rect 2329 15521 2363 15555
rect 3249 15521 3283 15555
rect 5825 15521 5859 15555
rect 6092 15521 6126 15555
rect 8033 15521 8067 15555
rect 8861 15521 8895 15555
rect 10057 15521 10091 15555
rect 10149 15521 10183 15555
rect 10885 15521 10919 15555
rect 11621 15521 11655 15555
rect 12357 15521 12391 15555
rect 1685 15453 1719 15487
rect 2513 15453 2547 15487
rect 5089 15453 5123 15487
rect 5273 15453 5307 15487
rect 8217 15453 8251 15487
rect 10241 15453 10275 15487
rect 13093 15453 13127 15487
rect 13737 15453 13771 15487
rect 4629 15317 4663 15351
rect 7665 15317 7699 15351
rect 9689 15317 9723 15351
rect 3709 15113 3743 15147
rect 8677 15113 8711 15147
rect 11069 15045 11103 15079
rect 2053 14977 2087 15011
rect 4169 14977 4203 15011
rect 4353 14977 4387 15011
rect 6837 14977 6871 15011
rect 9229 14977 9263 15011
rect 10425 14977 10459 15011
rect 11529 14977 11563 15011
rect 11621 14977 11655 15011
rect 12449 14977 12483 15011
rect 1777 14909 1811 14943
rect 2697 14909 2731 14943
rect 4905 14909 4939 14943
rect 9045 14909 9079 14943
rect 2973 14841 3007 14875
rect 4077 14841 4111 14875
rect 5172 14841 5206 14875
rect 7082 14841 7116 14875
rect 10333 14841 10367 14875
rect 6285 14773 6319 14807
rect 8217 14773 8251 14807
rect 9137 14773 9171 14807
rect 9873 14773 9907 14807
rect 10241 14773 10275 14807
rect 11437 14773 11471 14807
rect 13093 14773 13127 14807
rect 13737 14773 13771 14807
rect 14381 14773 14415 14807
rect 2789 14569 2823 14603
rect 4445 14569 4479 14603
rect 4905 14569 4939 14603
rect 7021 14569 7055 14603
rect 9689 14569 9723 14603
rect 14105 14569 14139 14603
rect 2145 14501 2179 14535
rect 3249 14501 3283 14535
rect 5886 14501 5920 14535
rect 11345 14501 11379 14535
rect 1869 14433 1903 14467
rect 3157 14433 3191 14467
rect 4813 14433 4847 14467
rect 7748 14433 7782 14467
rect 9505 14433 9539 14467
rect 10057 14433 10091 14467
rect 11253 14433 11287 14467
rect 12081 14433 12115 14467
rect 13369 14433 13403 14467
rect 3433 14365 3467 14399
rect 5089 14365 5123 14399
rect 5641 14365 5675 14399
rect 7481 14365 7515 14399
rect 10149 14365 10183 14399
rect 10241 14365 10275 14399
rect 11437 14365 11471 14399
rect 12265 14365 12299 14399
rect 8861 14297 8895 14331
rect 10885 14297 10919 14331
rect 9321 14229 9355 14263
rect 13553 14229 13587 14263
rect 3709 14025 3743 14059
rect 10517 14025 10551 14059
rect 2513 13957 2547 13991
rect 6285 13957 6319 13991
rect 8217 13957 8251 13991
rect 12449 13957 12483 13991
rect 14013 13957 14047 13991
rect 1777 13889 1811 13923
rect 3157 13889 3191 13923
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 11069 13889 11103 13923
rect 13001 13889 13035 13923
rect 1593 13821 1627 13855
rect 2973 13821 3007 13855
rect 4905 13821 4939 13855
rect 6837 13821 6871 13855
rect 7104 13821 7138 13855
rect 8677 13821 8711 13855
rect 8933 13821 8967 13855
rect 10977 13821 11011 13855
rect 13829 13821 13863 13855
rect 5172 13753 5206 13787
rect 10885 13753 10919 13787
rect 11713 13753 11747 13787
rect 12817 13753 12851 13787
rect 14565 13753 14599 13787
rect 2881 13685 2915 13719
rect 4077 13685 4111 13719
rect 10057 13685 10091 13719
rect 12909 13685 12943 13719
rect 1961 13481 1995 13515
rect 5733 13481 5767 13515
rect 8033 13481 8067 13515
rect 11529 13481 11563 13515
rect 11897 13481 11931 13515
rect 13185 13481 13219 13515
rect 3157 13413 3191 13447
rect 6438 13413 6472 13447
rect 11989 13413 12023 13447
rect 4353 13345 4387 13379
rect 4620 13345 4654 13379
rect 6193 13345 6227 13379
rect 8401 13345 8435 13379
rect 9413 13345 9447 13379
rect 9956 13345 9990 13379
rect 13093 13345 13127 13379
rect 13921 13345 13955 13379
rect 2053 13277 2087 13311
rect 2237 13277 2271 13311
rect 3249 13277 3283 13311
rect 3433 13277 3467 13311
rect 8493 13277 8527 13311
rect 8677 13277 8711 13311
rect 9505 13277 9539 13311
rect 9689 13277 9723 13311
rect 12173 13277 12207 13311
rect 13369 13277 13403 13311
rect 14105 13277 14139 13311
rect 1593 13209 1627 13243
rect 11069 13209 11103 13243
rect 12725 13209 12759 13243
rect 2789 13141 2823 13175
rect 7573 13141 7607 13175
rect 9229 13141 9263 13175
rect 9505 13141 9539 13175
rect 6285 12937 6319 12971
rect 8217 12937 8251 12971
rect 13645 12937 13679 12971
rect 1869 12869 1903 12903
rect 4445 12869 4479 12903
rect 10517 12869 10551 12903
rect 12449 12869 12483 12903
rect 2513 12801 2547 12835
rect 8677 12801 8711 12835
rect 11069 12801 11103 12835
rect 13001 12801 13035 12835
rect 2237 12733 2271 12767
rect 3065 12733 3099 12767
rect 4905 12733 4939 12767
rect 5172 12733 5206 12767
rect 6837 12733 6871 12767
rect 7104 12733 7138 12767
rect 10885 12733 10919 12767
rect 13829 12733 13863 12767
rect 13921 12733 13955 12767
rect 14841 12733 14875 12767
rect 3332 12665 3366 12699
rect 8922 12665 8956 12699
rect 10977 12665 11011 12699
rect 14197 12665 14231 12699
rect 2329 12597 2363 12631
rect 10057 12597 10091 12631
rect 11713 12597 11747 12631
rect 12817 12597 12851 12631
rect 12909 12597 12943 12631
rect 15025 12597 15059 12631
rect 2789 12393 2823 12427
rect 3157 12393 3191 12427
rect 3249 12393 3283 12427
rect 6929 12393 6963 12427
rect 9229 12393 9263 12427
rect 11253 12393 11287 12427
rect 12541 12393 12575 12427
rect 2053 12325 2087 12359
rect 4721 12325 4755 12359
rect 5794 12325 5828 12359
rect 7656 12325 7690 12359
rect 10057 12325 10091 12359
rect 11345 12325 11379 12359
rect 12449 12325 12483 12359
rect 1961 12257 1995 12291
rect 5549 12257 5583 12291
rect 9413 12257 9447 12291
rect 13461 12257 13495 12291
rect 13553 12257 13587 12291
rect 14473 12257 14507 12291
rect 2237 12189 2271 12223
rect 3433 12189 3467 12223
rect 4813 12189 4847 12223
rect 4905 12189 4939 12223
rect 7389 12189 7423 12223
rect 10149 12189 10183 12223
rect 10333 12189 10367 12223
rect 11437 12189 11471 12223
rect 12633 12189 12667 12223
rect 13829 12189 13863 12223
rect 13277 12121 13311 12155
rect 1593 12053 1627 12087
rect 4353 12053 4387 12087
rect 8769 12053 8803 12087
rect 9689 12053 9723 12087
rect 10885 12053 10919 12087
rect 12081 12053 12115 12087
rect 14657 12053 14691 12087
rect 2513 11849 2547 11883
rect 3709 11849 3743 11883
rect 10425 11849 10459 11883
rect 12449 11781 12483 11815
rect 3157 11713 3191 11747
rect 4261 11713 4295 11747
rect 7389 11713 7423 11747
rect 9781 11713 9815 11747
rect 10885 11713 10919 11747
rect 11069 11713 11103 11747
rect 13001 11713 13035 11747
rect 13921 11713 13955 11747
rect 1593 11645 1627 11679
rect 2881 11645 2915 11679
rect 4077 11645 4111 11679
rect 4905 11645 4939 11679
rect 7656 11645 7690 11679
rect 10793 11645 10827 11679
rect 11621 11645 11655 11679
rect 13645 11645 13679 11679
rect 14565 11645 14599 11679
rect 1869 11577 1903 11611
rect 2973 11577 3007 11611
rect 5172 11577 5206 11611
rect 9597 11577 9631 11611
rect 12817 11577 12851 11611
rect 14841 11577 14875 11611
rect 4169 11509 4203 11543
rect 6285 11509 6319 11543
rect 8769 11509 8803 11543
rect 9229 11509 9263 11543
rect 9689 11509 9723 11543
rect 11805 11509 11839 11543
rect 12909 11509 12943 11543
rect 1593 11305 1627 11339
rect 3157 11305 3191 11339
rect 4629 11305 4663 11339
rect 10149 11305 10183 11339
rect 11345 11305 11379 11339
rect 13277 11305 13311 11339
rect 4997 11237 5031 11271
rect 10057 11237 10091 11271
rect 12541 11237 12575 11271
rect 1961 11169 1995 11203
rect 2053 11169 2087 11203
rect 5089 11169 5123 11203
rect 5825 11169 5859 11203
rect 6092 11169 6126 11203
rect 7932 11169 7966 11203
rect 11253 11169 11287 11203
rect 12449 11169 12483 11203
rect 13645 11169 13679 11203
rect 14473 11169 14507 11203
rect 2145 11101 2179 11135
rect 3249 11101 3283 11135
rect 3433 11101 3467 11135
rect 5273 11101 5307 11135
rect 7665 11101 7699 11135
rect 10333 11101 10367 11135
rect 11437 11101 11471 11135
rect 12633 11101 12667 11135
rect 13737 11101 13771 11135
rect 13829 11101 13863 11135
rect 2789 11033 2823 11067
rect 9689 11033 9723 11067
rect 10885 11033 10919 11067
rect 12081 11033 12115 11067
rect 14657 11033 14691 11067
rect 7205 10965 7239 10999
rect 9045 10965 9079 10999
rect 3709 10761 3743 10795
rect 6837 10761 6871 10795
rect 8033 10761 8067 10795
rect 10333 10761 10367 10795
rect 11713 10761 11747 10795
rect 13645 10761 13679 10795
rect 2513 10693 2547 10727
rect 12265 10693 12299 10727
rect 2973 10625 3007 10659
rect 3157 10625 3191 10659
rect 4353 10625 4387 10659
rect 4905 10625 4939 10659
rect 7297 10625 7331 10659
rect 7481 10625 7515 10659
rect 10885 10625 10919 10659
rect 1593 10557 1627 10591
rect 4077 10557 4111 10591
rect 4169 10557 4203 10591
rect 8217 10557 8251 10591
rect 8493 10557 8527 10591
rect 10701 10557 10735 10591
rect 11529 10557 11563 10591
rect 1869 10489 1903 10523
rect 5150 10489 5184 10523
rect 7205 10489 7239 10523
rect 8760 10489 8794 10523
rect 12909 10625 12943 10659
rect 13001 10625 13035 10659
rect 14197 10625 14231 10659
rect 12817 10557 12851 10591
rect 14013 10557 14047 10591
rect 14841 10557 14875 10591
rect 14105 10489 14139 10523
rect 2881 10421 2915 10455
rect 6285 10421 6319 10455
rect 9873 10421 9907 10455
rect 10793 10421 10827 10455
rect 12265 10421 12299 10455
rect 12449 10421 12483 10455
rect 15025 10421 15059 10455
rect 1961 10217 1995 10251
rect 2789 10217 2823 10251
rect 4261 10217 4295 10251
rect 4721 10217 4755 10251
rect 10885 10217 10919 10251
rect 11345 10217 11379 10251
rect 12541 10217 12575 10251
rect 13277 10217 13311 10251
rect 4629 10149 4663 10183
rect 7542 10149 7576 10183
rect 10057 10149 10091 10183
rect 11253 10149 11287 10183
rect 12449 10149 12483 10183
rect 2053 10081 2087 10115
rect 3157 10081 3191 10115
rect 3249 10081 3283 10115
rect 5724 10081 5758 10115
rect 7297 10081 7331 10115
rect 9321 10081 9355 10115
rect 10149 10081 10183 10115
rect 13645 10081 13679 10115
rect 13737 10081 13771 10115
rect 14473 10081 14507 10115
rect 2237 10013 2271 10047
rect 3433 10013 3467 10047
rect 4813 10013 4847 10047
rect 5457 10013 5491 10047
rect 10333 10013 10367 10047
rect 11529 10013 11563 10047
rect 12725 10013 12759 10047
rect 13829 10013 13863 10047
rect 8677 9945 8711 9979
rect 14657 9945 14691 9979
rect 1593 9877 1627 9911
rect 6837 9877 6871 9911
rect 9137 9877 9171 9911
rect 9689 9877 9723 9911
rect 12081 9877 12115 9911
rect 5181 9673 5215 9707
rect 2145 9605 2179 9639
rect 2973 9605 3007 9639
rect 8677 9605 8711 9639
rect 9873 9605 9907 9639
rect 12265 9605 12299 9639
rect 12449 9605 12483 9639
rect 2605 9537 2639 9571
rect 2789 9537 2823 9571
rect 3617 9537 3651 9571
rect 6837 9537 6871 9571
rect 9229 9537 9263 9571
rect 10425 9537 10459 9571
rect 11529 9537 11563 9571
rect 11713 9537 11747 9571
rect 13001 9537 13035 9571
rect 14105 9537 14139 9571
rect 14197 9537 14231 9571
rect 1593 9469 1627 9503
rect 1869 9469 1903 9503
rect 3801 9469 3835 9503
rect 5273 9469 5307 9503
rect 9137 9469 9171 9503
rect 10241 9469 10275 9503
rect 11437 9469 11471 9503
rect 12265 9469 12299 9503
rect 14841 9469 14875 9503
rect 2513 9401 2547 9435
rect 4068 9401 4102 9435
rect 5540 9401 5574 9435
rect 7082 9401 7116 9435
rect 12817 9401 12851 9435
rect 3341 9333 3375 9367
rect 3433 9333 3467 9367
rect 6653 9333 6687 9367
rect 8217 9333 8251 9367
rect 9045 9333 9079 9367
rect 10333 9333 10367 9367
rect 11069 9333 11103 9367
rect 12909 9333 12943 9367
rect 13645 9333 13679 9367
rect 14013 9333 14047 9367
rect 15025 9333 15059 9367
rect 2789 9129 2823 9163
rect 4169 9129 4203 9163
rect 4261 9129 4295 9163
rect 7757 9129 7791 9163
rect 10057 9129 10091 9163
rect 11345 9129 11379 9163
rect 12081 9129 12115 9163
rect 12449 9129 12483 9163
rect 13277 9129 13311 9163
rect 13737 9129 13771 9163
rect 4629 9061 4663 9095
rect 10149 9061 10183 9095
rect 1961 8993 1995 9027
rect 3157 8993 3191 9027
rect 4169 8993 4203 9027
rect 4721 8993 4755 9027
rect 5917 8993 5951 9027
rect 7665 8993 7699 9027
rect 8125 8993 8159 9027
rect 8217 8993 8251 9027
rect 8585 8993 8619 9027
rect 11253 8993 11287 9027
rect 12541 8993 12575 9027
rect 13645 8993 13679 9027
rect 14473 8993 14507 9027
rect 949 8925 983 8959
rect 2053 8925 2087 8959
rect 2237 8925 2271 8959
rect 3249 8925 3283 8959
rect 3433 8925 3467 8959
rect 4905 8925 4939 8959
rect 8401 8925 8435 8959
rect 8769 8925 8803 8959
rect 10241 8925 10275 8959
rect 11437 8925 11471 8959
rect 12633 8925 12667 8959
rect 13829 8925 13863 8959
rect 10885 8857 10919 8891
rect 1593 8789 1627 8823
rect 9689 8789 9723 8823
rect 14657 8789 14691 8823
rect 11069 8585 11103 8619
rect 12449 8585 12483 8619
rect 13645 8585 13679 8619
rect 3709 8517 3743 8551
rect 6285 8517 6319 8551
rect 2973 8449 3007 8483
rect 3157 8449 3191 8483
rect 4353 8449 4387 8483
rect 9229 8449 9263 8483
rect 10425 8449 10459 8483
rect 11713 8449 11747 8483
rect 13001 8449 13035 8483
rect 14289 8449 14323 8483
rect 1593 8381 1627 8415
rect 2881 8381 2915 8415
rect 4905 8381 4939 8415
rect 5172 8381 5206 8415
rect 6837 8381 6871 8415
rect 11529 8381 11563 8415
rect 14105 8381 14139 8415
rect 14841 8381 14875 8415
rect 1869 8313 1903 8347
rect 4077 8313 4111 8347
rect 4169 8313 4203 8347
rect 7082 8313 7116 8347
rect 10333 8313 10367 8347
rect 12909 8313 12943 8347
rect 14013 8313 14047 8347
rect 2513 8245 2547 8279
rect 8217 8245 8251 8279
rect 8677 8245 8711 8279
rect 9045 8245 9079 8279
rect 9137 8245 9171 8279
rect 9873 8245 9907 8279
rect 10241 8245 10275 8279
rect 11437 8245 11471 8279
rect 12817 8245 12851 8279
rect 15025 8245 15059 8279
rect 1961 8041 1995 8075
rect 7297 8041 7331 8075
rect 9137 8041 9171 8075
rect 9689 8041 9723 8075
rect 10149 8041 10183 8075
rect 10885 8041 10919 8075
rect 12081 8041 12115 8075
rect 12449 8041 12483 8075
rect 3157 7973 3191 8007
rect 11253 7973 11287 8007
rect 4077 7905 4111 7939
rect 4344 7905 4378 7939
rect 6173 7905 6207 7939
rect 8024 7905 8058 7939
rect 10057 7905 10091 7939
rect 13645 7905 13679 7939
rect 14473 7905 14507 7939
rect 2053 7837 2087 7871
rect 2237 7837 2271 7871
rect 3249 7837 3283 7871
rect 3433 7837 3467 7871
rect 5917 7837 5951 7871
rect 7757 7837 7791 7871
rect 10241 7837 10275 7871
rect 11345 7837 11379 7871
rect 11529 7837 11563 7871
rect 12541 7837 12575 7871
rect 12725 7837 12759 7871
rect 13737 7837 13771 7871
rect 13921 7837 13955 7871
rect 13277 7769 13311 7803
rect 1593 7701 1627 7735
rect 2789 7701 2823 7735
rect 5457 7701 5491 7735
rect 14657 7701 14691 7735
rect 1869 7497 1903 7531
rect 4445 7429 4479 7463
rect 8217 7429 8251 7463
rect 10517 7429 10551 7463
rect 2329 7361 2363 7395
rect 2513 7361 2547 7395
rect 10977 7361 11011 7395
rect 11069 7361 11103 7395
rect 12909 7361 12943 7395
rect 13093 7361 13127 7395
rect 14197 7361 14231 7395
rect 3065 7293 3099 7327
rect 4905 7293 4939 7327
rect 6837 7293 6871 7327
rect 7093 7293 7127 7327
rect 8677 7293 8711 7327
rect 8933 7293 8967 7327
rect 10885 7293 10919 7327
rect 11713 7293 11747 7327
rect 14841 7293 14875 7327
rect 3332 7225 3366 7259
rect 5172 7225 5206 7259
rect 14105 7225 14139 7259
rect 2237 7157 2271 7191
rect 6285 7157 6319 7191
rect 10057 7157 10091 7191
rect 12449 7157 12483 7191
rect 12817 7157 12851 7191
rect 13645 7157 13679 7191
rect 14013 7157 14047 7191
rect 15025 7157 15059 7191
rect 7113 6953 7147 6987
rect 8953 6953 8987 6987
rect 10057 6953 10091 6987
rect 12081 6953 12115 6987
rect 13277 6953 13311 6987
rect 11253 6885 11287 6919
rect 12449 6885 12483 6919
rect 13645 6885 13679 6919
rect 1409 6817 1443 6851
rect 2412 6817 2446 6851
rect 4261 6817 4295 6851
rect 5089 6817 5123 6851
rect 6000 6817 6034 6851
rect 7573 6817 7607 6851
rect 7829 6817 7863 6851
rect 14473 6817 14507 6851
rect 2145 6749 2179 6783
rect 5733 6749 5767 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 11345 6749 11379 6783
rect 11437 6749 11471 6783
rect 12541 6749 12575 6783
rect 12633 6749 12667 6783
rect 13737 6749 13771 6783
rect 13921 6749 13955 6783
rect 3525 6681 3559 6715
rect 1593 6613 1627 6647
rect 9689 6613 9723 6647
rect 10885 6613 10919 6647
rect 14657 6613 14691 6647
rect 1869 6409 1903 6443
rect 4445 6409 4479 6443
rect 15025 6409 15059 6443
rect 6285 6341 6319 6375
rect 8217 6341 8251 6375
rect 13645 6341 13679 6375
rect 2513 6273 2547 6307
rect 4905 6273 4939 6307
rect 6837 6273 6871 6307
rect 10977 6273 11011 6307
rect 11161 6273 11195 6307
rect 13001 6273 13035 6307
rect 14105 6273 14139 6307
rect 14289 6273 14323 6307
rect 3065 6205 3099 6239
rect 8677 6205 8711 6239
rect 10885 6205 10919 6239
rect 14841 6205 14875 6239
rect 2237 6137 2271 6171
rect 3332 6137 3366 6171
rect 5172 6137 5206 6171
rect 7104 6137 7138 6171
rect 8922 6137 8956 6171
rect 12817 6137 12851 6171
rect 2329 6069 2363 6103
rect 10057 6069 10091 6103
rect 10517 6069 10551 6103
rect 11713 6069 11747 6103
rect 12449 6069 12483 6103
rect 12909 6069 12943 6103
rect 14013 6069 14047 6103
rect 3525 5865 3559 5899
rect 4629 5865 4663 5899
rect 9137 5865 9171 5899
rect 11069 5865 11103 5899
rect 12725 5865 12759 5899
rect 13093 5865 13127 5899
rect 13185 5865 13219 5899
rect 4721 5797 4755 5831
rect 1409 5729 1443 5763
rect 2145 5729 2179 5763
rect 2412 5729 2446 5763
rect 5457 5729 5491 5763
rect 5724 5729 5758 5763
rect 7564 5729 7598 5763
rect 9321 5729 9355 5763
rect 9945 5729 9979 5763
rect 11897 5729 11931 5763
rect 14289 5729 14323 5763
rect 4905 5661 4939 5695
rect 7297 5661 7331 5695
rect 9689 5661 9723 5695
rect 11989 5661 12023 5695
rect 12081 5661 12115 5695
rect 13369 5661 13403 5695
rect 14381 5661 14415 5695
rect 14473 5661 14507 5695
rect 1593 5525 1627 5559
rect 4261 5525 4295 5559
rect 6837 5525 6871 5559
rect 8677 5525 8711 5559
rect 11529 5525 11563 5559
rect 13921 5525 13955 5559
rect 8217 5321 8251 5355
rect 12449 5321 12483 5355
rect 13645 5321 13679 5355
rect 4445 5253 4479 5287
rect 10057 5253 10091 5287
rect 15025 5253 15059 5287
rect 2513 5185 2547 5219
rect 10977 5185 11011 5219
rect 11069 5185 11103 5219
rect 11713 5185 11747 5219
rect 13001 5185 13035 5219
rect 14289 5185 14323 5219
rect 2237 5117 2271 5151
rect 3065 5117 3099 5151
rect 3332 5117 3366 5151
rect 4905 5117 4939 5151
rect 5172 5117 5206 5151
rect 6837 5117 6871 5151
rect 8677 5117 8711 5151
rect 14841 5117 14875 5151
rect 7104 5049 7138 5083
rect 8944 5049 8978 5083
rect 13461 5049 13495 5083
rect 14013 5049 14047 5083
rect 14105 5049 14139 5083
rect 1869 4981 1903 5015
rect 2329 4981 2363 5015
rect 6285 4981 6319 5015
rect 10517 4981 10551 5015
rect 10885 4981 10919 5015
rect 12817 4981 12851 5015
rect 12909 4981 12943 5015
rect 8953 4777 8987 4811
rect 11253 4777 11287 4811
rect 12449 4777 12483 4811
rect 13277 4777 13311 4811
rect 4537 4709 4571 4743
rect 10057 4709 10091 4743
rect 10149 4709 10183 4743
rect 12541 4709 12575 4743
rect 1409 4641 1443 4675
rect 2145 4641 2179 4675
rect 2401 4641 2435 4675
rect 4445 4641 4479 4675
rect 5540 4641 5574 4675
rect 7113 4641 7147 4675
rect 7380 4641 7414 4675
rect 13645 4641 13679 4675
rect 14473 4641 14507 4675
rect 4721 4573 4755 4607
rect 5273 4573 5307 4607
rect 10241 4573 10275 4607
rect 11345 4573 11379 4607
rect 11437 4573 11471 4607
rect 12633 4573 12667 4607
rect 13737 4573 13771 4607
rect 13829 4573 13863 4607
rect 3525 4505 3559 4539
rect 8493 4505 8527 4539
rect 12081 4505 12115 4539
rect 1593 4437 1627 4471
rect 4077 4437 4111 4471
rect 6653 4437 6687 4471
rect 9689 4437 9723 4471
rect 10885 4437 10919 4471
rect 14657 4437 14691 4471
rect 9873 4233 9907 4267
rect 11069 4233 11103 4267
rect 1869 4165 1903 4199
rect 4445 4165 4479 4199
rect 13645 4165 13679 4199
rect 15025 4165 15059 4199
rect 2421 4097 2455 4131
rect 4905 4097 4939 4131
rect 9321 4097 9355 4131
rect 10425 4097 10459 4131
rect 11621 4097 11655 4131
rect 12909 4097 12943 4131
rect 13093 4097 13127 4131
rect 14105 4097 14139 4131
rect 14289 4097 14323 4131
rect 3065 4029 3099 4063
rect 6837 4029 6871 4063
rect 9137 4029 9171 4063
rect 10241 4029 10275 4063
rect 11437 4029 11471 4063
rect 12817 4029 12851 4063
rect 14841 4029 14875 4063
rect 3332 3961 3366 3995
rect 5172 3961 5206 3995
rect 7082 3961 7116 3995
rect 11529 3961 11563 3995
rect 14013 3961 14047 3995
rect 2237 3893 2271 3927
rect 2329 3893 2363 3927
rect 6285 3893 6319 3927
rect 8217 3893 8251 3927
rect 8677 3893 8711 3927
rect 9045 3893 9079 3927
rect 10333 3893 10367 3927
rect 12449 3893 12483 3927
rect 1593 3689 1627 3723
rect 1961 3689 1995 3723
rect 2053 3689 2087 3723
rect 2789 3689 2823 3723
rect 8953 3689 8987 3723
rect 12449 3689 12483 3723
rect 3157 3621 3191 3655
rect 4905 3621 4939 3655
rect 6000 3621 6034 3655
rect 12541 3621 12575 3655
rect 13645 3621 13679 3655
rect 3249 3553 3283 3587
rect 4997 3553 5031 3587
rect 7573 3553 7607 3587
rect 7840 3553 7874 3587
rect 10057 3553 10091 3587
rect 10149 3553 10183 3587
rect 11253 3553 11287 3587
rect 13737 3553 13771 3587
rect 14473 3553 14507 3587
rect 2145 3485 2179 3519
rect 3433 3485 3467 3519
rect 5135 3485 5169 3519
rect 5733 3485 5767 3519
rect 10241 3485 10275 3519
rect 11345 3485 11379 3519
rect 11529 3485 11563 3519
rect 12633 3485 12667 3519
rect 13921 3485 13955 3519
rect 9689 3417 9723 3451
rect 14657 3417 14691 3451
rect 4537 3349 4571 3383
rect 7113 3349 7147 3383
rect 10885 3349 10919 3383
rect 12081 3349 12115 3383
rect 13277 3349 13311 3383
rect 2513 3145 2547 3179
rect 3709 3145 3743 3179
rect 9873 3145 9907 3179
rect 13645 3145 13679 3179
rect 8217 3077 8251 3111
rect 15025 3077 15059 3111
rect 3157 3009 3191 3043
rect 4169 3009 4203 3043
rect 4353 3009 4387 3043
rect 6837 3009 6871 3043
rect 9137 3009 9171 3043
rect 9321 3009 9355 3043
rect 10425 3009 10459 3043
rect 11621 3009 11655 3043
rect 13093 3009 13127 3043
rect 14105 3009 14139 3043
rect 14289 3009 14323 3043
rect 1593 2941 1627 2975
rect 4077 2941 4111 2975
rect 4905 2941 4939 2975
rect 5161 2941 5195 2975
rect 11529 2941 11563 2975
rect 14841 2941 14875 2975
rect 1869 2873 1903 2907
rect 2973 2873 3007 2907
rect 7082 2873 7116 2907
rect 10333 2873 10367 2907
rect 12817 2873 12851 2907
rect 2881 2805 2915 2839
rect 6285 2805 6319 2839
rect 8677 2805 8711 2839
rect 9045 2805 9079 2839
rect 9781 2805 9815 2839
rect 10241 2805 10275 2839
rect 11069 2805 11103 2839
rect 11437 2805 11471 2839
rect 12449 2805 12483 2839
rect 12909 2805 12943 2839
rect 14013 2805 14047 2839
rect 6377 2601 6411 2635
rect 6929 2601 6963 2635
rect 7389 2601 7423 2635
rect 8125 2601 8159 2635
rect 10241 2601 10275 2635
rect 10977 2601 11011 2635
rect 11345 2601 11379 2635
rect 12173 2601 12207 2635
rect 13093 2601 13127 2635
rect 14289 2601 14323 2635
rect 5242 2533 5276 2567
rect 10149 2533 10183 2567
rect 13001 2533 13035 2567
rect 1409 2465 1443 2499
rect 2145 2465 2179 2499
rect 2412 2465 2446 2499
rect 4077 2465 4111 2499
rect 7297 2465 7331 2499
rect 8493 2465 8527 2499
rect 9505 2465 9539 2499
rect 12357 2465 12391 2499
rect 14197 2465 14231 2499
rect 15209 2465 15243 2499
rect 4353 2397 4387 2431
rect 4997 2397 5031 2431
rect 7481 2397 7515 2431
rect 8585 2397 8619 2431
rect 8677 2397 8711 2431
rect 10333 2397 10367 2431
rect 11437 2397 11471 2431
rect 11529 2397 11563 2431
rect 13185 2397 13219 2431
rect 14381 2397 14415 2431
rect 12633 2329 12667 2363
rect 1593 2261 1627 2295
rect 3525 2261 3559 2295
rect 9321 2261 9355 2295
rect 9781 2261 9815 2295
rect 13829 2261 13863 2295
rect 15025 2261 15059 2295
rect 949 1989 983 2023
<< metal1 >>
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 12342 18068 12348 18080
rect 9824 18040 12348 18068
rect 9824 18028 9830 18040
rect 12342 18028 12348 18040
rect 12400 18028 12406 18080
rect 8864 17972 9904 18000
rect 4062 17892 4068 17944
rect 4120 17932 4126 17944
rect 8864 17932 8892 17972
rect 4120 17904 8892 17932
rect 4120 17892 4126 17904
rect 8938 17892 8944 17944
rect 8996 17932 9002 17944
rect 9769 17935 9827 17941
rect 9769 17932 9781 17935
rect 8996 17904 9781 17932
rect 8996 17892 9002 17904
rect 9769 17901 9781 17904
rect 9815 17901 9827 17935
rect 9876 17932 9904 17972
rect 10502 17960 10508 18012
rect 10560 18000 10566 18012
rect 13354 18000 13360 18012
rect 10560 17972 13360 18000
rect 10560 17960 10566 17972
rect 13354 17960 13360 17972
rect 13412 17960 13418 18012
rect 10045 17935 10103 17941
rect 9876 17904 9996 17932
rect 9769 17895 9827 17901
rect 3510 17824 3516 17876
rect 3568 17864 3574 17876
rect 9490 17864 9496 17876
rect 3568 17836 9496 17864
rect 3568 17824 3574 17836
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 9968 17864 9996 17904
rect 10045 17901 10057 17935
rect 10091 17932 10103 17935
rect 12802 17932 12808 17944
rect 10091 17904 12808 17932
rect 10091 17901 10103 17904
rect 10045 17895 10103 17901
rect 12802 17892 12808 17904
rect 12860 17892 12866 17944
rect 9968 17836 11376 17864
rect 7834 17756 7840 17808
rect 7892 17796 7898 17808
rect 11149 17799 11207 17805
rect 11149 17796 11161 17799
rect 7892 17768 11161 17796
rect 7892 17756 7898 17768
rect 11149 17765 11161 17768
rect 11195 17765 11207 17799
rect 11149 17759 11207 17765
rect 5534 17688 5540 17740
rect 5592 17728 5598 17740
rect 11238 17728 11244 17740
rect 5592 17700 11244 17728
rect 5592 17688 5598 17700
rect 11238 17688 11244 17700
rect 11296 17688 11302 17740
rect 11348 17728 11376 17836
rect 11517 17799 11575 17805
rect 11517 17765 11529 17799
rect 11563 17796 11575 17799
rect 14550 17796 14556 17808
rect 11563 17768 14556 17796
rect 11563 17765 11575 17768
rect 11517 17759 11575 17765
rect 14550 17756 14556 17768
rect 14608 17756 14614 17808
rect 13170 17728 13176 17740
rect 11348 17700 13176 17728
rect 13170 17688 13176 17700
rect 13228 17688 13234 17740
rect 6914 17620 6920 17672
rect 6972 17660 6978 17672
rect 14274 17660 14280 17672
rect 6972 17632 14280 17660
rect 6972 17620 6978 17632
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 5442 17552 5448 17604
rect 5500 17592 5506 17604
rect 12710 17592 12716 17604
rect 5500 17564 12716 17592
rect 5500 17552 5506 17564
rect 12710 17552 12716 17564
rect 12768 17552 12774 17604
rect 3142 17484 3148 17536
rect 3200 17524 3206 17536
rect 4246 17524 4252 17536
rect 3200 17496 4252 17524
rect 3200 17484 3206 17496
rect 4246 17484 4252 17496
rect 4304 17484 4310 17536
rect 7190 17484 7196 17536
rect 7248 17524 7254 17536
rect 12894 17524 12900 17536
rect 7248 17496 12900 17524
rect 7248 17484 7254 17496
rect 12894 17484 12900 17496
rect 12952 17484 12958 17536
rect 1104 17434 15824 17456
rect 1104 17382 3447 17434
rect 3499 17382 3511 17434
rect 3563 17382 3575 17434
rect 3627 17382 3639 17434
rect 3691 17382 8378 17434
rect 8430 17382 8442 17434
rect 8494 17382 8506 17434
rect 8558 17382 8570 17434
rect 8622 17382 13308 17434
rect 13360 17382 13372 17434
rect 13424 17382 13436 17434
rect 13488 17382 13500 17434
rect 13552 17382 15824 17434
rect 1104 17360 15824 17382
rect 7558 17280 7564 17332
rect 7616 17320 7622 17332
rect 12805 17323 12863 17329
rect 12805 17320 12817 17323
rect 7616 17292 12817 17320
rect 7616 17280 7622 17292
rect 12805 17289 12817 17292
rect 12851 17289 12863 17323
rect 12805 17283 12863 17289
rect 12894 17280 12900 17332
rect 12952 17320 12958 17332
rect 13541 17323 13599 17329
rect 13541 17320 13553 17323
rect 12952 17292 13553 17320
rect 12952 17280 12958 17292
rect 13541 17289 13553 17292
rect 13587 17289 13599 17323
rect 13541 17283 13599 17289
rect 2406 17212 2412 17264
rect 2464 17252 2470 17264
rect 2464 17224 2636 17252
rect 2464 17212 2470 17224
rect 750 17144 756 17196
rect 808 17184 814 17196
rect 1765 17187 1823 17193
rect 808 17156 1624 17184
rect 808 17144 814 17156
rect 1486 17116 1492 17128
rect 1447 17088 1492 17116
rect 1486 17076 1492 17088
rect 1544 17076 1550 17128
rect 1596 17116 1624 17156
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 2130 17184 2136 17196
rect 1811 17156 2136 17184
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 2130 17144 2136 17156
rect 2188 17144 2194 17196
rect 2608 17193 2636 17224
rect 4062 17212 4068 17264
rect 4120 17212 4126 17264
rect 6178 17212 6184 17264
rect 6236 17252 6242 17264
rect 10226 17252 10232 17264
rect 6236 17224 10232 17252
rect 6236 17212 6242 17224
rect 10226 17212 10232 17224
rect 10284 17212 10290 17264
rect 10689 17255 10747 17261
rect 10689 17221 10701 17255
rect 10735 17221 10747 17255
rect 10689 17215 10747 17221
rect 2593 17187 2651 17193
rect 2593 17153 2605 17187
rect 2639 17153 2651 17187
rect 2593 17147 2651 17153
rect 2406 17116 2412 17128
rect 1596 17088 2412 17116
rect 2406 17076 2412 17088
rect 2464 17076 2470 17128
rect 3694 17076 3700 17128
rect 3752 17116 3758 17128
rect 4080 17125 4108 17212
rect 4246 17184 4252 17196
rect 4207 17156 4252 17184
rect 4246 17144 4252 17156
rect 4304 17144 4310 17196
rect 6273 17187 6331 17193
rect 6273 17153 6285 17187
rect 6319 17184 6331 17187
rect 7282 17184 7288 17196
rect 6319 17156 7288 17184
rect 6319 17153 6331 17156
rect 6273 17147 6331 17153
rect 7282 17144 7288 17156
rect 7340 17144 7346 17196
rect 7466 17184 7472 17196
rect 7427 17156 7472 17184
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 8665 17187 8723 17193
rect 8665 17184 8677 17187
rect 8128 17156 8677 17184
rect 4065 17119 4123 17125
rect 4065 17116 4077 17119
rect 3752 17088 4077 17116
rect 3752 17076 3758 17088
rect 4065 17085 4077 17088
rect 4111 17085 4123 17119
rect 7300 17116 7328 17144
rect 8128 17116 8156 17156
rect 8665 17153 8677 17156
rect 8711 17153 8723 17187
rect 10134 17184 10140 17196
rect 8665 17147 8723 17153
rect 9324 17156 10140 17184
rect 7300 17088 8156 17116
rect 8481 17119 8539 17125
rect 4065 17079 4123 17085
rect 8481 17085 8493 17119
rect 8527 17116 8539 17119
rect 9324 17116 9352 17156
rect 10134 17144 10140 17156
rect 10192 17144 10198 17196
rect 9490 17116 9496 17128
rect 8527 17088 9352 17116
rect 9451 17088 9496 17116
rect 8527 17085 8539 17088
rect 8481 17079 8539 17085
rect 9490 17076 9496 17088
rect 9548 17076 9554 17128
rect 9769 17119 9827 17125
rect 9769 17085 9781 17119
rect 9815 17116 9827 17119
rect 10042 17116 10048 17128
rect 9815 17088 10048 17116
rect 9815 17085 9827 17088
rect 9769 17079 9827 17085
rect 10042 17076 10048 17088
rect 10100 17076 10106 17128
rect 10410 17076 10416 17128
rect 10468 17116 10474 17128
rect 10505 17119 10563 17125
rect 10505 17116 10517 17119
rect 10468 17088 10517 17116
rect 10468 17076 10474 17088
rect 10505 17085 10517 17088
rect 10551 17085 10563 17119
rect 10704 17116 10732 17215
rect 10505 17079 10563 17085
rect 10612 17088 10732 17116
rect 11241 17119 11299 17125
rect 3142 17008 3148 17060
rect 3200 17048 3206 17060
rect 6270 17048 6276 17060
rect 3200 17020 6276 17048
rect 3200 17008 3206 17020
rect 6270 17008 6276 17020
rect 6328 17008 6334 17060
rect 7377 17051 7435 17057
rect 7377 17017 7389 17051
rect 7423 17048 7435 17051
rect 9122 17048 9128 17060
rect 7423 17020 9128 17048
rect 7423 17017 7435 17020
rect 7377 17011 7435 17017
rect 9122 17008 9128 17020
rect 9180 17008 9186 17060
rect 9674 17008 9680 17060
rect 9732 17048 9738 17060
rect 10612 17048 10640 17088
rect 11241 17085 11253 17119
rect 11287 17116 11299 17119
rect 12434 17116 12440 17128
rect 11287 17088 12440 17116
rect 11287 17085 11299 17088
rect 11241 17079 11299 17085
rect 12434 17076 12440 17088
rect 12492 17076 12498 17128
rect 12621 17119 12679 17125
rect 12621 17085 12633 17119
rect 12667 17116 12679 17119
rect 12894 17116 12900 17128
rect 12667 17088 12900 17116
rect 12667 17085 12679 17088
rect 12621 17079 12679 17085
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 13354 17116 13360 17128
rect 13315 17088 13360 17116
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 9732 17020 10640 17048
rect 9732 17008 9738 17020
rect 3237 16983 3295 16989
rect 3237 16949 3249 16983
rect 3283 16980 3295 16983
rect 3326 16980 3332 16992
rect 3283 16952 3332 16980
rect 3283 16949 3295 16952
rect 3237 16943 3295 16949
rect 3326 16940 3332 16952
rect 3384 16940 3390 16992
rect 4893 16983 4951 16989
rect 4893 16949 4905 16983
rect 4939 16980 4951 16983
rect 4982 16980 4988 16992
rect 4939 16952 4988 16980
rect 4939 16949 4951 16952
rect 4893 16943 4951 16949
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 5626 16980 5632 16992
rect 5587 16952 5632 16980
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 5718 16940 5724 16992
rect 5776 16980 5782 16992
rect 5997 16983 6055 16989
rect 5997 16980 6009 16983
rect 5776 16952 6009 16980
rect 5776 16940 5782 16952
rect 5997 16949 6009 16952
rect 6043 16949 6055 16983
rect 5997 16943 6055 16949
rect 6089 16983 6147 16989
rect 6089 16949 6101 16983
rect 6135 16980 6147 16983
rect 6917 16983 6975 16989
rect 6917 16980 6929 16983
rect 6135 16952 6929 16980
rect 6135 16949 6147 16952
rect 6089 16943 6147 16949
rect 6917 16949 6929 16952
rect 6963 16949 6975 16983
rect 6917 16943 6975 16949
rect 7285 16983 7343 16989
rect 7285 16949 7297 16983
rect 7331 16980 7343 16983
rect 7650 16980 7656 16992
rect 7331 16952 7656 16980
rect 7331 16949 7343 16952
rect 7285 16943 7343 16949
rect 7650 16940 7656 16952
rect 7708 16940 7714 16992
rect 8110 16980 8116 16992
rect 8071 16952 8116 16980
rect 8110 16940 8116 16952
rect 8168 16940 8174 16992
rect 8570 16980 8576 16992
rect 8531 16952 8576 16980
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 9306 16980 9312 16992
rect 9267 16952 9312 16980
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 9398 16940 9404 16992
rect 9456 16980 9462 16992
rect 9953 16983 10011 16989
rect 9953 16980 9965 16983
rect 9456 16952 9965 16980
rect 9456 16940 9462 16952
rect 9953 16949 9965 16952
rect 9999 16949 10011 16983
rect 9953 16943 10011 16949
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 11425 16983 11483 16989
rect 11425 16980 11437 16983
rect 10284 16952 11437 16980
rect 10284 16940 10290 16952
rect 11425 16949 11437 16952
rect 11471 16949 11483 16983
rect 11425 16943 11483 16949
rect 1104 16890 15824 16912
rect 1104 16838 5912 16890
rect 5964 16838 5976 16890
rect 6028 16838 6040 16890
rect 6092 16838 6104 16890
rect 6156 16838 10843 16890
rect 10895 16838 10907 16890
rect 10959 16838 10971 16890
rect 11023 16838 11035 16890
rect 11087 16838 15824 16890
rect 1104 16816 15824 16838
rect 2501 16779 2559 16785
rect 2501 16745 2513 16779
rect 2547 16745 2559 16779
rect 2501 16739 2559 16745
rect 1670 16708 1676 16720
rect 1631 16680 1676 16708
rect 1670 16668 1676 16680
rect 1728 16668 1734 16720
rect 2516 16708 2544 16739
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 3697 16779 3755 16785
rect 2832 16748 3096 16776
rect 2832 16736 2838 16748
rect 3068 16717 3096 16748
rect 3697 16745 3709 16779
rect 3743 16776 3755 16779
rect 4890 16776 4896 16788
rect 3743 16748 4896 16776
rect 3743 16745 3755 16748
rect 3697 16739 3755 16745
rect 4890 16736 4896 16748
rect 4948 16736 4954 16788
rect 4985 16779 5043 16785
rect 4985 16745 4997 16779
rect 5031 16745 5043 16779
rect 4985 16739 5043 16745
rect 3053 16711 3111 16717
rect 2516 16680 3004 16708
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 2682 16640 2688 16652
rect 1443 16612 2544 16640
rect 2643 16612 2688 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 2516 16572 2544 16612
rect 2682 16600 2688 16612
rect 2740 16600 2746 16652
rect 2774 16600 2780 16652
rect 2832 16640 2838 16652
rect 2976 16640 3004 16680
rect 3053 16677 3065 16711
rect 3099 16677 3111 16711
rect 3053 16671 3111 16677
rect 3712 16680 4200 16708
rect 3712 16640 3740 16680
rect 3878 16640 3884 16652
rect 2832 16612 2877 16640
rect 2976 16612 3740 16640
rect 3839 16612 3884 16640
rect 2832 16600 2838 16612
rect 3878 16600 3884 16612
rect 3936 16600 3942 16652
rect 3970 16600 3976 16652
rect 4028 16640 4034 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 4028 16612 4077 16640
rect 4028 16600 4034 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 3326 16572 3332 16584
rect 2516 16544 3332 16572
rect 3326 16532 3332 16544
rect 3384 16572 3390 16584
rect 3694 16572 3700 16584
rect 3384 16544 3700 16572
rect 3384 16532 3390 16544
rect 3694 16532 3700 16544
rect 3752 16532 3758 16584
rect 4172 16572 4200 16680
rect 4430 16668 4436 16720
rect 4488 16708 4494 16720
rect 5000 16708 5028 16739
rect 5350 16736 5356 16788
rect 5408 16776 5414 16788
rect 5445 16779 5503 16785
rect 5445 16776 5457 16779
rect 5408 16748 5457 16776
rect 5408 16736 5414 16748
rect 5445 16745 5457 16748
rect 5491 16745 5503 16779
rect 6270 16776 6276 16788
rect 6231 16748 6276 16776
rect 5445 16739 5503 16745
rect 6270 16736 6276 16748
rect 6328 16736 6334 16788
rect 6641 16779 6699 16785
rect 6641 16745 6653 16779
rect 6687 16776 6699 16779
rect 7469 16779 7527 16785
rect 7469 16776 7481 16779
rect 6687 16748 7481 16776
rect 6687 16745 6699 16748
rect 6641 16739 6699 16745
rect 7469 16745 7481 16748
rect 7515 16745 7527 16779
rect 7834 16776 7840 16788
rect 7795 16748 7840 16776
rect 7469 16739 7527 16745
rect 7834 16736 7840 16748
rect 7892 16736 7898 16788
rect 7929 16779 7987 16785
rect 7929 16745 7941 16779
rect 7975 16776 7987 16779
rect 8938 16776 8944 16788
rect 7975 16748 8944 16776
rect 7975 16745 7987 16748
rect 7929 16739 7987 16745
rect 8938 16736 8944 16748
rect 8996 16736 9002 16788
rect 9582 16736 9588 16788
rect 9640 16776 9646 16788
rect 9861 16779 9919 16785
rect 9861 16776 9873 16779
rect 9640 16748 9873 16776
rect 9640 16736 9646 16748
rect 9861 16745 9873 16748
rect 9907 16745 9919 16779
rect 9861 16739 9919 16745
rect 10597 16779 10655 16785
rect 10597 16745 10609 16779
rect 10643 16745 10655 16779
rect 10597 16739 10655 16745
rect 6733 16711 6791 16717
rect 4488 16680 5028 16708
rect 5276 16680 6684 16708
rect 4488 16668 4494 16680
rect 4246 16600 4252 16652
rect 4304 16640 4310 16652
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 4304 16612 4353 16640
rect 4304 16600 4310 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 4522 16600 4528 16652
rect 4580 16640 4586 16652
rect 5276 16640 5304 16680
rect 4580 16612 5304 16640
rect 5353 16643 5411 16649
rect 4580 16600 4586 16612
rect 5353 16609 5365 16643
rect 5399 16640 5411 16643
rect 5442 16640 5448 16652
rect 5399 16612 5448 16640
rect 5399 16609 5411 16612
rect 5353 16603 5411 16609
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 6656 16640 6684 16680
rect 6733 16677 6745 16711
rect 6779 16708 6791 16711
rect 8110 16708 8116 16720
rect 6779 16680 8116 16708
rect 6779 16677 6791 16680
rect 6733 16671 6791 16677
rect 8110 16668 8116 16680
rect 8168 16668 8174 16720
rect 10612 16708 10640 16739
rect 12158 16736 12164 16788
rect 12216 16776 12222 16788
rect 13541 16779 13599 16785
rect 13541 16776 13553 16779
rect 12216 16748 13553 16776
rect 12216 16736 12222 16748
rect 13541 16745 13553 16748
rect 13587 16745 13599 16779
rect 14274 16776 14280 16788
rect 14235 16748 14280 16776
rect 13541 16739 13599 16745
rect 14274 16736 14280 16748
rect 14332 16736 14338 16788
rect 8496 16680 10640 16708
rect 8496 16640 8524 16680
rect 12066 16668 12072 16720
rect 12124 16708 12130 16720
rect 12124 16680 13400 16708
rect 12124 16668 12130 16680
rect 8662 16640 8668 16652
rect 6656 16612 8524 16640
rect 8623 16612 8668 16640
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 8846 16600 8852 16652
rect 8904 16640 8910 16652
rect 8941 16643 8999 16649
rect 8941 16640 8953 16643
rect 8904 16612 8953 16640
rect 8904 16600 8910 16612
rect 8941 16609 8953 16612
rect 8987 16609 8999 16643
rect 8941 16603 8999 16609
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16640 10471 16643
rect 10502 16640 10508 16652
rect 10459 16612 10508 16640
rect 10459 16609 10471 16612
rect 10413 16603 10471 16609
rect 4706 16572 4712 16584
rect 4172 16544 4712 16572
rect 4706 16532 4712 16544
rect 4764 16532 4770 16584
rect 5074 16532 5080 16584
rect 5132 16572 5138 16584
rect 5537 16575 5595 16581
rect 5537 16572 5549 16575
rect 5132 16544 5549 16572
rect 5132 16532 5138 16544
rect 5537 16541 5549 16544
rect 5583 16541 5595 16575
rect 5537 16535 5595 16541
rect 6086 16532 6092 16584
rect 6144 16572 6150 16584
rect 6825 16575 6883 16581
rect 6825 16572 6837 16575
rect 6144 16544 6837 16572
rect 6144 16532 6150 16544
rect 6825 16541 6837 16544
rect 6871 16541 6883 16575
rect 6825 16535 6883 16541
rect 7282 16532 7288 16584
rect 7340 16572 7346 16584
rect 7742 16572 7748 16584
rect 7340 16544 7748 16572
rect 7340 16532 7346 16544
rect 7742 16532 7748 16544
rect 7800 16572 7806 16584
rect 8021 16575 8079 16581
rect 8021 16572 8033 16575
rect 7800 16544 8033 16572
rect 7800 16532 7806 16544
rect 8021 16541 8033 16544
rect 8067 16541 8079 16575
rect 8021 16535 8079 16541
rect 8110 16532 8116 16584
rect 8168 16572 8174 16584
rect 9030 16572 9036 16584
rect 8168 16544 9036 16572
rect 8168 16532 8174 16544
rect 9030 16532 9036 16544
rect 9088 16532 9094 16584
rect 1486 16464 1492 16516
rect 1544 16504 1550 16516
rect 3786 16504 3792 16516
rect 1544 16476 3792 16504
rect 1544 16464 1550 16476
rect 3786 16464 3792 16476
rect 3844 16464 3850 16516
rect 4338 16464 4344 16516
rect 4396 16504 4402 16516
rect 9398 16504 9404 16516
rect 4396 16476 9404 16504
rect 4396 16464 4402 16476
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 2314 16396 2320 16448
rect 2372 16436 2378 16448
rect 4430 16436 4436 16448
rect 2372 16408 4436 16436
rect 2372 16396 2378 16408
rect 4430 16396 4436 16408
rect 4488 16396 4494 16448
rect 4798 16396 4804 16448
rect 4856 16436 4862 16448
rect 9582 16436 9588 16448
rect 4856 16408 9588 16436
rect 4856 16396 4862 16408
rect 9582 16396 9588 16408
rect 9640 16396 9646 16448
rect 9692 16436 9720 16603
rect 10502 16600 10508 16612
rect 10560 16600 10566 16652
rect 10962 16600 10968 16652
rect 11020 16640 11026 16652
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 11020 16612 11161 16640
rect 11020 16600 11026 16612
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 11149 16603 11207 16609
rect 11256 16612 11897 16640
rect 9858 16532 9864 16584
rect 9916 16572 9922 16584
rect 10778 16572 10784 16584
rect 9916 16544 10784 16572
rect 9916 16532 9922 16544
rect 10778 16532 10784 16544
rect 10836 16532 10842 16584
rect 11256 16572 11284 16612
rect 11885 16609 11897 16612
rect 11931 16609 11943 16643
rect 11885 16603 11943 16609
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 13372 16649 13400 16680
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 12584 16612 12633 16640
rect 12584 16600 12590 16612
rect 12621 16609 12633 16612
rect 12667 16609 12679 16643
rect 12621 16603 12679 16609
rect 13357 16643 13415 16649
rect 13357 16609 13369 16643
rect 13403 16609 13415 16643
rect 13357 16603 13415 16609
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 11164 16544 11284 16572
rect 11164 16516 11192 16544
rect 11422 16532 11428 16584
rect 11480 16572 11486 16584
rect 14108 16572 14136 16603
rect 11480 16544 14136 16572
rect 11480 16532 11486 16544
rect 11146 16464 11152 16516
rect 11204 16464 11210 16516
rect 11238 16464 11244 16516
rect 11296 16504 11302 16516
rect 11333 16507 11391 16513
rect 11333 16504 11345 16507
rect 11296 16476 11345 16504
rect 11296 16464 11302 16476
rect 11333 16473 11345 16476
rect 11379 16473 11391 16507
rect 11333 16467 11391 16473
rect 11882 16464 11888 16516
rect 11940 16504 11946 16516
rect 12069 16507 12127 16513
rect 12069 16504 12081 16507
rect 11940 16476 12081 16504
rect 11940 16464 11946 16476
rect 12069 16473 12081 16476
rect 12115 16473 12127 16507
rect 12802 16504 12808 16516
rect 12763 16476 12808 16504
rect 12069 16467 12127 16473
rect 12802 16464 12808 16476
rect 12860 16464 12866 16516
rect 10226 16436 10232 16448
rect 9692 16408 10232 16436
rect 10226 16396 10232 16408
rect 10284 16396 10290 16448
rect 10318 16396 10324 16448
rect 10376 16436 10382 16448
rect 14366 16436 14372 16448
rect 10376 16408 14372 16436
rect 10376 16396 10382 16408
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 1104 16346 15824 16368
rect 1104 16294 3447 16346
rect 3499 16294 3511 16346
rect 3563 16294 3575 16346
rect 3627 16294 3639 16346
rect 3691 16294 8378 16346
rect 8430 16294 8442 16346
rect 8494 16294 8506 16346
rect 8558 16294 8570 16346
rect 8622 16294 13308 16346
rect 13360 16294 13372 16346
rect 13424 16294 13436 16346
rect 13488 16294 13500 16346
rect 13552 16294 15824 16346
rect 1104 16272 15824 16294
rect 1118 16192 1124 16244
rect 1176 16232 1182 16244
rect 2498 16232 2504 16244
rect 1176 16204 2504 16232
rect 1176 16192 1182 16204
rect 2498 16192 2504 16204
rect 2556 16232 2562 16244
rect 2774 16232 2780 16244
rect 2556 16204 2780 16232
rect 2556 16192 2562 16204
rect 2774 16192 2780 16204
rect 2832 16192 2838 16244
rect 5537 16235 5595 16241
rect 5537 16201 5549 16235
rect 5583 16201 5595 16235
rect 5537 16195 5595 16201
rect 3418 16124 3424 16176
rect 3476 16164 3482 16176
rect 5552 16164 5580 16195
rect 6638 16192 6644 16244
rect 6696 16232 6702 16244
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 6696 16204 8033 16232
rect 6696 16192 6702 16204
rect 8021 16201 8033 16204
rect 8067 16201 8079 16235
rect 8021 16195 8079 16201
rect 8754 16192 8760 16244
rect 8812 16232 8818 16244
rect 8812 16204 9904 16232
rect 8812 16192 8818 16204
rect 3476 16136 5580 16164
rect 3476 16124 3482 16136
rect 7006 16124 7012 16176
rect 7064 16164 7070 16176
rect 7064 16136 8616 16164
rect 7064 16124 7070 16136
rect 1394 16056 1400 16108
rect 1452 16096 1458 16108
rect 1673 16099 1731 16105
rect 1673 16096 1685 16099
rect 1452 16068 1685 16096
rect 1452 16056 1458 16068
rect 1673 16065 1685 16068
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 1762 16056 1768 16108
rect 1820 16096 1826 16108
rect 2593 16099 2651 16105
rect 2593 16096 2605 16099
rect 1820 16068 2605 16096
rect 1820 16056 1826 16068
rect 2593 16065 2605 16068
rect 2639 16065 2651 16099
rect 2593 16059 2651 16065
rect 4062 16056 4068 16108
rect 4120 16096 4126 16108
rect 4985 16099 5043 16105
rect 4120 16068 4660 16096
rect 4120 16056 4126 16068
rect 106 15988 112 16040
rect 164 16028 170 16040
rect 1302 16028 1308 16040
rect 164 16000 1308 16028
rect 164 15988 170 16000
rect 1302 15988 1308 16000
rect 1360 16028 1366 16040
rect 1489 16031 1547 16037
rect 1489 16028 1501 16031
rect 1360 16000 1501 16028
rect 1360 15988 1366 16000
rect 1489 15997 1501 16000
rect 1535 15997 1547 16031
rect 1489 15991 1547 15997
rect 2409 16031 2467 16037
rect 2409 15997 2421 16031
rect 2455 16028 2467 16031
rect 3234 16028 3240 16040
rect 2455 16000 3240 16028
rect 2455 15997 2467 16000
rect 2409 15991 2467 15997
rect 382 15920 388 15972
rect 440 15960 446 15972
rect 2424 15960 2452 15991
rect 3234 15988 3240 16000
rect 3292 15988 3298 16040
rect 3329 16031 3387 16037
rect 3329 15997 3341 16031
rect 3375 16028 3387 16031
rect 4430 16028 4436 16040
rect 3375 16000 4436 16028
rect 3375 15997 3387 16000
rect 3329 15991 3387 15997
rect 4430 15988 4436 16000
rect 4488 15988 4494 16040
rect 3602 15960 3608 15972
rect 440 15932 2452 15960
rect 3563 15932 3608 15960
rect 440 15920 446 15932
rect 3602 15920 3608 15932
rect 3660 15920 3666 15972
rect 4246 15920 4252 15972
rect 4304 15960 4310 15972
rect 4632 15960 4660 16068
rect 4985 16065 4997 16099
rect 5031 16096 5043 16099
rect 5534 16096 5540 16108
rect 5031 16068 5540 16096
rect 5031 16065 5043 16068
rect 4985 16059 5043 16065
rect 5534 16056 5540 16068
rect 5592 16056 5598 16108
rect 5626 16056 5632 16108
rect 5684 16096 5690 16108
rect 5997 16099 6055 16105
rect 5997 16096 6009 16099
rect 5684 16068 6009 16096
rect 5684 16056 5690 16068
rect 5997 16065 6009 16068
rect 6043 16065 6055 16099
rect 5997 16059 6055 16065
rect 6086 16056 6092 16108
rect 6144 16096 6150 16108
rect 7374 16096 7380 16108
rect 6144 16068 6189 16096
rect 7335 16068 7380 16096
rect 6144 16056 6150 16068
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 8588 16105 8616 16136
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16065 8631 16099
rect 8573 16059 8631 16065
rect 9398 16056 9404 16108
rect 9456 16096 9462 16108
rect 9769 16099 9827 16105
rect 9769 16096 9781 16099
rect 9456 16068 9781 16096
rect 9456 16056 9462 16068
rect 9769 16065 9781 16068
rect 9815 16065 9827 16099
rect 9876 16096 9904 16204
rect 9950 16192 9956 16244
rect 10008 16232 10014 16244
rect 10597 16235 10655 16241
rect 10597 16232 10609 16235
rect 10008 16204 10609 16232
rect 10008 16192 10014 16204
rect 10597 16201 10609 16204
rect 10643 16201 10655 16235
rect 10597 16195 10655 16201
rect 10778 16192 10784 16244
rect 10836 16232 10842 16244
rect 13357 16235 13415 16241
rect 13357 16232 13369 16235
rect 10836 16204 13369 16232
rect 10836 16192 10842 16204
rect 13357 16201 13369 16204
rect 13403 16201 13415 16235
rect 13357 16195 13415 16201
rect 14182 16192 14188 16244
rect 14240 16232 14246 16244
rect 15102 16232 15108 16244
rect 14240 16204 15108 16232
rect 14240 16192 14246 16204
rect 15102 16192 15108 16204
rect 15160 16232 15166 16244
rect 16390 16232 16396 16244
rect 15160 16204 16396 16232
rect 15160 16192 15166 16204
rect 16390 16192 16396 16204
rect 16448 16192 16454 16244
rect 10502 16124 10508 16176
rect 10560 16164 10566 16176
rect 10962 16164 10968 16176
rect 10560 16136 10968 16164
rect 10560 16124 10566 16136
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 12621 16167 12679 16173
rect 12621 16133 12633 16167
rect 12667 16133 12679 16167
rect 12621 16127 12679 16133
rect 12636 16096 12664 16127
rect 9876 16068 12664 16096
rect 9769 16059 9827 16065
rect 4798 16028 4804 16040
rect 4759 16000 4804 16028
rect 4798 15988 4804 16000
rect 4856 15988 4862 16040
rect 4890 15988 4896 16040
rect 4948 16028 4954 16040
rect 5905 16031 5963 16037
rect 4948 16000 5120 16028
rect 4948 15988 4954 16000
rect 5092 15960 5120 16000
rect 5905 15997 5917 16031
rect 5951 16028 5963 16031
rect 7282 16028 7288 16040
rect 5951 16000 7144 16028
rect 7243 16000 7288 16028
rect 5951 15997 5963 16000
rect 5905 15991 5963 15997
rect 4304 15932 4476 15960
rect 4632 15932 5028 15960
rect 5092 15932 6868 15960
rect 4304 15920 4310 15932
rect 4338 15892 4344 15904
rect 4299 15864 4344 15892
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 4448 15892 4476 15932
rect 4709 15895 4767 15901
rect 4709 15892 4721 15895
rect 4448 15864 4721 15892
rect 4709 15861 4721 15864
rect 4755 15861 4767 15895
rect 5000 15892 5028 15932
rect 6730 15892 6736 15904
rect 5000 15864 6736 15892
rect 4709 15855 4767 15861
rect 6730 15852 6736 15864
rect 6788 15852 6794 15904
rect 6840 15901 6868 15932
rect 6825 15895 6883 15901
rect 6825 15861 6837 15895
rect 6871 15861 6883 15895
rect 7116 15892 7144 16000
rect 7282 15988 7288 16000
rect 7340 15988 7346 16040
rect 8481 16031 8539 16037
rect 8481 15997 8493 16031
rect 8527 16028 8539 16031
rect 9582 16028 9588 16040
rect 8527 16000 9076 16028
rect 9543 16000 9588 16028
rect 8527 15997 8539 16000
rect 8481 15991 8539 15997
rect 7193 15963 7251 15969
rect 7193 15929 7205 15963
rect 7239 15960 7251 15963
rect 8389 15963 8447 15969
rect 7239 15932 8340 15960
rect 7239 15929 7251 15932
rect 7193 15923 7251 15929
rect 7834 15892 7840 15904
rect 7116 15864 7840 15892
rect 6825 15855 6883 15861
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 8312 15892 8340 15932
rect 8389 15929 8401 15963
rect 8435 15960 8447 15963
rect 8754 15960 8760 15972
rect 8435 15932 8760 15960
rect 8435 15929 8447 15932
rect 8389 15923 8447 15929
rect 8754 15920 8760 15932
rect 8812 15920 8818 15972
rect 9048 15960 9076 16000
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 16028 9735 16031
rect 10318 16028 10324 16040
rect 9723 16000 10324 16028
rect 9723 15997 9735 16000
rect 9677 15991 9735 15997
rect 10318 15988 10324 16000
rect 10376 15988 10382 16040
rect 10413 16031 10471 16037
rect 10413 15997 10425 16031
rect 10459 16028 10471 16031
rect 11149 16031 11207 16037
rect 10459 16000 11100 16028
rect 10459 15997 10471 16000
rect 10413 15991 10471 15997
rect 9766 15960 9772 15972
rect 9048 15932 9772 15960
rect 9766 15920 9772 15932
rect 9824 15920 9830 15972
rect 11072 15960 11100 16000
rect 11149 15997 11161 16031
rect 11195 16028 11207 16031
rect 11790 16028 11796 16040
rect 11195 16000 11796 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 11790 15988 11796 16000
rect 11848 15988 11854 16040
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 16028 12495 16031
rect 12710 16028 12716 16040
rect 12483 16000 12716 16028
rect 12483 15997 12495 16000
rect 12437 15991 12495 15997
rect 12710 15988 12716 16000
rect 12768 15988 12774 16040
rect 13170 16028 13176 16040
rect 13131 16000 13176 16028
rect 13170 15988 13176 16000
rect 13228 15988 13234 16040
rect 12342 15960 12348 15972
rect 11072 15932 12348 15960
rect 12342 15920 12348 15932
rect 12400 15920 12406 15972
rect 8938 15892 8944 15904
rect 8312 15864 8944 15892
rect 8938 15852 8944 15864
rect 8996 15852 9002 15904
rect 9030 15852 9036 15904
rect 9088 15892 9094 15904
rect 9217 15895 9275 15901
rect 9217 15892 9229 15895
rect 9088 15864 9229 15892
rect 9088 15852 9094 15864
rect 9217 15861 9229 15864
rect 9263 15861 9275 15895
rect 9217 15855 9275 15861
rect 11146 15852 11152 15904
rect 11204 15892 11210 15904
rect 11333 15895 11391 15901
rect 11333 15892 11345 15895
rect 11204 15864 11345 15892
rect 11204 15852 11210 15864
rect 11333 15861 11345 15864
rect 11379 15861 11391 15895
rect 11333 15855 11391 15861
rect 1104 15802 15824 15824
rect 1104 15750 5912 15802
rect 5964 15750 5976 15802
rect 6028 15750 6040 15802
rect 6092 15750 6104 15802
rect 6156 15750 10843 15802
rect 10895 15750 10907 15802
rect 10959 15750 10971 15802
rect 11023 15750 11035 15802
rect 11087 15750 15824 15802
rect 1104 15728 15824 15750
rect 2958 15648 2964 15700
rect 3016 15688 3022 15700
rect 3421 15691 3479 15697
rect 3421 15688 3433 15691
rect 3016 15660 3433 15688
rect 3016 15648 3022 15660
rect 3421 15657 3433 15660
rect 3467 15657 3479 15691
rect 3421 15651 3479 15657
rect 5166 15648 5172 15700
rect 5224 15688 5230 15700
rect 7193 15691 7251 15697
rect 7193 15688 7205 15691
rect 5224 15660 7205 15688
rect 5224 15648 5230 15660
rect 7193 15657 7205 15660
rect 7239 15688 7251 15691
rect 7374 15688 7380 15700
rect 7239 15660 7380 15688
rect 7239 15657 7251 15660
rect 7193 15651 7251 15657
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 8110 15688 8116 15700
rect 8071 15660 8116 15688
rect 8110 15648 8116 15660
rect 8168 15648 8174 15700
rect 9033 15691 9091 15697
rect 9033 15688 9045 15691
rect 8220 15660 9045 15688
rect 1302 15580 1308 15632
rect 1360 15620 1366 15632
rect 4614 15620 4620 15632
rect 1360 15592 4620 15620
rect 1360 15580 1366 15592
rect 4614 15580 4620 15592
rect 4672 15580 4678 15632
rect 4985 15623 5043 15629
rect 4985 15589 4997 15623
rect 5031 15620 5043 15623
rect 6822 15620 6828 15632
rect 5031 15592 6828 15620
rect 5031 15589 5043 15592
rect 4985 15583 5043 15589
rect 6822 15580 6828 15592
rect 6880 15580 6886 15632
rect 6914 15580 6920 15632
rect 6972 15620 6978 15632
rect 8220 15620 8248 15660
rect 9033 15657 9045 15660
rect 9079 15657 9091 15691
rect 9033 15651 9091 15657
rect 9214 15648 9220 15700
rect 9272 15688 9278 15700
rect 11057 15691 11115 15697
rect 11057 15688 11069 15691
rect 9272 15660 11069 15688
rect 9272 15648 9278 15660
rect 11057 15657 11069 15660
rect 11103 15657 11115 15691
rect 11057 15651 11115 15657
rect 11793 15691 11851 15697
rect 11793 15657 11805 15691
rect 11839 15657 11851 15691
rect 11793 15651 11851 15657
rect 6972 15592 8248 15620
rect 6972 15580 6978 15592
rect 8294 15580 8300 15632
rect 8352 15620 8358 15632
rect 11808 15620 11836 15651
rect 12158 15648 12164 15700
rect 12216 15688 12222 15700
rect 12529 15691 12587 15697
rect 12529 15688 12541 15691
rect 12216 15660 12541 15688
rect 12216 15648 12222 15660
rect 12529 15657 12541 15660
rect 12575 15657 12587 15691
rect 12529 15651 12587 15657
rect 8352 15592 11836 15620
rect 8352 15580 8358 15592
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15521 1455 15555
rect 1397 15515 1455 15521
rect 1302 15444 1308 15496
rect 1360 15484 1366 15496
rect 1412 15484 1440 15515
rect 1486 15512 1492 15564
rect 1544 15552 1550 15564
rect 2317 15555 2375 15561
rect 2317 15552 2329 15555
rect 1544 15524 2329 15552
rect 1544 15512 1550 15524
rect 2317 15521 2329 15524
rect 2363 15521 2375 15555
rect 2317 15515 2375 15521
rect 3237 15555 3295 15561
rect 3237 15521 3249 15555
rect 3283 15552 3295 15555
rect 3326 15552 3332 15564
rect 3283 15524 3332 15552
rect 3283 15521 3295 15524
rect 3237 15515 3295 15521
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 4706 15512 4712 15564
rect 4764 15552 4770 15564
rect 5813 15555 5871 15561
rect 5813 15552 5825 15555
rect 4764 15524 5825 15552
rect 4764 15512 4770 15524
rect 5813 15521 5825 15524
rect 5859 15521 5871 15555
rect 5813 15515 5871 15521
rect 6080 15555 6138 15561
rect 6080 15521 6092 15555
rect 6126 15552 6138 15555
rect 8021 15555 8079 15561
rect 6126 15524 7972 15552
rect 6126 15521 6138 15524
rect 6080 15515 6138 15521
rect 1360 15456 1440 15484
rect 1673 15487 1731 15493
rect 1360 15444 1366 15456
rect 1673 15453 1685 15487
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 1688 15416 1716 15447
rect 2038 15444 2044 15496
rect 2096 15484 2102 15496
rect 2501 15487 2559 15493
rect 2501 15484 2513 15487
rect 2096 15456 2513 15484
rect 2096 15444 2102 15456
rect 2501 15453 2513 15456
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 2590 15444 2596 15496
rect 2648 15484 2654 15496
rect 5077 15487 5135 15493
rect 5077 15484 5089 15487
rect 2648 15456 5089 15484
rect 2648 15444 2654 15456
rect 5077 15453 5089 15456
rect 5123 15453 5135 15487
rect 5077 15447 5135 15453
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15484 5319 15487
rect 5442 15484 5448 15496
rect 5307 15456 5448 15484
rect 5307 15453 5319 15456
rect 5261 15447 5319 15453
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 7944 15484 7972 15524
rect 8021 15521 8033 15555
rect 8067 15552 8079 15555
rect 8110 15552 8116 15564
rect 8067 15524 8116 15552
rect 8067 15521 8079 15524
rect 8021 15515 8079 15521
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 8849 15555 8907 15561
rect 8849 15521 8861 15555
rect 8895 15552 8907 15555
rect 9122 15552 9128 15564
rect 8895 15524 9128 15552
rect 8895 15521 8907 15524
rect 8849 15515 8907 15521
rect 9122 15512 9128 15524
rect 9180 15512 9186 15564
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9732 15524 10057 15552
rect 9732 15512 9738 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10045 15515 10103 15521
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15552 10195 15555
rect 10502 15552 10508 15564
rect 10183 15524 10508 15552
rect 10183 15521 10195 15524
rect 10137 15515 10195 15521
rect 10502 15512 10508 15524
rect 10560 15512 10566 15564
rect 10686 15512 10692 15564
rect 10744 15552 10750 15564
rect 10870 15552 10876 15564
rect 10744 15524 10876 15552
rect 10744 15512 10750 15524
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 11514 15512 11520 15564
rect 11572 15552 11578 15564
rect 11609 15555 11667 15561
rect 11609 15552 11621 15555
rect 11572 15524 11621 15552
rect 11572 15512 11578 15524
rect 11609 15521 11621 15524
rect 11655 15521 11667 15555
rect 11609 15515 11667 15521
rect 11698 15512 11704 15564
rect 11756 15552 11762 15564
rect 12345 15555 12403 15561
rect 12345 15552 12357 15555
rect 11756 15524 12357 15552
rect 11756 15512 11762 15524
rect 12345 15521 12357 15524
rect 12391 15521 12403 15555
rect 12345 15515 12403 15521
rect 8205 15487 8263 15493
rect 8205 15484 8217 15487
rect 7944 15456 8217 15484
rect 8205 15453 8217 15456
rect 8251 15484 8263 15487
rect 9214 15484 9220 15496
rect 8251 15456 9220 15484
rect 8251 15453 8263 15456
rect 8205 15447 8263 15453
rect 9214 15444 9220 15456
rect 9272 15444 9278 15496
rect 9766 15484 9772 15496
rect 9600 15456 9772 15484
rect 2222 15416 2228 15428
rect 1688 15388 2228 15416
rect 2222 15376 2228 15388
rect 2280 15376 2286 15428
rect 3234 15376 3240 15428
rect 3292 15416 3298 15428
rect 5718 15416 5724 15428
rect 3292 15388 5724 15416
rect 3292 15376 3298 15388
rect 5718 15376 5724 15388
rect 5776 15376 5782 15428
rect 9600 15416 9628 15456
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 9968 15456 10241 15484
rect 9968 15428 9996 15456
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15453 13139 15487
rect 13081 15447 13139 15453
rect 7484 15388 9628 15416
rect 4154 15308 4160 15360
rect 4212 15348 4218 15360
rect 4617 15351 4675 15357
rect 4617 15348 4629 15351
rect 4212 15320 4629 15348
rect 4212 15308 4218 15320
rect 4617 15317 4629 15320
rect 4663 15317 4675 15351
rect 4617 15311 4675 15317
rect 5258 15308 5264 15360
rect 5316 15348 5322 15360
rect 7484 15348 7512 15388
rect 9950 15376 9956 15428
rect 10008 15376 10014 15428
rect 12526 15416 12532 15428
rect 10520 15388 12532 15416
rect 7650 15348 7656 15360
rect 5316 15320 7512 15348
rect 7611 15320 7656 15348
rect 5316 15308 5322 15320
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 7742 15308 7748 15360
rect 7800 15348 7806 15360
rect 9398 15348 9404 15360
rect 7800 15320 9404 15348
rect 7800 15308 7806 15320
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 9677 15351 9735 15357
rect 9677 15317 9689 15351
rect 9723 15348 9735 15351
rect 10520 15348 10548 15388
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 9723 15320 10548 15348
rect 9723 15317 9735 15320
rect 9677 15311 9735 15317
rect 10594 15308 10600 15360
rect 10652 15348 10658 15360
rect 13096 15348 13124 15447
rect 13170 15444 13176 15496
rect 13228 15484 13234 15496
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 13228 15456 13737 15484
rect 13228 15444 13234 15456
rect 13725 15453 13737 15456
rect 13771 15453 13783 15487
rect 13725 15447 13783 15453
rect 10652 15320 13124 15348
rect 10652 15308 10658 15320
rect 1104 15258 15824 15280
rect 1104 15206 3447 15258
rect 3499 15206 3511 15258
rect 3563 15206 3575 15258
rect 3627 15206 3639 15258
rect 3691 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 13308 15258
rect 13360 15206 13372 15258
rect 13424 15206 13436 15258
rect 13488 15206 13500 15258
rect 13552 15206 15824 15258
rect 1104 15184 15824 15206
rect 3697 15147 3755 15153
rect 3697 15113 3709 15147
rect 3743 15144 3755 15147
rect 4798 15144 4804 15156
rect 3743 15116 4804 15144
rect 3743 15113 3755 15116
rect 3697 15107 3755 15113
rect 4798 15104 4804 15116
rect 4856 15104 4862 15156
rect 5902 15104 5908 15156
rect 5960 15144 5966 15156
rect 8110 15144 8116 15156
rect 5960 15116 8116 15144
rect 5960 15104 5966 15116
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 8665 15147 8723 15153
rect 8665 15113 8677 15147
rect 8711 15144 8723 15147
rect 8938 15144 8944 15156
rect 8711 15116 8944 15144
rect 8711 15113 8723 15116
rect 8665 15107 8723 15113
rect 8938 15104 8944 15116
rect 8996 15104 9002 15156
rect 9398 15104 9404 15156
rect 9456 15144 9462 15156
rect 10502 15144 10508 15156
rect 9456 15116 10508 15144
rect 9456 15104 9462 15116
rect 10502 15104 10508 15116
rect 10560 15104 10566 15156
rect 12250 15104 12256 15156
rect 12308 15144 12314 15156
rect 12308 15116 12480 15144
rect 12308 15104 12314 15116
rect 7834 15036 7840 15088
rect 7892 15076 7898 15088
rect 11057 15079 11115 15085
rect 11057 15076 11069 15079
rect 7892 15048 11069 15076
rect 7892 15036 7898 15048
rect 11057 15045 11069 15048
rect 11103 15045 11115 15079
rect 11057 15039 11115 15045
rect 11164 15048 11652 15076
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 15008 2099 15011
rect 3234 15008 3240 15020
rect 2087 14980 3240 15008
rect 2087 14977 2099 14980
rect 2041 14971 2099 14977
rect 3234 14968 3240 14980
rect 3292 14968 3298 15020
rect 4154 15008 4160 15020
rect 4115 14980 4160 15008
rect 4154 14968 4160 14980
rect 4212 14968 4218 15020
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 15008 4399 15011
rect 4522 15008 4528 15020
rect 4387 14980 4528 15008
rect 4387 14977 4399 14980
rect 4341 14971 4399 14977
rect 4522 14968 4528 14980
rect 4580 14968 4586 15020
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 6825 15011 6883 15017
rect 6825 15008 6837 15011
rect 6788 14980 6837 15008
rect 6788 14968 6794 14980
rect 6825 14977 6837 14980
rect 6871 14977 6883 15011
rect 9214 15008 9220 15020
rect 9175 14980 9220 15008
rect 6825 14971 6883 14977
rect 9214 14968 9220 14980
rect 9272 14968 9278 15020
rect 9398 14968 9404 15020
rect 9456 15008 9462 15020
rect 10413 15011 10471 15017
rect 10413 15008 10425 15011
rect 9456 14980 10425 15008
rect 9456 14968 9462 14980
rect 10413 14977 10425 14980
rect 10459 14977 10471 15011
rect 10413 14971 10471 14977
rect 10502 14968 10508 15020
rect 10560 15008 10566 15020
rect 11164 15008 11192 15048
rect 10560 14980 11192 15008
rect 10560 14968 10566 14980
rect 11330 14968 11336 15020
rect 11388 15008 11394 15020
rect 11624 15017 11652 15048
rect 12452 15017 12480 15116
rect 11517 15011 11575 15017
rect 11517 15008 11529 15011
rect 11388 14980 11529 15008
rect 11388 14968 11394 14980
rect 11517 14977 11529 14980
rect 11563 14977 11575 15011
rect 11517 14971 11575 14977
rect 11609 15011 11667 15017
rect 11609 14977 11621 15011
rect 11655 14977 11667 15011
rect 11609 14971 11667 14977
rect 12437 15011 12495 15017
rect 12437 14977 12449 15011
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 1854 14900 1860 14952
rect 1912 14940 1918 14952
rect 2685 14943 2743 14949
rect 2685 14940 2697 14943
rect 1912 14912 2697 14940
rect 1912 14900 1918 14912
rect 2685 14909 2697 14912
rect 2731 14909 2743 14943
rect 2685 14903 2743 14909
rect 4798 14900 4804 14952
rect 4856 14940 4862 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4856 14912 4905 14940
rect 4856 14900 4862 14912
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 9033 14943 9091 14949
rect 4893 14903 4951 14909
rect 6840 14912 7236 14940
rect 2958 14872 2964 14884
rect 2919 14844 2964 14872
rect 2958 14832 2964 14844
rect 3016 14832 3022 14884
rect 4065 14875 4123 14881
rect 4065 14841 4077 14875
rect 4111 14872 4123 14875
rect 4338 14872 4344 14884
rect 4111 14844 4344 14872
rect 4111 14841 4123 14844
rect 4065 14835 4123 14841
rect 4338 14832 4344 14844
rect 4396 14832 4402 14884
rect 4706 14832 4712 14884
rect 4764 14872 4770 14884
rect 5160 14875 5218 14881
rect 5160 14872 5172 14875
rect 4764 14844 5172 14872
rect 4764 14832 4770 14844
rect 5160 14841 5172 14844
rect 5206 14872 5218 14875
rect 6840 14872 6868 14912
rect 5206 14844 6868 14872
rect 5206 14841 5218 14844
rect 5160 14835 5218 14841
rect 6914 14832 6920 14884
rect 6972 14872 6978 14884
rect 7070 14875 7128 14881
rect 7070 14872 7082 14875
rect 6972 14844 7082 14872
rect 6972 14832 6978 14844
rect 7070 14841 7082 14844
rect 7116 14841 7128 14875
rect 7208 14872 7236 14912
rect 9033 14909 9045 14943
rect 9079 14940 9091 14943
rect 11422 14940 11428 14952
rect 9079 14912 11428 14940
rect 9079 14909 9091 14912
rect 9033 14903 9091 14909
rect 11422 14900 11428 14912
rect 11480 14900 11486 14952
rect 7208 14844 8248 14872
rect 7070 14835 7128 14841
rect 5258 14764 5264 14816
rect 5316 14804 5322 14816
rect 6273 14807 6331 14813
rect 6273 14804 6285 14807
rect 5316 14776 6285 14804
rect 5316 14764 5322 14776
rect 6273 14773 6285 14776
rect 6319 14804 6331 14807
rect 7926 14804 7932 14816
rect 6319 14776 7932 14804
rect 6319 14773 6331 14776
rect 6273 14767 6331 14773
rect 7926 14764 7932 14776
rect 7984 14764 7990 14816
rect 8220 14813 8248 14844
rect 9674 14832 9680 14884
rect 9732 14872 9738 14884
rect 10321 14875 10379 14881
rect 10321 14872 10333 14875
rect 9732 14844 10333 14872
rect 9732 14832 9738 14844
rect 10321 14841 10333 14844
rect 10367 14841 10379 14875
rect 10778 14872 10784 14884
rect 10321 14835 10379 14841
rect 10520 14844 10784 14872
rect 10520 14816 10548 14844
rect 10778 14832 10784 14844
rect 10836 14832 10842 14884
rect 11698 14872 11704 14884
rect 11440 14844 11704 14872
rect 8205 14807 8263 14813
rect 8205 14773 8217 14807
rect 8251 14773 8263 14807
rect 8205 14767 8263 14773
rect 9125 14807 9183 14813
rect 9125 14773 9137 14807
rect 9171 14804 9183 14807
rect 9582 14804 9588 14816
rect 9171 14776 9588 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 9582 14764 9588 14776
rect 9640 14764 9646 14816
rect 9858 14804 9864 14816
rect 9819 14776 9864 14804
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 10229 14807 10287 14813
rect 10229 14773 10241 14807
rect 10275 14804 10287 14807
rect 10502 14804 10508 14816
rect 10275 14776 10508 14804
rect 10275 14773 10287 14776
rect 10229 14767 10287 14773
rect 10502 14764 10508 14776
rect 10560 14764 10566 14816
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 11440 14813 11468 14844
rect 11698 14832 11704 14844
rect 11756 14832 11762 14884
rect 12158 14832 12164 14884
rect 12216 14872 12222 14884
rect 14090 14872 14096 14884
rect 12216 14844 14096 14872
rect 12216 14832 12222 14844
rect 14090 14832 14096 14844
rect 14148 14832 14154 14884
rect 11425 14807 11483 14813
rect 11425 14804 11437 14807
rect 11204 14776 11437 14804
rect 11204 14764 11210 14776
rect 11425 14773 11437 14776
rect 11471 14773 11483 14807
rect 11425 14767 11483 14773
rect 11606 14764 11612 14816
rect 11664 14804 11670 14816
rect 12250 14804 12256 14816
rect 11664 14776 12256 14804
rect 11664 14764 11670 14776
rect 12250 14764 12256 14776
rect 12308 14764 12314 14816
rect 13078 14804 13084 14816
rect 13039 14776 13084 14804
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 13722 14804 13728 14816
rect 13683 14776 13728 14804
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 14366 14804 14372 14816
rect 14327 14776 14372 14804
rect 14366 14764 14372 14776
rect 14424 14764 14430 14816
rect 1104 14714 15824 14736
rect 1104 14662 5912 14714
rect 5964 14662 5976 14714
rect 6028 14662 6040 14714
rect 6092 14662 6104 14714
rect 6156 14662 10843 14714
rect 10895 14662 10907 14714
rect 10959 14662 10971 14714
rect 11023 14662 11035 14714
rect 11087 14662 15824 14714
rect 1104 14640 15824 14662
rect 2777 14603 2835 14609
rect 2777 14569 2789 14603
rect 2823 14600 2835 14603
rect 4246 14600 4252 14612
rect 2823 14572 4252 14600
rect 2823 14569 2835 14572
rect 2777 14563 2835 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 4430 14600 4436 14612
rect 4391 14572 4436 14600
rect 4430 14560 4436 14572
rect 4488 14560 4494 14612
rect 4890 14600 4896 14612
rect 4851 14572 4896 14600
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 7009 14603 7067 14609
rect 7009 14569 7021 14603
rect 7055 14600 7067 14603
rect 7466 14600 7472 14612
rect 7055 14572 7472 14600
rect 7055 14569 7067 14572
rect 7009 14563 7067 14569
rect 7466 14560 7472 14572
rect 7524 14560 7530 14612
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 9030 14600 9036 14612
rect 7616 14572 9036 14600
rect 7616 14560 7622 14572
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 9122 14560 9128 14612
rect 9180 14600 9186 14612
rect 9677 14603 9735 14609
rect 9677 14600 9689 14603
rect 9180 14572 9689 14600
rect 9180 14560 9186 14572
rect 9677 14569 9689 14572
rect 9723 14569 9735 14603
rect 9677 14563 9735 14569
rect 10134 14560 10140 14612
rect 10192 14600 10198 14612
rect 14090 14600 14096 14612
rect 10192 14572 13400 14600
rect 14051 14572 14096 14600
rect 10192 14560 10198 14572
rect 2133 14535 2191 14541
rect 2133 14501 2145 14535
rect 2179 14532 2191 14535
rect 2866 14532 2872 14544
rect 2179 14504 2872 14532
rect 2179 14501 2191 14504
rect 2133 14495 2191 14501
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 3237 14535 3295 14541
rect 3237 14501 3249 14535
rect 3283 14532 3295 14535
rect 3283 14504 5488 14532
rect 3283 14501 3295 14504
rect 3237 14495 3295 14501
rect 1857 14467 1915 14473
rect 1857 14433 1869 14467
rect 1903 14433 1915 14467
rect 1857 14427 1915 14433
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14433 3203 14467
rect 4798 14464 4804 14476
rect 4759 14436 4804 14464
rect 3145 14427 3203 14433
rect 1872 14328 1900 14427
rect 3050 14328 3056 14340
rect 1872 14300 3056 14328
rect 3050 14288 3056 14300
rect 3108 14288 3114 14340
rect 3160 14260 3188 14427
rect 4798 14424 4804 14436
rect 4856 14424 4862 14476
rect 5460 14464 5488 14504
rect 5534 14492 5540 14544
rect 5592 14532 5598 14544
rect 5874 14535 5932 14541
rect 5874 14532 5886 14535
rect 5592 14504 5886 14532
rect 5592 14492 5598 14504
rect 5874 14501 5886 14504
rect 5920 14532 5932 14535
rect 6270 14532 6276 14544
rect 5920 14504 6276 14532
rect 5920 14501 5932 14504
rect 5874 14495 5932 14501
rect 6270 14492 6276 14504
rect 6328 14492 6334 14544
rect 6822 14492 6828 14544
rect 6880 14532 6886 14544
rect 10778 14532 10784 14544
rect 6880 14504 10784 14532
rect 6880 14492 6886 14504
rect 10778 14492 10784 14504
rect 10836 14492 10842 14544
rect 11333 14535 11391 14541
rect 11333 14532 11345 14535
rect 10888 14504 11345 14532
rect 7558 14464 7564 14476
rect 5460 14436 7564 14464
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 7742 14473 7748 14476
rect 7736 14464 7748 14473
rect 7703 14436 7748 14464
rect 7736 14427 7748 14436
rect 7742 14424 7748 14427
rect 7800 14424 7806 14476
rect 8110 14424 8116 14476
rect 8168 14464 8174 14476
rect 8168 14436 8892 14464
rect 8168 14424 8174 14436
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 4522 14396 4528 14408
rect 3467 14368 4528 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 5077 14399 5135 14405
rect 4672 14368 5028 14396
rect 4672 14356 4678 14368
rect 4246 14288 4252 14340
rect 4304 14328 4310 14340
rect 4706 14328 4712 14340
rect 4304 14300 4712 14328
rect 4304 14288 4310 14300
rect 4706 14288 4712 14300
rect 4764 14288 4770 14340
rect 5000 14328 5028 14368
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5534 14396 5540 14408
rect 5123 14368 5540 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 5644 14328 5672 14359
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 7469 14399 7527 14405
rect 7469 14396 7481 14399
rect 7432 14368 7481 14396
rect 7432 14356 7438 14368
rect 7469 14365 7481 14368
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 8864 14337 8892 14436
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 9493 14467 9551 14473
rect 9493 14464 9505 14467
rect 9088 14436 9505 14464
rect 9088 14424 9094 14436
rect 9493 14433 9505 14436
rect 9539 14433 9551 14467
rect 9493 14427 9551 14433
rect 9582 14424 9588 14476
rect 9640 14464 9646 14476
rect 9766 14464 9772 14476
rect 9640 14436 9772 14464
rect 9640 14424 9646 14436
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 10042 14464 10048 14476
rect 10003 14436 10048 14464
rect 10042 14424 10048 14436
rect 10100 14464 10106 14476
rect 10888 14464 10916 14504
rect 11333 14501 11345 14504
rect 11379 14501 11391 14535
rect 11333 14495 11391 14501
rect 10100 14436 10916 14464
rect 10100 14424 10106 14436
rect 11146 14424 11152 14476
rect 11204 14464 11210 14476
rect 11241 14467 11299 14473
rect 11241 14464 11253 14467
rect 11204 14436 11253 14464
rect 11204 14424 11210 14436
rect 11241 14433 11253 14436
rect 11287 14433 11299 14467
rect 11241 14427 11299 14433
rect 11606 14424 11612 14476
rect 11664 14464 11670 14476
rect 13372 14473 13400 14572
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 12069 14467 12127 14473
rect 12069 14464 12081 14467
rect 11664 14436 12081 14464
rect 11664 14424 11670 14436
rect 12069 14433 12081 14436
rect 12115 14433 12127 14467
rect 12069 14427 12127 14433
rect 13357 14467 13415 14473
rect 13357 14433 13369 14467
rect 13403 14464 13415 14467
rect 13630 14464 13636 14476
rect 13403 14436 13636 14464
rect 13403 14433 13415 14436
rect 13357 14427 13415 14433
rect 13630 14424 13636 14436
rect 13688 14424 13694 14476
rect 8938 14356 8944 14408
rect 8996 14396 9002 14408
rect 9858 14396 9864 14408
rect 8996 14368 9864 14396
rect 8996 14356 9002 14368
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 10134 14396 10140 14408
rect 10095 14368 10140 14396
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 5000 14300 5672 14328
rect 8849 14331 8907 14337
rect 8849 14297 8861 14331
rect 8895 14297 8907 14331
rect 9214 14328 9220 14340
rect 8849 14291 8907 14297
rect 8956 14300 9220 14328
rect 8956 14272 8984 14300
rect 9214 14288 9220 14300
rect 9272 14328 9278 14340
rect 10244 14328 10272 14359
rect 10410 14356 10416 14408
rect 10468 14396 10474 14408
rect 11054 14396 11060 14408
rect 10468 14368 11060 14396
rect 10468 14356 10474 14368
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 11422 14396 11428 14408
rect 11383 14368 11428 14396
rect 11422 14356 11428 14368
rect 11480 14356 11486 14408
rect 12253 14399 12311 14405
rect 12253 14365 12265 14399
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 9272 14300 10272 14328
rect 9272 14288 9278 14300
rect 10778 14288 10784 14340
rect 10836 14328 10842 14340
rect 10873 14331 10931 14337
rect 10873 14328 10885 14331
rect 10836 14300 10885 14328
rect 10836 14288 10842 14300
rect 10873 14297 10885 14300
rect 10919 14297 10931 14331
rect 10873 14291 10931 14297
rect 11330 14288 11336 14340
rect 11388 14328 11394 14340
rect 12268 14328 12296 14359
rect 11388 14300 12296 14328
rect 11388 14288 11394 14300
rect 8110 14260 8116 14272
rect 3160 14232 8116 14260
rect 8110 14220 8116 14232
rect 8168 14220 8174 14272
rect 8938 14220 8944 14272
rect 8996 14220 9002 14272
rect 9122 14220 9128 14272
rect 9180 14260 9186 14272
rect 9309 14263 9367 14269
rect 9309 14260 9321 14263
rect 9180 14232 9321 14260
rect 9180 14220 9186 14232
rect 9309 14229 9321 14232
rect 9355 14229 9367 14263
rect 9309 14223 9367 14229
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 11698 14260 11704 14272
rect 9916 14232 11704 14260
rect 9916 14220 9922 14232
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 13541 14263 13599 14269
rect 13541 14229 13553 14263
rect 13587 14260 13599 14263
rect 15470 14260 15476 14272
rect 13587 14232 15476 14260
rect 13587 14229 13599 14232
rect 13541 14223 13599 14229
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 1104 14170 15824 14192
rect 1104 14118 3447 14170
rect 3499 14118 3511 14170
rect 3563 14118 3575 14170
rect 3627 14118 3639 14170
rect 3691 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 13308 14170
rect 13360 14118 13372 14170
rect 13424 14118 13436 14170
rect 13488 14118 13500 14170
rect 13552 14118 15824 14170
rect 1104 14096 15824 14118
rect 3697 14059 3755 14065
rect 3697 14025 3709 14059
rect 3743 14056 3755 14059
rect 4798 14056 4804 14068
rect 3743 14028 4804 14056
rect 3743 14025 3755 14028
rect 3697 14019 3755 14025
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 8018 14056 8024 14068
rect 4915 14028 8024 14056
rect 2501 13991 2559 13997
rect 2501 13957 2513 13991
rect 2547 13988 2559 13991
rect 3970 13988 3976 14000
rect 2547 13960 3976 13988
rect 2547 13957 2559 13960
rect 2501 13951 2559 13957
rect 3970 13948 3976 13960
rect 4028 13948 4034 14000
rect 4915 13988 4943 14028
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 8110 14016 8116 14068
rect 8168 14056 8174 14068
rect 8168 14028 9628 14056
rect 8168 14016 8174 14028
rect 6270 13988 6276 14000
rect 4172 13960 4943 13988
rect 6231 13960 6276 13988
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 1765 13923 1823 13929
rect 1765 13920 1777 13923
rect 1452 13892 1777 13920
rect 1452 13880 1458 13892
rect 1765 13889 1777 13892
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 4062 13920 4068 13932
rect 3191 13892 4068 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4172 13929 4200 13960
rect 6270 13948 6276 13960
rect 6328 13948 6334 14000
rect 7834 13948 7840 14000
rect 7892 13988 7898 14000
rect 8205 13991 8263 13997
rect 8205 13988 8217 13991
rect 7892 13960 8217 13988
rect 7892 13948 7898 13960
rect 8205 13957 8217 13960
rect 8251 13957 8263 13991
rect 9600 13988 9628 14028
rect 10134 14016 10140 14068
rect 10192 14056 10198 14068
rect 10505 14059 10563 14065
rect 10505 14056 10517 14059
rect 10192 14028 10517 14056
rect 10192 14016 10198 14028
rect 10505 14025 10517 14028
rect 10551 14025 10563 14059
rect 10505 14019 10563 14025
rect 12802 14016 12808 14068
rect 12860 14056 12866 14068
rect 12860 14028 13492 14056
rect 12860 14016 12866 14028
rect 13464 14000 13492 14028
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 14182 14056 14188 14068
rect 13872 14028 14188 14056
rect 13872 14016 13878 14028
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 12437 13991 12495 13997
rect 12437 13988 12449 13991
rect 9600 13960 12449 13988
rect 8205 13951 8263 13957
rect 12437 13957 12449 13960
rect 12483 13957 12495 13991
rect 12437 13951 12495 13957
rect 13446 13948 13452 14000
rect 13504 13948 13510 14000
rect 14001 13991 14059 13997
rect 14001 13957 14013 13991
rect 14047 13988 14059 13991
rect 14918 13988 14924 14000
rect 14047 13960 14924 13988
rect 14047 13957 14059 13960
rect 14001 13951 14059 13957
rect 14918 13948 14924 13960
rect 14976 13948 14982 14000
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13889 4215 13923
rect 4157 13883 4215 13889
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4387 13892 4476 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13852 3019 13855
rect 3326 13852 3332 13864
rect 3007 13824 3332 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 4448 13796 4476 13892
rect 7926 13880 7932 13932
rect 7984 13920 7990 13932
rect 11057 13923 11115 13929
rect 11057 13920 11069 13923
rect 7984 13892 8800 13920
rect 7984 13880 7990 13892
rect 4614 13812 4620 13864
rect 4672 13852 4678 13864
rect 4893 13855 4951 13861
rect 4893 13852 4905 13855
rect 4672 13824 4905 13852
rect 4672 13812 4678 13824
rect 4893 13821 4905 13824
rect 4939 13821 4951 13855
rect 4893 13815 4951 13821
rect 6730 13812 6736 13864
rect 6788 13852 6794 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6788 13824 6837 13852
rect 6788 13812 6794 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 7092 13855 7150 13861
rect 7092 13821 7104 13855
rect 7138 13852 7150 13855
rect 7466 13852 7472 13864
rect 7138 13824 7472 13852
rect 7138 13821 7150 13824
rect 7092 13815 7150 13821
rect 4430 13744 4436 13796
rect 4488 13744 4494 13796
rect 4522 13744 4528 13796
rect 4580 13784 4586 13796
rect 5160 13787 5218 13793
rect 5160 13784 5172 13787
rect 4580 13756 5172 13784
rect 4580 13744 4586 13756
rect 5160 13753 5172 13756
rect 5206 13784 5218 13787
rect 5442 13784 5448 13796
rect 5206 13756 5448 13784
rect 5206 13753 5218 13756
rect 5160 13747 5218 13753
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 6840 13784 6868 13815
rect 7466 13812 7472 13824
rect 7524 13812 7530 13864
rect 8662 13852 8668 13864
rect 7576 13824 8668 13852
rect 7374 13784 7380 13796
rect 6840 13756 7380 13784
rect 7374 13744 7380 13756
rect 7432 13784 7438 13796
rect 7576 13784 7604 13824
rect 8662 13812 8668 13824
rect 8720 13812 8726 13864
rect 8772 13852 8800 13892
rect 9692 13892 11069 13920
rect 8921 13855 8979 13861
rect 8921 13852 8933 13855
rect 8772 13824 8933 13852
rect 8921 13821 8933 13824
rect 8967 13821 8979 13855
rect 8921 13815 8979 13821
rect 7432 13756 7604 13784
rect 7432 13744 7438 13756
rect 8110 13744 8116 13796
rect 8168 13784 8174 13796
rect 9692 13784 9720 13892
rect 11057 13889 11069 13892
rect 11103 13889 11115 13923
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 11057 13883 11115 13889
rect 11624 13892 13001 13920
rect 9858 13812 9864 13864
rect 9916 13852 9922 13864
rect 10226 13852 10232 13864
rect 9916 13824 10232 13852
rect 9916 13812 9922 13824
rect 10226 13812 10232 13824
rect 10284 13852 10290 13864
rect 10965 13855 11023 13861
rect 10965 13852 10977 13855
rect 10284 13824 10977 13852
rect 10284 13812 10290 13824
rect 10965 13821 10977 13824
rect 11011 13821 11023 13855
rect 10965 13815 11023 13821
rect 8168 13756 9720 13784
rect 8168 13744 8174 13756
rect 10134 13744 10140 13796
rect 10192 13784 10198 13796
rect 10410 13784 10416 13796
rect 10192 13756 10416 13784
rect 10192 13744 10198 13756
rect 10410 13744 10416 13756
rect 10468 13744 10474 13796
rect 10502 13744 10508 13796
rect 10560 13784 10566 13796
rect 10686 13784 10692 13796
rect 10560 13756 10692 13784
rect 10560 13744 10566 13756
rect 10686 13744 10692 13756
rect 10744 13784 10750 13796
rect 10873 13787 10931 13793
rect 10873 13784 10885 13787
rect 10744 13756 10885 13784
rect 10744 13744 10750 13756
rect 10873 13753 10885 13756
rect 10919 13753 10931 13787
rect 10873 13747 10931 13753
rect 11624 13728 11652 13892
rect 12989 13889 13001 13892
rect 13035 13920 13047 13923
rect 13538 13920 13544 13932
rect 13035 13892 13544 13920
rect 13035 13889 13047 13892
rect 12989 13883 13047 13889
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 13262 13852 13268 13864
rect 12584 13824 13268 13852
rect 12584 13812 12590 13824
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13814 13852 13820 13864
rect 13775 13824 13820 13852
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 11701 13787 11759 13793
rect 11701 13753 11713 13787
rect 11747 13784 11759 13787
rect 12805 13787 12863 13793
rect 12805 13784 12817 13787
rect 11747 13756 12817 13784
rect 11747 13753 11759 13756
rect 11701 13747 11759 13753
rect 12805 13753 12817 13756
rect 12851 13753 12863 13787
rect 14550 13784 14556 13796
rect 14511 13756 14556 13784
rect 12805 13747 12863 13753
rect 14550 13744 14556 13756
rect 14608 13744 14614 13796
rect 2869 13719 2927 13725
rect 2869 13685 2881 13719
rect 2915 13716 2927 13719
rect 3142 13716 3148 13728
rect 2915 13688 3148 13716
rect 2915 13685 2927 13688
rect 2869 13679 2927 13685
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 4065 13719 4123 13725
rect 4065 13685 4077 13719
rect 4111 13716 4123 13719
rect 7650 13716 7656 13728
rect 4111 13688 7656 13716
rect 4111 13685 4123 13688
rect 4065 13679 4123 13685
rect 7650 13676 7656 13688
rect 7708 13676 7714 13728
rect 8662 13676 8668 13728
rect 8720 13716 8726 13728
rect 9306 13716 9312 13728
rect 8720 13688 9312 13716
rect 8720 13676 8726 13688
rect 9306 13676 9312 13688
rect 9364 13676 9370 13728
rect 9950 13676 9956 13728
rect 10008 13716 10014 13728
rect 10045 13719 10103 13725
rect 10045 13716 10057 13719
rect 10008 13688 10057 13716
rect 10008 13676 10014 13688
rect 10045 13685 10057 13688
rect 10091 13716 10103 13719
rect 11422 13716 11428 13728
rect 10091 13688 11428 13716
rect 10091 13685 10103 13688
rect 10045 13679 10103 13685
rect 11422 13676 11428 13688
rect 11480 13676 11486 13728
rect 11606 13676 11612 13728
rect 11664 13676 11670 13728
rect 12897 13719 12955 13725
rect 12897 13685 12909 13719
rect 12943 13716 12955 13719
rect 14090 13716 14096 13728
rect 12943 13688 14096 13716
rect 12943 13685 12955 13688
rect 12897 13679 12955 13685
rect 14090 13676 14096 13688
rect 14148 13716 14154 13728
rect 15746 13716 15752 13728
rect 14148 13688 15752 13716
rect 14148 13676 14154 13688
rect 15746 13676 15752 13688
rect 15804 13676 15810 13728
rect 1104 13626 15824 13648
rect 1104 13574 5912 13626
rect 5964 13574 5976 13626
rect 6028 13574 6040 13626
rect 6092 13574 6104 13626
rect 6156 13574 10843 13626
rect 10895 13574 10907 13626
rect 10959 13574 10971 13626
rect 11023 13574 11035 13626
rect 11087 13574 15824 13626
rect 1104 13552 15824 13574
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 4338 13512 4344 13524
rect 1995 13484 4344 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 4338 13472 4344 13484
rect 4396 13472 4402 13524
rect 4430 13472 4436 13524
rect 4488 13512 4494 13524
rect 5166 13512 5172 13524
rect 4488 13484 5172 13512
rect 4488 13472 4494 13484
rect 5166 13472 5172 13484
rect 5224 13472 5230 13524
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 8018 13512 8024 13524
rect 7979 13484 8024 13512
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 9398 13512 9404 13524
rect 8352 13484 9404 13512
rect 8352 13472 8358 13484
rect 9398 13472 9404 13484
rect 9456 13472 9462 13524
rect 9766 13472 9772 13524
rect 9824 13512 9830 13524
rect 11517 13515 11575 13521
rect 11517 13512 11529 13515
rect 9824 13484 11529 13512
rect 9824 13472 9830 13484
rect 11517 13481 11529 13484
rect 11563 13481 11575 13515
rect 11517 13475 11575 13481
rect 11885 13515 11943 13521
rect 11885 13481 11897 13515
rect 11931 13512 11943 13515
rect 13078 13512 13084 13524
rect 11931 13484 13084 13512
rect 11931 13481 11943 13484
rect 11885 13475 11943 13481
rect 13078 13472 13084 13484
rect 13136 13472 13142 13524
rect 13173 13515 13231 13521
rect 13173 13481 13185 13515
rect 13219 13512 13231 13515
rect 13262 13512 13268 13524
rect 13219 13484 13268 13512
rect 13219 13481 13231 13484
rect 13173 13475 13231 13481
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 3145 13447 3203 13453
rect 3145 13413 3157 13447
rect 3191 13444 3203 13447
rect 3326 13444 3332 13456
rect 3191 13416 3332 13444
rect 3191 13413 3203 13416
rect 3145 13407 3203 13413
rect 3326 13404 3332 13416
rect 3384 13404 3390 13456
rect 5258 13444 5264 13456
rect 3436 13416 5264 13444
rect 2240 13348 3372 13376
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13308 2099 13311
rect 2130 13308 2136 13320
rect 2087 13280 2136 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 2130 13268 2136 13280
rect 2188 13268 2194 13320
rect 2240 13317 2268 13348
rect 2225 13311 2283 13317
rect 2225 13277 2237 13311
rect 2271 13277 2283 13311
rect 2225 13271 2283 13277
rect 2774 13268 2780 13320
rect 2832 13308 2838 13320
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 2832 13280 3249 13308
rect 2832 13268 2838 13280
rect 3237 13277 3249 13280
rect 3283 13277 3295 13311
rect 3237 13271 3295 13277
rect 1581 13243 1639 13249
rect 1581 13209 1593 13243
rect 1627 13240 1639 13243
rect 2590 13240 2596 13252
rect 1627 13212 2596 13240
rect 1627 13209 1639 13212
rect 1581 13203 1639 13209
rect 2590 13200 2596 13212
rect 2648 13200 2654 13252
rect 2777 13175 2835 13181
rect 2777 13141 2789 13175
rect 2823 13172 2835 13175
rect 2866 13172 2872 13184
rect 2823 13144 2872 13172
rect 2823 13141 2835 13144
rect 2777 13135 2835 13141
rect 2866 13132 2872 13144
rect 2924 13132 2930 13184
rect 3344 13172 3372 13348
rect 3436 13317 3464 13416
rect 5258 13404 5264 13416
rect 5316 13404 5322 13456
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 6270 13444 6276 13456
rect 5592 13416 6276 13444
rect 5592 13404 5598 13416
rect 6270 13404 6276 13416
rect 6328 13444 6334 13456
rect 6426 13447 6484 13453
rect 6426 13444 6438 13447
rect 6328 13416 6438 13444
rect 6328 13404 6334 13416
rect 6426 13413 6438 13416
rect 6472 13413 6484 13447
rect 6426 13407 6484 13413
rect 7466 13404 7472 13456
rect 7524 13444 7530 13456
rect 7524 13416 9536 13444
rect 7524 13404 7530 13416
rect 4341 13379 4399 13385
rect 4341 13345 4353 13379
rect 4387 13376 4399 13379
rect 4430 13376 4436 13388
rect 4387 13348 4436 13376
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 4430 13336 4436 13348
rect 4488 13336 4494 13388
rect 4608 13379 4666 13385
rect 4608 13345 4620 13379
rect 4654 13376 4666 13379
rect 5810 13376 5816 13388
rect 4654 13348 5816 13376
rect 4654 13345 4666 13348
rect 4608 13339 4666 13345
rect 5810 13336 5816 13348
rect 5868 13336 5874 13388
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13376 6239 13379
rect 6730 13376 6736 13388
rect 6227 13348 6736 13376
rect 6227 13345 6239 13348
rect 6181 13339 6239 13345
rect 6730 13336 6736 13348
rect 6788 13336 6794 13388
rect 6822 13336 6828 13388
rect 6880 13376 6886 13388
rect 8294 13376 8300 13388
rect 6880 13348 8300 13376
rect 6880 13336 6886 13348
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 8386 13336 8392 13388
rect 8444 13376 8450 13388
rect 9398 13376 9404 13388
rect 8444 13348 8489 13376
rect 9359 13348 9404 13376
rect 8444 13336 8450 13348
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 9508 13376 9536 13416
rect 9674 13404 9680 13456
rect 9732 13444 9738 13456
rect 11054 13444 11060 13456
rect 9732 13416 11060 13444
rect 9732 13404 9738 13416
rect 11054 13404 11060 13416
rect 11112 13404 11118 13456
rect 11977 13447 12035 13453
rect 11977 13413 11989 13447
rect 12023 13444 12035 13447
rect 12023 13416 12296 13444
rect 12023 13413 12035 13416
rect 11977 13407 12035 13413
rect 9950 13385 9956 13388
rect 9944 13376 9956 13385
rect 9508 13348 9956 13376
rect 9944 13339 9956 13348
rect 9950 13336 9956 13339
rect 10008 13336 10014 13388
rect 10410 13336 10416 13388
rect 10468 13376 10474 13388
rect 12268 13376 12296 13416
rect 12526 13376 12532 13388
rect 10468 13348 11008 13376
rect 12268 13348 12532 13376
rect 10468 13336 10474 13348
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13277 8539 13311
rect 8481 13271 8539 13277
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 8938 13308 8944 13320
rect 8711 13280 8944 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 8496 13240 8524 13271
rect 8938 13268 8944 13280
rect 8996 13268 9002 13320
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13308 9551 13311
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9539 13280 9689 13308
rect 9539 13277 9551 13280
rect 9493 13271 9551 13277
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 10980 13240 11008 13348
rect 12526 13336 12532 13348
rect 12584 13336 12590 13388
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 12802 13376 12808 13388
rect 12676 13348 12808 13376
rect 12676 13336 12682 13348
rect 12802 13336 12808 13348
rect 12860 13376 12866 13388
rect 13081 13379 13139 13385
rect 13081 13376 13093 13379
rect 12860 13348 13093 13376
rect 12860 13336 12866 13348
rect 13081 13345 13093 13348
rect 13127 13345 13139 13379
rect 13906 13376 13912 13388
rect 13867 13348 13912 13376
rect 13081 13339 13139 13345
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 11388 13280 12173 13308
rect 11388 13268 11394 13280
rect 12161 13277 12173 13280
rect 12207 13308 12219 13311
rect 13357 13311 13415 13317
rect 12207 13280 12848 13308
rect 12207 13277 12219 13280
rect 12161 13271 12219 13277
rect 12820 13252 12848 13280
rect 13357 13277 13369 13311
rect 13403 13308 13415 13311
rect 13538 13308 13544 13320
rect 13403 13280 13544 13308
rect 13403 13277 13415 13280
rect 13357 13271 13415 13277
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 13722 13268 13728 13320
rect 13780 13308 13786 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 13780 13280 14105 13308
rect 13780 13268 13786 13280
rect 14093 13277 14105 13280
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 11057 13243 11115 13249
rect 11057 13240 11069 13243
rect 8496 13212 9720 13240
rect 10980 13212 11069 13240
rect 7466 13172 7472 13184
rect 3344 13144 7472 13172
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 7561 13175 7619 13181
rect 7561 13141 7573 13175
rect 7607 13172 7619 13175
rect 7650 13172 7656 13184
rect 7607 13144 7656 13172
rect 7607 13141 7619 13144
rect 7561 13135 7619 13141
rect 7650 13132 7656 13144
rect 7708 13132 7714 13184
rect 9214 13172 9220 13184
rect 9175 13144 9220 13172
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 9306 13132 9312 13184
rect 9364 13172 9370 13184
rect 9493 13175 9551 13181
rect 9493 13172 9505 13175
rect 9364 13144 9505 13172
rect 9364 13132 9370 13144
rect 9493 13141 9505 13144
rect 9539 13141 9551 13175
rect 9692 13172 9720 13212
rect 11057 13209 11069 13212
rect 11103 13240 11115 13243
rect 11606 13240 11612 13252
rect 11103 13212 11612 13240
rect 11103 13209 11115 13212
rect 11057 13203 11115 13209
rect 11606 13200 11612 13212
rect 11664 13200 11670 13252
rect 11698 13200 11704 13252
rect 11756 13240 11762 13252
rect 12713 13243 12771 13249
rect 12713 13240 12725 13243
rect 11756 13212 12725 13240
rect 11756 13200 11762 13212
rect 12713 13209 12725 13212
rect 12759 13209 12771 13243
rect 12713 13203 12771 13209
rect 12802 13200 12808 13252
rect 12860 13200 12866 13252
rect 13906 13200 13912 13252
rect 13964 13240 13970 13252
rect 14274 13240 14280 13252
rect 13964 13212 14280 13240
rect 13964 13200 13970 13212
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 14182 13172 14188 13184
rect 9692 13144 14188 13172
rect 9493 13135 9551 13141
rect 14182 13132 14188 13144
rect 14240 13172 14246 13184
rect 15102 13172 15108 13184
rect 14240 13144 15108 13172
rect 14240 13132 14246 13144
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 1104 13082 15824 13104
rect 1104 13030 3447 13082
rect 3499 13030 3511 13082
rect 3563 13030 3575 13082
rect 3627 13030 3639 13082
rect 3691 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 13308 13082
rect 13360 13030 13372 13082
rect 13424 13030 13436 13082
rect 13488 13030 13500 13082
rect 13552 13030 15824 13082
rect 1104 13008 15824 13030
rect 3050 12928 3056 12980
rect 3108 12968 3114 12980
rect 6270 12968 6276 12980
rect 3108 12940 6132 12968
rect 6231 12940 6276 12968
rect 3108 12928 3114 12940
rect 1857 12903 1915 12909
rect 1857 12869 1869 12903
rect 1903 12900 1915 12903
rect 2406 12900 2412 12912
rect 1903 12872 2412 12900
rect 1903 12869 1915 12872
rect 1857 12863 1915 12869
rect 2406 12860 2412 12872
rect 2464 12860 2470 12912
rect 4433 12903 4491 12909
rect 4433 12869 4445 12903
rect 4479 12869 4491 12903
rect 6104 12900 6132 12940
rect 6270 12928 6276 12940
rect 6328 12928 6334 12980
rect 8205 12971 8263 12977
rect 6748 12940 8156 12968
rect 6748 12900 6776 12940
rect 6104 12872 6776 12900
rect 4433 12863 4491 12869
rect 2498 12832 2504 12844
rect 2459 12804 2504 12832
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 4448 12832 4476 12863
rect 6822 12860 6828 12912
rect 6880 12860 6886 12912
rect 8128 12900 8156 12940
rect 8205 12937 8217 12971
rect 8251 12968 8263 12971
rect 8938 12968 8944 12980
rect 8251 12940 8944 12968
rect 8251 12937 8263 12940
rect 8205 12931 8263 12937
rect 8938 12928 8944 12940
rect 8996 12928 9002 12980
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 9364 12940 9628 12968
rect 9364 12928 9370 12940
rect 8478 12900 8484 12912
rect 8128 12872 8484 12900
rect 8478 12860 8484 12872
rect 8536 12860 8542 12912
rect 9600 12900 9628 12940
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 13633 12971 13691 12977
rect 13633 12968 13645 12971
rect 9732 12940 13645 12968
rect 9732 12928 9738 12940
rect 13633 12937 13645 12940
rect 13679 12937 13691 12971
rect 13633 12931 13691 12937
rect 9950 12900 9956 12912
rect 9600 12872 9956 12900
rect 9950 12860 9956 12872
rect 10008 12860 10014 12912
rect 10226 12860 10232 12912
rect 10284 12900 10290 12912
rect 10505 12903 10563 12909
rect 10505 12900 10517 12903
rect 10284 12872 10517 12900
rect 10284 12860 10290 12872
rect 10505 12869 10517 12872
rect 10551 12869 10563 12903
rect 10505 12863 10563 12869
rect 11422 12860 11428 12912
rect 11480 12900 11486 12912
rect 12437 12903 12495 12909
rect 12437 12900 12449 12903
rect 11480 12872 12449 12900
rect 11480 12860 11486 12872
rect 12437 12869 12449 12872
rect 12483 12869 12495 12903
rect 12437 12863 12495 12869
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 14274 12900 14280 12912
rect 12584 12872 14280 12900
rect 12584 12860 12590 12872
rect 14274 12860 14280 12872
rect 14332 12900 14338 12912
rect 15378 12900 15384 12912
rect 14332 12872 15384 12900
rect 14332 12860 14338 12872
rect 15378 12860 15384 12872
rect 15436 12860 15442 12912
rect 6840 12832 6868 12860
rect 4448 12804 5028 12832
rect 2225 12767 2283 12773
rect 2225 12733 2237 12767
rect 2271 12764 2283 12767
rect 2590 12764 2596 12776
rect 2271 12736 2596 12764
rect 2271 12733 2283 12736
rect 2225 12727 2283 12733
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 3053 12767 3111 12773
rect 3053 12733 3065 12767
rect 3099 12764 3111 12767
rect 4614 12764 4620 12776
rect 3099 12736 4620 12764
rect 3099 12733 3111 12736
rect 3053 12727 3111 12733
rect 4614 12724 4620 12736
rect 4672 12764 4678 12776
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 4672 12736 4905 12764
rect 4672 12724 4678 12736
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 4893 12727 4951 12733
rect 3320 12699 3378 12705
rect 3320 12665 3332 12699
rect 3366 12696 3378 12699
rect 3510 12696 3516 12708
rect 3366 12668 3516 12696
rect 3366 12665 3378 12668
rect 3320 12659 3378 12665
rect 3510 12656 3516 12668
rect 3568 12656 3574 12708
rect 5000 12696 5028 12804
rect 5920 12804 6868 12832
rect 5166 12773 5172 12776
rect 5160 12764 5172 12773
rect 5127 12736 5172 12764
rect 5160 12727 5172 12736
rect 5166 12724 5172 12727
rect 5224 12724 5230 12776
rect 5920 12764 5948 12804
rect 7834 12792 7840 12844
rect 7892 12832 7898 12844
rect 8662 12832 8668 12844
rect 7892 12804 8524 12832
rect 8623 12804 8668 12832
rect 7892 12792 7898 12804
rect 5276 12736 5948 12764
rect 6825 12767 6883 12773
rect 5276 12708 5304 12736
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 6825 12727 6883 12733
rect 5258 12696 5264 12708
rect 4356 12668 4660 12696
rect 5000 12668 5264 12696
rect 2317 12631 2375 12637
rect 2317 12597 2329 12631
rect 2363 12628 2375 12631
rect 4356 12628 4384 12668
rect 2363 12600 4384 12628
rect 4632 12628 4660 12668
rect 5258 12656 5264 12668
rect 5316 12656 5322 12708
rect 5534 12656 5540 12708
rect 5592 12696 5598 12708
rect 6840 12696 6868 12727
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 7092 12767 7150 12773
rect 7092 12764 7104 12767
rect 6972 12736 7104 12764
rect 6972 12724 6978 12736
rect 7092 12733 7104 12736
rect 7138 12764 7150 12767
rect 8110 12764 8116 12776
rect 7138 12736 8116 12764
rect 7138 12733 7150 12736
rect 7092 12727 7150 12733
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 8496 12764 8524 12804
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 10686 12792 10692 12844
rect 10744 12832 10750 12844
rect 11057 12835 11115 12841
rect 11057 12832 11069 12835
rect 10744 12804 11069 12832
rect 10744 12792 10750 12804
rect 11057 12801 11069 12804
rect 11103 12801 11115 12835
rect 11057 12795 11115 12801
rect 12802 12792 12808 12844
rect 12860 12832 12866 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12860 12804 13001 12832
rect 12860 12792 12866 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13630 12792 13636 12844
rect 13688 12832 13694 12844
rect 13688 12804 13952 12832
rect 13688 12792 13694 12804
rect 9214 12764 9220 12776
rect 8496 12736 9220 12764
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 9306 12724 9312 12776
rect 9364 12764 9370 12776
rect 10873 12767 10931 12773
rect 10873 12764 10885 12767
rect 9364 12736 10885 12764
rect 9364 12724 9370 12736
rect 10873 12733 10885 12736
rect 10919 12733 10931 12767
rect 10873 12727 10931 12733
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 13924 12773 13952 12804
rect 14182 12792 14188 12844
rect 14240 12832 14246 12844
rect 15010 12832 15016 12844
rect 14240 12804 15016 12832
rect 14240 12792 14246 12804
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 13817 12767 13875 12773
rect 13817 12764 13829 12767
rect 11204 12736 13829 12764
rect 11204 12724 11210 12736
rect 13817 12733 13829 12736
rect 13863 12733 13875 12767
rect 13817 12727 13875 12733
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12733 13967 12767
rect 14826 12764 14832 12776
rect 14787 12736 14832 12764
rect 13909 12727 13967 12733
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 7374 12696 7380 12708
rect 5592 12668 7380 12696
rect 5592 12656 5598 12668
rect 7374 12656 7380 12668
rect 7432 12696 7438 12708
rect 7432 12668 7687 12696
rect 7432 12656 7438 12668
rect 7558 12628 7564 12640
rect 4632 12600 7564 12628
rect 2363 12597 2375 12600
rect 2317 12591 2375 12597
rect 7558 12588 7564 12600
rect 7616 12588 7622 12640
rect 7659 12628 7687 12668
rect 8202 12656 8208 12708
rect 8260 12696 8266 12708
rect 8910 12699 8968 12705
rect 8910 12696 8922 12699
rect 8260 12668 8922 12696
rect 8260 12656 8266 12668
rect 8910 12665 8922 12668
rect 8956 12665 8968 12699
rect 8910 12659 8968 12665
rect 9766 12656 9772 12708
rect 9824 12696 9830 12708
rect 10965 12699 11023 12705
rect 10965 12696 10977 12699
rect 9824 12668 10977 12696
rect 9824 12656 9830 12668
rect 10965 12665 10977 12668
rect 11011 12665 11023 12699
rect 11330 12696 11336 12708
rect 10965 12659 11023 12665
rect 11072 12668 11336 12696
rect 9582 12628 9588 12640
rect 7659 12600 9588 12628
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10045 12631 10103 12637
rect 10045 12628 10057 12631
rect 10008 12600 10057 12628
rect 10008 12588 10014 12600
rect 10045 12597 10057 12600
rect 10091 12628 10103 12631
rect 11072 12628 11100 12668
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 14185 12699 14243 12705
rect 14185 12665 14197 12699
rect 14231 12696 14243 12699
rect 15746 12696 15752 12708
rect 14231 12668 15752 12696
rect 14231 12665 14243 12668
rect 14185 12659 14243 12665
rect 15746 12656 15752 12668
rect 15804 12656 15810 12708
rect 11698 12628 11704 12640
rect 10091 12600 11100 12628
rect 11659 12600 11704 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 12066 12588 12072 12640
rect 12124 12628 12130 12640
rect 12250 12628 12256 12640
rect 12124 12600 12256 12628
rect 12124 12588 12130 12600
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 12802 12628 12808 12640
rect 12763 12600 12808 12628
rect 12802 12588 12808 12600
rect 12860 12588 12866 12640
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13998 12628 14004 12640
rect 12943 12600 14004 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13998 12588 14004 12600
rect 14056 12628 14062 12640
rect 14826 12628 14832 12640
rect 14056 12600 14832 12628
rect 14056 12588 14062 12600
rect 14826 12588 14832 12600
rect 14884 12588 14890 12640
rect 15010 12628 15016 12640
rect 14971 12600 15016 12628
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 1104 12538 15824 12560
rect 1104 12486 5912 12538
rect 5964 12486 5976 12538
rect 6028 12486 6040 12538
rect 6092 12486 6104 12538
rect 6156 12486 10843 12538
rect 10895 12486 10907 12538
rect 10959 12486 10971 12538
rect 11023 12486 11035 12538
rect 11087 12486 15824 12538
rect 1104 12464 15824 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 2832 12396 2877 12424
rect 2832 12384 2838 12396
rect 3050 12384 3056 12436
rect 3108 12424 3114 12436
rect 3145 12427 3203 12433
rect 3145 12424 3157 12427
rect 3108 12396 3157 12424
rect 3108 12384 3114 12396
rect 3145 12393 3157 12396
rect 3191 12393 3203 12427
rect 3145 12387 3203 12393
rect 3237 12427 3295 12433
rect 3237 12393 3249 12427
rect 3283 12424 3295 12427
rect 6638 12424 6644 12436
rect 3283 12396 6644 12424
rect 3283 12393 3295 12396
rect 3237 12387 3295 12393
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 6914 12424 6920 12436
rect 6875 12396 6920 12424
rect 6914 12384 6920 12396
rect 6972 12384 6978 12436
rect 9217 12427 9275 12433
rect 7024 12396 7972 12424
rect 2041 12359 2099 12365
rect 2041 12325 2053 12359
rect 2087 12356 2099 12359
rect 2590 12356 2596 12368
rect 2087 12328 2596 12356
rect 2087 12325 2099 12328
rect 2041 12319 2099 12325
rect 2590 12316 2596 12328
rect 2648 12316 2654 12368
rect 4706 12356 4712 12368
rect 4619 12328 4712 12356
rect 4706 12316 4712 12328
rect 4764 12356 4770 12368
rect 4764 12328 5672 12356
rect 4764 12316 4770 12328
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 3142 12288 3148 12300
rect 1995 12260 3148 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 4614 12288 4620 12300
rect 3344 12260 4620 12288
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12220 2283 12223
rect 3344 12220 3372 12260
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 5534 12288 5540 12300
rect 5495 12260 5540 12288
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 5644 12288 5672 12328
rect 5718 12316 5724 12368
rect 5776 12365 5782 12368
rect 5776 12359 5840 12365
rect 5776 12325 5794 12359
rect 5828 12325 5840 12359
rect 5776 12319 5840 12325
rect 5776 12316 5782 12319
rect 6546 12316 6552 12368
rect 6604 12356 6610 12368
rect 7024 12356 7052 12396
rect 6604 12328 7052 12356
rect 7644 12359 7702 12365
rect 6604 12316 6610 12328
rect 7644 12325 7656 12359
rect 7690 12356 7702 12359
rect 7742 12356 7748 12368
rect 7690 12328 7748 12356
rect 7690 12325 7702 12328
rect 7644 12319 7702 12325
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 7944 12356 7972 12396
rect 9217 12393 9229 12427
rect 9263 12424 9275 12427
rect 9490 12424 9496 12436
rect 9263 12396 9496 12424
rect 9263 12393 9275 12396
rect 9217 12387 9275 12393
rect 9490 12384 9496 12396
rect 9548 12424 9554 12436
rect 11146 12424 11152 12436
rect 9548 12396 11152 12424
rect 9548 12384 9554 12396
rect 11146 12384 11152 12396
rect 11204 12384 11210 12436
rect 11241 12427 11299 12433
rect 11241 12393 11253 12427
rect 11287 12424 11299 12427
rect 11698 12424 11704 12436
rect 11287 12396 11704 12424
rect 11287 12393 11299 12396
rect 11241 12387 11299 12393
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 12526 12424 12532 12436
rect 12487 12396 12532 12424
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 7944 12328 9536 12356
rect 9398 12288 9404 12300
rect 5644 12260 8432 12288
rect 9359 12260 9404 12288
rect 2271 12192 3372 12220
rect 3421 12223 3479 12229
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 3421 12189 3433 12223
rect 3467 12220 3479 12223
rect 4062 12220 4068 12232
rect 3467 12192 4068 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 3050 12112 3056 12164
rect 3108 12152 3114 12164
rect 3510 12152 3516 12164
rect 3108 12124 3516 12152
rect 3108 12112 3114 12124
rect 3510 12112 3516 12124
rect 3568 12112 3574 12164
rect 4816 12152 4844 12183
rect 4890 12180 4896 12232
rect 4948 12220 4954 12232
rect 7374 12220 7380 12232
rect 4948 12192 4993 12220
rect 7335 12192 7380 12220
rect 4948 12180 4954 12192
rect 7374 12180 7380 12192
rect 7432 12180 7438 12232
rect 8404 12220 8432 12260
rect 9398 12248 9404 12260
rect 9456 12248 9462 12300
rect 9508 12288 9536 12328
rect 9582 12316 9588 12368
rect 9640 12356 9646 12368
rect 10045 12359 10103 12365
rect 10045 12356 10057 12359
rect 9640 12328 10057 12356
rect 9640 12316 9646 12328
rect 10045 12325 10057 12328
rect 10091 12325 10103 12359
rect 10045 12319 10103 12325
rect 10226 12316 10232 12368
rect 10284 12356 10290 12368
rect 10870 12356 10876 12368
rect 10284 12328 10876 12356
rect 10284 12316 10290 12328
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 10962 12316 10968 12368
rect 11020 12356 11026 12368
rect 11330 12356 11336 12368
rect 11020 12328 11192 12356
rect 11243 12328 11336 12356
rect 11020 12316 11026 12328
rect 11054 12288 11060 12300
rect 9508 12260 11060 12288
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 11164 12288 11192 12328
rect 11330 12316 11336 12328
rect 11388 12356 11394 12368
rect 12250 12356 12256 12368
rect 11388 12328 12256 12356
rect 11388 12316 11394 12328
rect 12250 12316 12256 12328
rect 12308 12316 12314 12368
rect 12342 12316 12348 12368
rect 12400 12356 12406 12368
rect 12437 12359 12495 12365
rect 12437 12356 12449 12359
rect 12400 12328 12449 12356
rect 12400 12316 12406 12328
rect 12437 12325 12449 12328
rect 12483 12325 12495 12359
rect 12437 12319 12495 12325
rect 11164 12260 11560 12288
rect 9858 12220 9864 12232
rect 8404 12192 9864 12220
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 10134 12220 10140 12232
rect 10095 12192 10140 12220
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 10284 12192 10333 12220
rect 10284 12180 10290 12192
rect 10321 12189 10333 12192
rect 10367 12220 10379 12223
rect 11425 12223 11483 12229
rect 11425 12220 11437 12223
rect 10367 12192 11437 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 11425 12189 11437 12192
rect 11471 12189 11483 12223
rect 11532 12220 11560 12260
rect 11974 12248 11980 12300
rect 12032 12288 12038 12300
rect 12360 12288 12388 12316
rect 13446 12288 13452 12300
rect 12032 12260 12388 12288
rect 13407 12260 13452 12288
rect 12032 12248 12038 12260
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 13541 12291 13599 12297
rect 13541 12257 13553 12291
rect 13587 12288 13599 12291
rect 14461 12291 14519 12297
rect 14461 12288 14473 12291
rect 13587 12260 14473 12288
rect 13587 12257 13599 12260
rect 13541 12251 13599 12257
rect 14461 12257 14473 12260
rect 14507 12257 14519 12291
rect 14461 12251 14519 12257
rect 12621 12223 12679 12229
rect 12621 12220 12633 12223
rect 11532 12192 12633 12220
rect 11425 12183 11483 12189
rect 12621 12189 12633 12192
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 13170 12180 13176 12232
rect 13228 12220 13234 12232
rect 13556 12220 13584 12251
rect 14550 12248 14556 12300
rect 14608 12288 14614 12300
rect 14826 12288 14832 12300
rect 14608 12260 14832 12288
rect 14608 12248 14614 12260
rect 14826 12248 14832 12260
rect 14884 12248 14890 12300
rect 13228 12192 13584 12220
rect 13817 12223 13875 12229
rect 13228 12180 13234 12192
rect 13817 12189 13829 12223
rect 13863 12220 13875 12223
rect 15378 12220 15384 12232
rect 13863 12192 15384 12220
rect 13863 12189 13875 12192
rect 13817 12183 13875 12189
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 5534 12152 5540 12164
rect 4816 12124 5540 12152
rect 5534 12112 5540 12124
rect 5592 12112 5598 12164
rect 8386 12112 8392 12164
rect 8444 12152 8450 12164
rect 13265 12155 13323 12161
rect 13265 12152 13277 12155
rect 8444 12124 13277 12152
rect 8444 12112 8450 12124
rect 13265 12121 13277 12124
rect 13311 12121 13323 12155
rect 13265 12115 13323 12121
rect 14550 12112 14556 12164
rect 14608 12152 14614 12164
rect 14734 12152 14740 12164
rect 14608 12124 14740 12152
rect 14608 12112 14614 12124
rect 14734 12112 14740 12124
rect 14792 12112 14798 12164
rect 1581 12087 1639 12093
rect 1581 12053 1593 12087
rect 1627 12084 1639 12087
rect 2866 12084 2872 12096
rect 1627 12056 2872 12084
rect 1627 12053 1639 12056
rect 1581 12047 1639 12053
rect 2866 12044 2872 12056
rect 2924 12044 2930 12096
rect 4338 12084 4344 12096
rect 4299 12056 4344 12084
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 5442 12044 5448 12096
rect 5500 12084 5506 12096
rect 8757 12087 8815 12093
rect 8757 12084 8769 12087
rect 5500 12056 8769 12084
rect 5500 12044 5506 12056
rect 8757 12053 8769 12056
rect 8803 12053 8815 12087
rect 8757 12047 8815 12053
rect 8938 12044 8944 12096
rect 8996 12084 9002 12096
rect 9490 12084 9496 12096
rect 8996 12056 9496 12084
rect 8996 12044 9002 12056
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 9674 12084 9680 12096
rect 9635 12056 9680 12084
rect 9674 12044 9680 12056
rect 9732 12044 9738 12096
rect 9858 12044 9864 12096
rect 9916 12084 9922 12096
rect 10042 12084 10048 12096
rect 9916 12056 10048 12084
rect 9916 12044 9922 12056
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 10134 12044 10140 12096
rect 10192 12084 10198 12096
rect 10873 12087 10931 12093
rect 10873 12084 10885 12087
rect 10192 12056 10885 12084
rect 10192 12044 10198 12056
rect 10873 12053 10885 12056
rect 10919 12053 10931 12087
rect 10873 12047 10931 12053
rect 11698 12044 11704 12096
rect 11756 12084 11762 12096
rect 12069 12087 12127 12093
rect 12069 12084 12081 12087
rect 11756 12056 12081 12084
rect 11756 12044 11762 12056
rect 12069 12053 12081 12056
rect 12115 12053 12127 12087
rect 12069 12047 12127 12053
rect 12250 12044 12256 12096
rect 12308 12084 12314 12096
rect 12802 12084 12808 12096
rect 12308 12056 12808 12084
rect 12308 12044 12314 12056
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 14090 12044 14096 12096
rect 14148 12084 14154 12096
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 14148 12056 14657 12084
rect 14148 12044 14154 12056
rect 14645 12053 14657 12056
rect 14691 12053 14703 12087
rect 14645 12047 14703 12053
rect 1104 11994 15824 12016
rect 1104 11942 3447 11994
rect 3499 11942 3511 11994
rect 3563 11942 3575 11994
rect 3627 11942 3639 11994
rect 3691 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 13308 11994
rect 13360 11942 13372 11994
rect 13424 11942 13436 11994
rect 13488 11942 13500 11994
rect 13552 11942 15824 11994
rect 1104 11920 15824 11942
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 2501 11883 2559 11889
rect 2501 11880 2513 11883
rect 1820 11852 2513 11880
rect 1820 11840 1826 11852
rect 2501 11849 2513 11852
rect 2547 11849 2559 11883
rect 2501 11843 2559 11849
rect 3326 11840 3332 11892
rect 3384 11880 3390 11892
rect 3697 11883 3755 11889
rect 3697 11880 3709 11883
rect 3384 11852 3709 11880
rect 3384 11840 3390 11852
rect 3697 11849 3709 11852
rect 3743 11849 3755 11883
rect 3697 11843 3755 11849
rect 4080 11852 8340 11880
rect 1302 11772 1308 11824
rect 1360 11812 1366 11824
rect 3970 11812 3976 11824
rect 1360 11784 3976 11812
rect 1360 11772 1366 11784
rect 3970 11772 3976 11784
rect 4028 11772 4034 11824
rect 3050 11704 3056 11756
rect 3108 11744 3114 11756
rect 3145 11747 3203 11753
rect 3145 11744 3157 11747
rect 3108 11716 3157 11744
rect 3108 11704 3114 11716
rect 3145 11713 3157 11716
rect 3191 11744 3203 11747
rect 3326 11744 3332 11756
rect 3191 11716 3332 11744
rect 3191 11713 3203 11716
rect 3145 11707 3203 11713
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11676 1639 11679
rect 1762 11676 1768 11688
rect 1627 11648 1768 11676
rect 1627 11645 1639 11648
rect 1581 11639 1639 11645
rect 1762 11636 1768 11648
rect 1820 11636 1826 11688
rect 2866 11676 2872 11688
rect 2827 11648 2872 11676
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 4080 11685 4108 11852
rect 8312 11812 8340 11852
rect 8662 11840 8668 11892
rect 8720 11880 8726 11892
rect 10413 11883 10471 11889
rect 10413 11880 10425 11883
rect 8720 11852 10425 11880
rect 8720 11840 8726 11852
rect 10413 11849 10425 11852
rect 10459 11849 10471 11883
rect 10413 11843 10471 11849
rect 11054 11840 11060 11892
rect 11112 11880 11118 11892
rect 13170 11880 13176 11892
rect 11112 11852 13176 11880
rect 11112 11840 11118 11852
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 8938 11812 8944 11824
rect 8312 11784 8944 11812
rect 8938 11772 8944 11784
rect 8996 11772 9002 11824
rect 11422 11812 11428 11824
rect 9048 11784 11428 11812
rect 4246 11744 4252 11756
rect 4207 11716 4252 11744
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 7374 11744 7380 11756
rect 7335 11716 7380 11744
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 8662 11704 8668 11756
rect 8720 11744 8726 11756
rect 9048 11744 9076 11784
rect 11422 11772 11428 11784
rect 11480 11772 11486 11824
rect 12437 11815 12495 11821
rect 12437 11781 12449 11815
rect 12483 11812 12495 11815
rect 12710 11812 12716 11824
rect 12483 11784 12716 11812
rect 12483 11781 12495 11784
rect 12437 11775 12495 11781
rect 12710 11772 12716 11784
rect 12768 11772 12774 11824
rect 8720 11716 9076 11744
rect 9769 11747 9827 11753
rect 8720 11704 8726 11716
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 10870 11744 10876 11756
rect 10831 11716 10876 11744
rect 9769 11707 9827 11713
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11645 4123 11679
rect 4890 11676 4896 11688
rect 4803 11648 4896 11676
rect 4065 11639 4123 11645
rect 4890 11636 4896 11648
rect 4948 11676 4954 11688
rect 5718 11676 5724 11688
rect 4948 11648 5724 11676
rect 4948 11636 4954 11648
rect 5718 11636 5724 11648
rect 5776 11636 5782 11688
rect 7650 11685 7656 11688
rect 7644 11676 7656 11685
rect 7611 11648 7656 11676
rect 7644 11639 7656 11648
rect 7708 11676 7714 11688
rect 9784 11676 9812 11707
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 11057 11747 11115 11753
rect 11057 11713 11069 11747
rect 11103 11744 11115 11747
rect 11238 11744 11244 11756
rect 11103 11716 11244 11744
rect 11103 11713 11115 11716
rect 11057 11707 11115 11713
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 11348 11716 13001 11744
rect 10226 11676 10232 11688
rect 7708 11648 10232 11676
rect 7650 11636 7656 11639
rect 7708 11636 7714 11648
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 10502 11636 10508 11688
rect 10560 11676 10566 11688
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 10560 11648 10793 11676
rect 10560 11636 10566 11648
rect 10781 11645 10793 11648
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 1857 11611 1915 11617
rect 1857 11577 1869 11611
rect 1903 11608 1915 11611
rect 2961 11611 3019 11617
rect 1903 11580 2912 11608
rect 1903 11577 1915 11580
rect 1857 11571 1915 11577
rect 2884 11540 2912 11580
rect 2961 11577 2973 11611
rect 3007 11608 3019 11611
rect 4246 11608 4252 11620
rect 3007 11580 4252 11608
rect 3007 11577 3019 11580
rect 2961 11571 3019 11577
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 5166 11617 5172 11620
rect 5160 11608 5172 11617
rect 5127 11580 5172 11608
rect 5160 11571 5172 11580
rect 5166 11568 5172 11571
rect 5224 11568 5230 11620
rect 8662 11608 8668 11620
rect 6196 11580 8668 11608
rect 3050 11540 3056 11552
rect 2884 11512 3056 11540
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 4157 11543 4215 11549
rect 4157 11509 4169 11543
rect 4203 11540 4215 11543
rect 6196 11540 6224 11580
rect 8662 11568 8668 11580
rect 8720 11568 8726 11620
rect 9582 11608 9588 11620
rect 9543 11580 9588 11608
rect 9582 11568 9588 11580
rect 9640 11568 9646 11620
rect 4203 11512 6224 11540
rect 6273 11543 6331 11549
rect 4203 11509 4215 11512
rect 4157 11503 4215 11509
rect 6273 11509 6285 11543
rect 6319 11540 6331 11543
rect 6914 11540 6920 11552
rect 6319 11512 6920 11540
rect 6319 11509 6331 11512
rect 6273 11503 6331 11509
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 8757 11543 8815 11549
rect 8757 11509 8769 11543
rect 8803 11540 8815 11543
rect 8938 11540 8944 11552
rect 8803 11512 8944 11540
rect 8803 11509 8815 11512
rect 8757 11503 8815 11509
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9214 11540 9220 11552
rect 9175 11512 9220 11540
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 9677 11543 9735 11549
rect 9677 11509 9689 11543
rect 9723 11540 9735 11543
rect 9858 11540 9864 11552
rect 9723 11512 9864 11540
rect 9723 11509 9735 11512
rect 9677 11503 9735 11509
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 10226 11500 10232 11552
rect 10284 11540 10290 11552
rect 11348 11540 11376 11716
rect 12989 11713 13001 11716
rect 13035 11744 13047 11747
rect 13538 11744 13544 11756
rect 13035 11716 13544 11744
rect 13035 11713 13047 11716
rect 12989 11707 13047 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 13909 11747 13967 11753
rect 13909 11713 13921 11747
rect 13955 11744 13967 11747
rect 14918 11744 14924 11756
rect 13955 11716 14924 11744
rect 13955 11713 13967 11716
rect 13909 11707 13967 11713
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11676 11667 11679
rect 13633 11679 13691 11685
rect 11655 11648 13584 11676
rect 11655 11645 11667 11648
rect 11609 11639 11667 11645
rect 12805 11611 12863 11617
rect 12805 11577 12817 11611
rect 12851 11608 12863 11611
rect 13170 11608 13176 11620
rect 12851 11580 13176 11608
rect 12851 11577 12863 11580
rect 12805 11571 12863 11577
rect 13170 11568 13176 11580
rect 13228 11568 13234 11620
rect 13556 11608 13584 11648
rect 13633 11645 13645 11679
rect 13679 11676 13691 11679
rect 13722 11676 13728 11688
rect 13679 11648 13728 11676
rect 13679 11645 13691 11648
rect 13633 11639 13691 11645
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 13814 11636 13820 11688
rect 13872 11676 13878 11688
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 13872 11648 14565 11676
rect 13872 11636 13878 11648
rect 14553 11645 14565 11648
rect 14599 11645 14611 11679
rect 14553 11639 14611 11645
rect 13998 11608 14004 11620
rect 13556 11580 14004 11608
rect 13998 11568 14004 11580
rect 14056 11568 14062 11620
rect 14829 11611 14887 11617
rect 14829 11577 14841 11611
rect 14875 11608 14887 11611
rect 16390 11608 16396 11620
rect 14875 11580 16396 11608
rect 14875 11577 14887 11580
rect 14829 11571 14887 11577
rect 16390 11568 16396 11580
rect 16448 11568 16454 11620
rect 10284 11512 11376 11540
rect 11793 11543 11851 11549
rect 10284 11500 10290 11512
rect 11793 11509 11805 11543
rect 11839 11540 11851 11543
rect 12342 11540 12348 11552
rect 11839 11512 12348 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 12894 11540 12900 11552
rect 12855 11512 12900 11540
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 1104 11450 15824 11472
rect 1104 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 6104 11450
rect 6156 11398 10843 11450
rect 10895 11398 10907 11450
rect 10959 11398 10971 11450
rect 11023 11398 11035 11450
rect 11087 11398 15824 11450
rect 1104 11376 15824 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 4522 11336 4528 11348
rect 3191 11308 4528 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 4617 11339 4675 11345
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 8754 11336 8760 11348
rect 4663 11308 8760 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 8754 11296 8760 11308
rect 8812 11296 8818 11348
rect 9214 11296 9220 11348
rect 9272 11336 9278 11348
rect 10134 11336 10140 11348
rect 9272 11308 9720 11336
rect 10095 11308 10140 11336
rect 9272 11296 9278 11308
rect 4985 11271 5043 11277
rect 4985 11237 4997 11271
rect 5031 11268 5043 11271
rect 9582 11268 9588 11280
rect 5031 11240 9588 11268
rect 5031 11237 5043 11240
rect 4985 11231 5043 11237
rect 9582 11228 9588 11240
rect 9640 11228 9646 11280
rect 9692 11268 9720 11308
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 11333 11339 11391 11345
rect 11333 11305 11345 11339
rect 11379 11336 11391 11339
rect 11698 11336 11704 11348
rect 11379 11308 11704 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 13078 11296 13084 11348
rect 13136 11336 13142 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 13136 11308 13277 11336
rect 13136 11296 13142 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 10045 11271 10103 11277
rect 10045 11268 10057 11271
rect 9692 11240 10057 11268
rect 10045 11237 10057 11240
rect 10091 11237 10103 11271
rect 12529 11271 12587 11277
rect 12529 11268 12541 11271
rect 10045 11231 10103 11237
rect 10796 11240 12541 11268
rect 1946 11200 1952 11212
rect 1907 11172 1952 11200
rect 1946 11160 1952 11172
rect 2004 11160 2010 11212
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11200 2099 11203
rect 2406 11200 2412 11212
rect 2087 11172 2412 11200
rect 2087 11169 2099 11172
rect 2041 11163 2099 11169
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 2498 11160 2504 11212
rect 2556 11200 2562 11212
rect 5077 11203 5135 11209
rect 5077 11200 5089 11203
rect 2556 11172 5089 11200
rect 2556 11160 2562 11172
rect 5077 11169 5089 11172
rect 5123 11200 5135 11203
rect 5626 11200 5632 11212
rect 5123 11172 5632 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 5810 11200 5816 11212
rect 5771 11172 5816 11200
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 6080 11203 6138 11209
rect 6080 11169 6092 11203
rect 6126 11200 6138 11203
rect 6914 11200 6920 11212
rect 6126 11172 6920 11200
rect 6126 11169 6138 11172
rect 6080 11163 6138 11169
rect 6914 11160 6920 11172
rect 6972 11200 6978 11212
rect 7742 11200 7748 11212
rect 6972 11172 7748 11200
rect 6972 11160 6978 11172
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 7920 11203 7978 11209
rect 7920 11169 7932 11203
rect 7966 11200 7978 11203
rect 8938 11200 8944 11212
rect 7966 11172 8944 11200
rect 7966 11169 7978 11172
rect 7920 11163 7978 11169
rect 8938 11160 8944 11172
rect 8996 11200 9002 11212
rect 10686 11200 10692 11212
rect 8996 11172 10692 11200
rect 8996 11160 9002 11172
rect 1670 11092 1676 11144
rect 1728 11132 1734 11144
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 1728 11104 2145 11132
rect 1728 11092 1734 11104
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 3234 11132 3240 11144
rect 3195 11104 3240 11132
rect 2133 11095 2191 11101
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 4430 11132 4436 11144
rect 3467 11104 4436 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 4430 11092 4436 11104
rect 4488 11092 4494 11144
rect 5258 11132 5264 11144
rect 5171 11104 5264 11132
rect 5258 11092 5264 11104
rect 5316 11132 5322 11144
rect 5442 11132 5448 11144
rect 5316 11104 5448 11132
rect 5316 11092 5322 11104
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 7374 11092 7380 11144
rect 7432 11132 7438 11144
rect 7653 11135 7711 11141
rect 7653 11132 7665 11135
rect 7432 11104 7665 11132
rect 7432 11092 7438 11104
rect 7653 11101 7665 11104
rect 7699 11101 7711 11135
rect 7653 11095 7711 11101
rect 9030 11092 9036 11144
rect 9088 11092 9094 11144
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 9306 11132 9312 11144
rect 9180 11104 9312 11132
rect 9180 11092 9186 11104
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 10336 11141 10364 11172
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11101 10379 11135
rect 10796 11132 10824 11240
rect 12529 11237 12541 11240
rect 12575 11237 12587 11271
rect 12529 11231 12587 11237
rect 13722 11228 13728 11280
rect 13780 11268 13786 11280
rect 13780 11240 14504 11268
rect 13780 11228 13786 11240
rect 11054 11160 11060 11212
rect 11112 11200 11118 11212
rect 11241 11203 11299 11209
rect 11241 11200 11253 11203
rect 11112 11172 11253 11200
rect 11112 11160 11118 11172
rect 11241 11169 11253 11172
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 11330 11160 11336 11212
rect 11388 11200 11394 11212
rect 11388 11172 11468 11200
rect 11388 11160 11394 11172
rect 11440 11141 11468 11172
rect 11698 11160 11704 11212
rect 11756 11200 11762 11212
rect 11882 11200 11888 11212
rect 11756 11172 11888 11200
rect 11756 11160 11762 11172
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 12434 11200 12440 11212
rect 12395 11172 12440 11200
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 13630 11200 13636 11212
rect 13591 11172 13636 11200
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 14476 11209 14504 11240
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11169 14519 11203
rect 14461 11163 14519 11169
rect 10321 11095 10379 11101
rect 10416 11104 10824 11132
rect 11425 11135 11483 11141
rect 2777 11067 2835 11073
rect 2777 11033 2789 11067
rect 2823 11064 2835 11067
rect 4522 11064 4528 11076
rect 2823 11036 4528 11064
rect 2823 11033 2835 11036
rect 2777 11027 2835 11033
rect 4522 11024 4528 11036
rect 4580 11024 4586 11076
rect 9048 11064 9076 11092
rect 9582 11064 9588 11076
rect 9048 11036 9588 11064
rect 9582 11024 9588 11036
rect 9640 11024 9646 11076
rect 9677 11067 9735 11073
rect 9677 11033 9689 11067
rect 9723 11064 9735 11067
rect 9766 11064 9772 11076
rect 9723 11036 9772 11064
rect 9723 11033 9735 11036
rect 9677 11027 9735 11033
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 9950 11024 9956 11076
rect 10008 11064 10014 11076
rect 10416 11064 10444 11104
rect 11425 11101 11437 11135
rect 11471 11101 11483 11135
rect 12621 11135 12679 11141
rect 12621 11132 12633 11135
rect 11425 11095 11483 11101
rect 11624 11104 12633 11132
rect 10008 11036 10444 11064
rect 10008 11024 10014 11036
rect 10502 11024 10508 11076
rect 10560 11064 10566 11076
rect 10873 11067 10931 11073
rect 10873 11064 10885 11067
rect 10560 11036 10885 11064
rect 10560 11024 10566 11036
rect 10873 11033 10885 11036
rect 10919 11033 10931 11067
rect 10873 11027 10931 11033
rect 10962 11024 10968 11076
rect 11020 11064 11026 11076
rect 11624 11064 11652 11104
rect 12621 11101 12633 11104
rect 12667 11101 12679 11135
rect 13722 11132 13728 11144
rect 13683 11104 13728 11132
rect 12621 11095 12679 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13817 11135 13875 11141
rect 13817 11101 13829 11135
rect 13863 11101 13875 11135
rect 13817 11095 13875 11101
rect 11020 11036 11652 11064
rect 12069 11067 12127 11073
rect 11020 11024 11026 11036
rect 12069 11033 12081 11067
rect 12115 11064 12127 11067
rect 12710 11064 12716 11076
rect 12115 11036 12716 11064
rect 12115 11033 12127 11036
rect 12069 11027 12127 11033
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 13538 11024 13544 11076
rect 13596 11064 13602 11076
rect 13832 11064 13860 11095
rect 13596 11036 13860 11064
rect 14645 11067 14703 11073
rect 13596 11024 13602 11036
rect 14645 11033 14657 11067
rect 14691 11064 14703 11067
rect 14826 11064 14832 11076
rect 14691 11036 14832 11064
rect 14691 11033 14703 11036
rect 14645 11027 14703 11033
rect 14826 11024 14832 11036
rect 14884 11024 14890 11076
rect 1578 10956 1584 11008
rect 1636 10996 1642 11008
rect 2682 10996 2688 11008
rect 1636 10968 2688 10996
rect 1636 10956 1642 10968
rect 2682 10956 2688 10968
rect 2740 10996 2746 11008
rect 6730 10996 6736 11008
rect 2740 10968 6736 10996
rect 2740 10956 2746 10968
rect 6730 10956 6736 10968
rect 6788 10956 6794 11008
rect 7190 10996 7196 11008
rect 7103 10968 7196 10996
rect 7190 10956 7196 10968
rect 7248 10996 7254 11008
rect 7650 10996 7656 11008
rect 7248 10968 7656 10996
rect 7248 10956 7254 10968
rect 7650 10956 7656 10968
rect 7708 10956 7714 11008
rect 9030 10996 9036 11008
rect 8943 10968 9036 10996
rect 9030 10956 9036 10968
rect 9088 10996 9094 11008
rect 10778 10996 10784 11008
rect 9088 10968 10784 10996
rect 9088 10956 9094 10968
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 11882 10956 11888 11008
rect 11940 10996 11946 11008
rect 15286 10996 15292 11008
rect 11940 10968 15292 10996
rect 11940 10956 11946 10968
rect 15286 10956 15292 10968
rect 15344 10956 15350 11008
rect 1104 10906 15824 10928
rect 1104 10854 3447 10906
rect 3499 10854 3511 10906
rect 3563 10854 3575 10906
rect 3627 10854 3639 10906
rect 3691 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 13308 10906
rect 13360 10854 13372 10906
rect 13424 10854 13436 10906
rect 13488 10854 13500 10906
rect 13552 10854 15824 10906
rect 1104 10832 15824 10854
rect 3142 10752 3148 10804
rect 3200 10792 3206 10804
rect 3697 10795 3755 10801
rect 3697 10792 3709 10795
rect 3200 10764 3709 10792
rect 3200 10752 3206 10764
rect 3697 10761 3709 10764
rect 3743 10761 3755 10795
rect 5166 10792 5172 10804
rect 3697 10755 3755 10761
rect 4172 10764 5172 10792
rect 2501 10727 2559 10733
rect 2501 10693 2513 10727
rect 2547 10693 2559 10727
rect 2501 10687 2559 10693
rect 1581 10591 1639 10597
rect 1581 10557 1593 10591
rect 1627 10588 1639 10591
rect 2516 10588 2544 10687
rect 2682 10616 2688 10668
rect 2740 10656 2746 10668
rect 2961 10659 3019 10665
rect 2961 10656 2973 10659
rect 2740 10628 2973 10656
rect 2740 10616 2746 10628
rect 2961 10625 2973 10628
rect 3007 10625 3019 10659
rect 2961 10619 3019 10625
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10656 3203 10659
rect 4172 10656 4200 10764
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 5592 10764 6837 10792
rect 5592 10752 5598 10764
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 6825 10755 6883 10761
rect 8021 10795 8079 10801
rect 8021 10761 8033 10795
rect 8067 10792 8079 10795
rect 9398 10792 9404 10804
rect 8067 10764 9404 10792
rect 8067 10761 8079 10764
rect 8021 10755 8079 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 10321 10795 10379 10801
rect 10321 10761 10333 10795
rect 10367 10792 10379 10795
rect 11054 10792 11060 10804
rect 10367 10764 11060 10792
rect 10367 10761 10379 10764
rect 10321 10755 10379 10761
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11388 10764 11713 10792
rect 11388 10752 11394 10764
rect 11701 10761 11713 10764
rect 11747 10761 11759 10795
rect 13630 10792 13636 10804
rect 13591 10764 13636 10792
rect 11701 10755 11759 10761
rect 13630 10752 13636 10764
rect 13688 10752 13694 10804
rect 10686 10684 10692 10736
rect 10744 10724 10750 10736
rect 10744 10696 10916 10724
rect 10744 10684 10750 10696
rect 3191 10628 4200 10656
rect 4341 10659 4399 10665
rect 3191 10625 3203 10628
rect 3145 10619 3203 10625
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4430 10656 4436 10668
rect 4387 10628 4436 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4430 10616 4436 10628
rect 4488 10616 4494 10668
rect 4890 10656 4896 10668
rect 4851 10628 4896 10656
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 7282 10656 7288 10668
rect 7243 10628 7288 10656
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 7926 10656 7932 10668
rect 7515 10628 7932 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 8128 10628 8616 10656
rect 4062 10588 4068 10600
rect 1627 10560 2544 10588
rect 4023 10560 4068 10588
rect 1627 10557 1639 10560
rect 1581 10551 1639 10557
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4157 10591 4215 10597
rect 4157 10557 4169 10591
rect 4203 10588 4215 10591
rect 8128 10588 8156 10628
rect 4203 10560 8156 10588
rect 4203 10557 4215 10560
rect 4157 10551 4215 10557
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 8481 10591 8539 10597
rect 8260 10560 8305 10588
rect 8260 10548 8266 10560
rect 8481 10557 8493 10591
rect 8527 10557 8539 10591
rect 8588 10588 8616 10628
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10502 10656 10508 10668
rect 10192 10628 10508 10656
rect 10192 10616 10198 10628
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 10594 10616 10600 10668
rect 10652 10656 10658 10668
rect 10888 10665 10916 10696
rect 10962 10684 10968 10736
rect 11020 10724 11026 10736
rect 11514 10724 11520 10736
rect 11020 10696 11520 10724
rect 11020 10684 11026 10696
rect 11514 10684 11520 10696
rect 11572 10684 11578 10736
rect 11882 10724 11888 10736
rect 11624 10696 11888 10724
rect 10873 10659 10931 10665
rect 10652 10628 10732 10656
rect 10652 10616 10658 10628
rect 10704 10597 10732 10628
rect 10873 10625 10885 10659
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11330 10656 11336 10668
rect 11112 10628 11336 10656
rect 11112 10616 11118 10628
rect 11330 10616 11336 10628
rect 11388 10616 11394 10668
rect 11624 10656 11652 10696
rect 11882 10684 11888 10696
rect 11940 10684 11946 10736
rect 12253 10727 12311 10733
rect 12253 10693 12265 10727
rect 12299 10724 12311 10727
rect 12299 10696 14872 10724
rect 12299 10693 12311 10696
rect 12253 10687 12311 10693
rect 11532 10628 11652 10656
rect 11532 10597 11560 10628
rect 12526 10616 12532 10668
rect 12584 10656 12590 10668
rect 12897 10659 12955 10665
rect 12897 10656 12909 10659
rect 12584 10628 12909 10656
rect 12584 10616 12590 10628
rect 12897 10625 12909 10628
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 10689 10591 10747 10597
rect 8588 10560 10548 10588
rect 8481 10551 8539 10557
rect 1854 10520 1860 10532
rect 1815 10492 1860 10520
rect 1854 10480 1860 10492
rect 1912 10480 1918 10532
rect 3326 10480 3332 10532
rect 3384 10520 3390 10532
rect 3384 10492 4108 10520
rect 3384 10480 3390 10492
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 2869 10455 2927 10461
rect 2869 10452 2881 10455
rect 2832 10424 2881 10452
rect 2832 10412 2838 10424
rect 2869 10421 2881 10424
rect 2915 10421 2927 10455
rect 2869 10415 2927 10421
rect 3142 10412 3148 10464
rect 3200 10452 3206 10464
rect 3878 10452 3884 10464
rect 3200 10424 3884 10452
rect 3200 10412 3206 10424
rect 3878 10412 3884 10424
rect 3936 10412 3942 10464
rect 4080 10452 4108 10492
rect 4614 10480 4620 10532
rect 4672 10520 4678 10532
rect 5138 10523 5196 10529
rect 5138 10520 5150 10523
rect 4672 10492 5150 10520
rect 4672 10480 4678 10492
rect 5138 10489 5150 10492
rect 5184 10489 5196 10523
rect 5138 10483 5196 10489
rect 7006 10480 7012 10532
rect 7064 10520 7070 10532
rect 7193 10523 7251 10529
rect 7193 10520 7205 10523
rect 7064 10492 7205 10520
rect 7064 10480 7070 10492
rect 7193 10489 7205 10492
rect 7239 10489 7251 10523
rect 7193 10483 7251 10489
rect 7374 10480 7380 10532
rect 7432 10520 7438 10532
rect 8496 10520 8524 10551
rect 7432 10492 8524 10520
rect 8748 10523 8806 10529
rect 7432 10480 7438 10492
rect 8748 10489 8760 10523
rect 8794 10520 8806 10523
rect 9030 10520 9036 10532
rect 8794 10492 9036 10520
rect 8794 10489 8806 10492
rect 8748 10483 8806 10489
rect 9030 10480 9036 10492
rect 9088 10480 9094 10532
rect 10410 10520 10416 10532
rect 9876 10492 10416 10520
rect 6273 10455 6331 10461
rect 6273 10452 6285 10455
rect 4080 10424 6285 10452
rect 6273 10421 6285 10424
rect 6319 10421 6331 10455
rect 6273 10415 6331 10421
rect 6362 10412 6368 10464
rect 6420 10452 6426 10464
rect 9766 10452 9772 10464
rect 6420 10424 9772 10452
rect 6420 10412 6426 10424
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 9876 10461 9904 10492
rect 10410 10480 10416 10492
rect 10468 10480 10474 10532
rect 10520 10520 10548 10560
rect 10689 10557 10701 10591
rect 10735 10557 10747 10591
rect 10689 10551 10747 10557
rect 11517 10591 11575 10597
rect 11517 10557 11529 10591
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 11532 10520 11560 10551
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12492 10560 12817 10588
rect 12492 10548 12498 10560
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 10520 10492 11560 10520
rect 11882 10480 11888 10532
rect 11940 10520 11946 10532
rect 13004 10520 13032 10619
rect 13630 10616 13636 10668
rect 13688 10656 13694 10668
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 13688 10628 14197 10656
rect 13688 10616 13694 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 14001 10591 14059 10597
rect 14001 10557 14013 10591
rect 14047 10588 14059 10591
rect 14366 10588 14372 10600
rect 14047 10560 14372 10588
rect 14047 10557 14059 10560
rect 14001 10551 14059 10557
rect 14366 10548 14372 10560
rect 14424 10548 14430 10600
rect 14844 10597 14872 10696
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 16758 10588 16764 10600
rect 14875 10560 16764 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 16758 10548 16764 10560
rect 16816 10548 16822 10600
rect 11940 10492 13032 10520
rect 14093 10523 14151 10529
rect 11940 10480 11946 10492
rect 14093 10489 14105 10523
rect 14139 10520 14151 10523
rect 14642 10520 14648 10532
rect 14139 10492 14648 10520
rect 14139 10489 14151 10492
rect 14093 10483 14151 10489
rect 14384 10464 14412 10492
rect 14642 10480 14648 10492
rect 14700 10480 14706 10532
rect 9861 10455 9919 10461
rect 9861 10421 9873 10455
rect 9907 10421 9919 10455
rect 9861 10415 9919 10421
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10008 10424 10793 10452
rect 10008 10412 10014 10424
rect 10781 10421 10793 10424
rect 10827 10452 10839 10455
rect 12253 10455 12311 10461
rect 12253 10452 12265 10455
rect 10827 10424 12265 10452
rect 10827 10421 10839 10424
rect 10781 10415 10839 10421
rect 12253 10421 12265 10424
rect 12299 10421 12311 10455
rect 12253 10415 12311 10421
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12492 10424 12537 10452
rect 12492 10412 12498 10424
rect 14366 10412 14372 10464
rect 14424 10412 14430 10464
rect 15010 10452 15016 10464
rect 14971 10424 15016 10452
rect 15010 10412 15016 10424
rect 15068 10412 15074 10464
rect 1104 10362 15824 10384
rect 1104 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 6104 10362
rect 6156 10310 10843 10362
rect 10895 10310 10907 10362
rect 10959 10310 10971 10362
rect 11023 10310 11035 10362
rect 11087 10310 15824 10362
rect 1104 10288 15824 10310
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 2498 10248 2504 10260
rect 1995 10220 2504 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 2832 10220 2877 10248
rect 2832 10208 2838 10220
rect 3786 10208 3792 10260
rect 3844 10248 3850 10260
rect 4062 10248 4068 10260
rect 3844 10220 4068 10248
rect 3844 10208 3850 10220
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4246 10248 4252 10260
rect 4207 10220 4252 10248
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 4338 10208 4344 10260
rect 4396 10248 4402 10260
rect 4709 10251 4767 10257
rect 4709 10248 4721 10251
rect 4396 10220 4721 10248
rect 4396 10208 4402 10220
rect 4709 10217 4721 10220
rect 4755 10217 4767 10251
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 4709 10211 4767 10217
rect 6441 10220 10885 10248
rect 4522 10140 4528 10192
rect 4580 10180 4586 10192
rect 4617 10183 4675 10189
rect 4617 10180 4629 10183
rect 4580 10152 4629 10180
rect 4580 10140 4586 10152
rect 4617 10149 4629 10152
rect 4663 10149 4675 10183
rect 6441 10180 6469 10220
rect 10873 10217 10885 10220
rect 10919 10217 10931 10251
rect 11330 10248 11336 10260
rect 11243 10220 11336 10248
rect 10873 10211 10931 10217
rect 11330 10208 11336 10220
rect 11388 10248 11394 10260
rect 11606 10248 11612 10260
rect 11388 10220 11612 10248
rect 11388 10208 11394 10220
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 11790 10208 11796 10260
rect 11848 10248 11854 10260
rect 12529 10251 12587 10257
rect 12529 10248 12541 10251
rect 11848 10220 12541 10248
rect 11848 10208 11854 10220
rect 12529 10217 12541 10220
rect 12575 10217 12587 10251
rect 12529 10211 12587 10217
rect 13265 10251 13323 10257
rect 13265 10217 13277 10251
rect 13311 10248 13323 10251
rect 13722 10248 13728 10260
rect 13311 10220 13728 10248
rect 13311 10217 13323 10220
rect 13265 10211 13323 10217
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 4617 10143 4675 10149
rect 5552 10152 6469 10180
rect 2041 10115 2099 10121
rect 2041 10081 2053 10115
rect 2087 10112 2099 10115
rect 2774 10112 2780 10124
rect 2087 10084 2780 10112
rect 2087 10081 2099 10084
rect 2041 10075 2099 10081
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 3145 10115 3203 10121
rect 3145 10081 3157 10115
rect 3191 10081 3203 10115
rect 3145 10075 3203 10081
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 5552 10112 5580 10152
rect 7466 10140 7472 10192
rect 7524 10189 7530 10192
rect 7524 10183 7588 10189
rect 7524 10149 7542 10183
rect 7576 10149 7588 10183
rect 7524 10143 7588 10149
rect 7524 10140 7530 10143
rect 7650 10140 7656 10192
rect 7708 10180 7714 10192
rect 9858 10180 9864 10192
rect 7708 10152 9864 10180
rect 7708 10140 7714 10152
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 10045 10183 10103 10189
rect 10045 10149 10057 10183
rect 10091 10180 10103 10183
rect 10686 10180 10692 10192
rect 10091 10152 10692 10180
rect 10091 10149 10103 10152
rect 10045 10143 10103 10149
rect 10686 10140 10692 10152
rect 10744 10180 10750 10192
rect 11054 10180 11060 10192
rect 10744 10152 11060 10180
rect 10744 10140 10750 10152
rect 11054 10140 11060 10152
rect 11112 10140 11118 10192
rect 11241 10183 11299 10189
rect 11241 10149 11253 10183
rect 11287 10180 11299 10183
rect 11514 10180 11520 10192
rect 11287 10152 11520 10180
rect 11287 10149 11299 10152
rect 11241 10143 11299 10149
rect 11514 10140 11520 10152
rect 11572 10180 11578 10192
rect 12066 10180 12072 10192
rect 11572 10152 12072 10180
rect 11572 10140 11578 10152
rect 12066 10140 12072 10152
rect 12124 10140 12130 10192
rect 12437 10183 12495 10189
rect 12437 10149 12449 10183
rect 12483 10180 12495 10183
rect 13446 10180 13452 10192
rect 12483 10152 13452 10180
rect 12483 10149 12495 10152
rect 12437 10143 12495 10149
rect 13446 10140 13452 10152
rect 13504 10180 13510 10192
rect 13814 10180 13820 10192
rect 13504 10152 13820 10180
rect 13504 10140 13510 10152
rect 13814 10140 13820 10152
rect 13872 10140 13878 10192
rect 15654 10180 15660 10192
rect 13924 10152 15660 10180
rect 5718 10121 5724 10124
rect 5712 10112 5724 10121
rect 3283 10084 5580 10112
rect 5631 10084 5724 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 5712 10075 5724 10084
rect 5776 10112 5782 10124
rect 7190 10112 7196 10124
rect 5776 10084 7196 10112
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 2866 10044 2872 10056
rect 2271 10016 2872 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3160 9976 3188 10075
rect 5718 10072 5724 10075
rect 5776 10072 5782 10084
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 9306 10112 9312 10124
rect 7340 10084 7385 10112
rect 9267 10084 9312 10112
rect 7340 10072 7346 10084
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 10134 10112 10140 10124
rect 9876 10084 10140 10112
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10044 3479 10047
rect 3878 10044 3884 10056
rect 3467 10016 3884 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 4801 10047 4859 10053
rect 4801 10044 4813 10047
rect 4672 10016 4813 10044
rect 4672 10004 4678 10016
rect 4801 10013 4813 10016
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 4522 9976 4528 9988
rect 3160 9948 4528 9976
rect 4522 9936 4528 9948
rect 4580 9936 4586 9988
rect 4816 9976 4844 10007
rect 4890 10004 4896 10056
rect 4948 10044 4954 10056
rect 5445 10047 5503 10053
rect 5445 10044 5457 10047
rect 4948 10016 5457 10044
rect 4948 10004 4954 10016
rect 5445 10013 5457 10016
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 6822 10004 6828 10056
rect 6880 10044 6886 10056
rect 7300 10044 7328 10072
rect 9876 10056 9904 10084
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 10410 10112 10416 10124
rect 10336 10084 10416 10112
rect 6880 10016 7328 10044
rect 6880 10004 6886 10016
rect 9858 10004 9864 10056
rect 9916 10004 9922 10056
rect 10336 10053 10364 10084
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 12342 10112 12348 10124
rect 10560 10084 12348 10112
rect 10560 10072 10566 10084
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 13354 10072 13360 10124
rect 13412 10112 13418 10124
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 13412 10084 13645 10112
rect 13412 10072 13418 10084
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 13722 10072 13728 10124
rect 13780 10112 13786 10124
rect 13924 10112 13952 10152
rect 15654 10140 15660 10152
rect 15712 10140 15718 10192
rect 13780 10084 13952 10112
rect 13780 10072 13786 10084
rect 14182 10072 14188 10124
rect 14240 10112 14246 10124
rect 14461 10115 14519 10121
rect 14461 10112 14473 10115
rect 14240 10084 14473 10112
rect 14240 10072 14246 10084
rect 14461 10081 14473 10084
rect 14507 10081 14519 10115
rect 14461 10075 14519 10081
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10013 10379 10047
rect 10321 10007 10379 10013
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10044 11575 10047
rect 11882 10044 11888 10056
rect 11563 10016 11888 10044
rect 11563 10013 11575 10016
rect 11517 10007 11575 10013
rect 8665 9979 8723 9985
rect 4816 9948 5028 9976
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 2590 9908 2596 9920
rect 1627 9880 2596 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 3786 9868 3792 9920
rect 3844 9908 3850 9920
rect 4890 9908 4896 9920
rect 3844 9880 4896 9908
rect 3844 9868 3850 9880
rect 4890 9868 4896 9880
rect 4948 9868 4954 9920
rect 5000 9908 5028 9948
rect 8665 9945 8677 9979
rect 8711 9976 8723 9979
rect 10410 9976 10416 9988
rect 8711 9948 10416 9976
rect 8711 9945 8723 9948
rect 8665 9939 8723 9945
rect 6825 9911 6883 9917
rect 6825 9908 6837 9911
rect 5000 9880 6837 9908
rect 6825 9877 6837 9880
rect 6871 9877 6883 9911
rect 6825 9871 6883 9877
rect 8018 9868 8024 9920
rect 8076 9908 8082 9920
rect 8680 9908 8708 9939
rect 10410 9936 10416 9948
rect 10468 9976 10474 9988
rect 11532 9976 11560 10007
rect 11882 10004 11888 10016
rect 11940 10004 11946 10056
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10044 12771 10047
rect 13538 10044 13544 10056
rect 12759 10016 13544 10044
rect 12759 10013 12771 10016
rect 12713 10007 12771 10013
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 13817 10047 13875 10053
rect 13817 10013 13829 10047
rect 13863 10013 13875 10047
rect 13817 10007 13875 10013
rect 10468 9948 11560 9976
rect 10468 9936 10474 9948
rect 13722 9936 13728 9988
rect 13780 9976 13786 9988
rect 13832 9976 13860 10007
rect 14642 9976 14648 9988
rect 13780 9948 13860 9976
rect 14603 9948 14648 9976
rect 13780 9936 13786 9948
rect 14642 9936 14648 9948
rect 14700 9936 14706 9988
rect 8076 9880 8708 9908
rect 9125 9911 9183 9917
rect 8076 9868 8082 9880
rect 9125 9877 9137 9911
rect 9171 9908 9183 9911
rect 9398 9908 9404 9920
rect 9171 9880 9404 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 9677 9911 9735 9917
rect 9677 9908 9689 9911
rect 9548 9880 9689 9908
rect 9548 9868 9554 9880
rect 9677 9877 9689 9880
rect 9723 9877 9735 9911
rect 9677 9871 9735 9877
rect 9766 9868 9772 9920
rect 9824 9908 9830 9920
rect 12069 9911 12127 9917
rect 12069 9908 12081 9911
rect 9824 9880 12081 9908
rect 9824 9868 9830 9880
rect 12069 9877 12081 9880
rect 12115 9877 12127 9911
rect 12069 9871 12127 9877
rect 13998 9868 14004 9920
rect 14056 9908 14062 9920
rect 14918 9908 14924 9920
rect 14056 9880 14924 9908
rect 14056 9868 14062 9880
rect 14918 9868 14924 9880
rect 14976 9868 14982 9920
rect 1104 9818 15824 9840
rect 1104 9766 3447 9818
rect 3499 9766 3511 9818
rect 3563 9766 3575 9818
rect 3627 9766 3639 9818
rect 3691 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 13308 9818
rect 13360 9766 13372 9818
rect 13424 9766 13436 9818
rect 13488 9766 13500 9818
rect 13552 9766 15824 9818
rect 1104 9744 15824 9766
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 5166 9704 5172 9716
rect 2924 9676 5028 9704
rect 5127 9676 5172 9704
rect 2924 9664 2930 9676
rect 2133 9639 2191 9645
rect 2133 9605 2145 9639
rect 2179 9636 2191 9639
rect 2682 9636 2688 9648
rect 2179 9608 2688 9636
rect 2179 9605 2191 9608
rect 2133 9599 2191 9605
rect 2682 9596 2688 9608
rect 2740 9596 2746 9648
rect 2961 9639 3019 9645
rect 2961 9605 2973 9639
rect 3007 9636 3019 9639
rect 3694 9636 3700 9648
rect 3007 9608 3700 9636
rect 3007 9605 3019 9608
rect 2961 9599 3019 9605
rect 3694 9596 3700 9608
rect 3752 9596 3758 9648
rect 5000 9636 5028 9676
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 11698 9704 11704 9716
rect 5316 9676 9260 9704
rect 5316 9664 5322 9676
rect 8665 9639 8723 9645
rect 5000 9608 5273 9636
rect 2314 9568 2320 9580
rect 1596 9540 2320 9568
rect 1596 9509 1624 9540
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 2590 9568 2596 9580
rect 2551 9540 2596 9568
rect 2590 9528 2596 9540
rect 2648 9528 2654 9580
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9568 2835 9571
rect 3605 9571 3663 9577
rect 2823 9540 3556 9568
rect 2823 9537 2835 9540
rect 2777 9531 2835 9537
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9469 1639 9503
rect 1581 9463 1639 9469
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9500 1915 9503
rect 2866 9500 2872 9512
rect 1903 9472 2872 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 3234 9500 3240 9512
rect 3016 9472 3240 9500
rect 3016 9460 3022 9472
rect 3234 9460 3240 9472
rect 3292 9460 3298 9512
rect 2498 9432 2504 9444
rect 2459 9404 2504 9432
rect 2498 9392 2504 9404
rect 2556 9392 2562 9444
rect 3528 9432 3556 9540
rect 3605 9537 3617 9571
rect 3651 9568 3663 9571
rect 3651 9540 3924 9568
rect 3651 9537 3663 9540
rect 3605 9531 3663 9537
rect 3786 9500 3792 9512
rect 3747 9472 3792 9500
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 3896 9500 3924 9540
rect 4982 9528 4988 9580
rect 5040 9528 5046 9580
rect 5245 9568 5273 9608
rect 8665 9605 8677 9639
rect 8711 9636 8723 9639
rect 9122 9636 9128 9648
rect 8711 9608 9128 9636
rect 8711 9605 8723 9608
rect 8665 9599 8723 9605
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 9232 9636 9260 9676
rect 10980 9676 11704 9704
rect 9861 9639 9919 9645
rect 9861 9636 9873 9639
rect 9232 9608 9873 9636
rect 9861 9605 9873 9608
rect 9907 9605 9919 9639
rect 9861 9599 9919 9605
rect 10226 9596 10232 9648
rect 10284 9596 10290 9648
rect 10686 9596 10692 9648
rect 10744 9636 10750 9648
rect 10980 9636 11008 9676
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 12584 9676 14136 9704
rect 12584 9664 12590 9676
rect 12253 9639 12311 9645
rect 12253 9636 12265 9639
rect 10744 9608 11008 9636
rect 11532 9608 12265 9636
rect 10744 9596 10750 9608
rect 6822 9568 6828 9580
rect 5245 9540 5396 9568
rect 6783 9540 6828 9568
rect 4522 9500 4528 9512
rect 3896 9472 4528 9500
rect 4522 9460 4528 9472
rect 4580 9460 4586 9512
rect 4798 9460 4804 9512
rect 4856 9500 4862 9512
rect 5000 9500 5028 9528
rect 5261 9503 5319 9509
rect 5261 9500 5273 9503
rect 4856 9472 5273 9500
rect 4856 9460 4862 9472
rect 5261 9469 5273 9472
rect 5307 9469 5319 9503
rect 5261 9463 5319 9469
rect 3878 9432 3884 9444
rect 3528 9404 3884 9432
rect 3878 9392 3884 9404
rect 3936 9432 3942 9444
rect 4056 9435 4114 9441
rect 4056 9432 4068 9435
rect 3936 9404 4068 9432
rect 3936 9392 3942 9404
rect 4056 9401 4068 9404
rect 4102 9432 4114 9435
rect 5368 9432 5396 9540
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 8110 9528 8116 9580
rect 8168 9568 8174 9580
rect 8754 9568 8760 9580
rect 8168 9540 8760 9568
rect 8168 9528 8174 9540
rect 8754 9528 8760 9540
rect 8812 9528 8818 9580
rect 8938 9528 8944 9580
rect 8996 9568 9002 9580
rect 9217 9571 9275 9577
rect 9217 9568 9229 9571
rect 8996 9540 9229 9568
rect 8996 9528 9002 9540
rect 9217 9537 9229 9540
rect 9263 9537 9275 9571
rect 9217 9531 9275 9537
rect 9398 9528 9404 9580
rect 9456 9568 9462 9580
rect 10244 9568 10272 9596
rect 10410 9568 10416 9580
rect 9456 9540 10272 9568
rect 10371 9540 10416 9568
rect 9456 9528 9462 9540
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 10502 9528 10508 9580
rect 10560 9568 10566 9580
rect 11238 9568 11244 9580
rect 10560 9540 11244 9568
rect 10560 9528 10566 9540
rect 11238 9528 11244 9540
rect 11296 9528 11302 9580
rect 11532 9577 11560 9608
rect 12253 9605 12265 9608
rect 12299 9605 12311 9639
rect 12253 9599 12311 9605
rect 12437 9639 12495 9645
rect 12437 9605 12449 9639
rect 12483 9636 12495 9639
rect 13446 9636 13452 9648
rect 12483 9608 13452 9636
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 13446 9596 13452 9608
rect 13504 9596 13510 9648
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9537 11759 9571
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 11701 9531 11759 9537
rect 11992 9540 13001 9568
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 9125 9503 9183 9509
rect 5868 9472 9076 9500
rect 5868 9460 5874 9472
rect 5528 9435 5586 9441
rect 5528 9432 5540 9435
rect 4102 9404 5212 9432
rect 5368 9404 5540 9432
rect 4102 9401 4114 9404
rect 4056 9395 4114 9401
rect 3326 9364 3332 9376
rect 3287 9336 3332 9364
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 3421 9367 3479 9373
rect 3421 9333 3433 9367
rect 3467 9364 3479 9367
rect 4982 9364 4988 9376
rect 3467 9336 4988 9364
rect 3467 9333 3479 9336
rect 3421 9327 3479 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5184 9364 5212 9404
rect 5528 9401 5540 9404
rect 5574 9432 5586 9435
rect 5626 9432 5632 9444
rect 5574 9404 5632 9432
rect 5574 9401 5586 9404
rect 5528 9395 5586 9401
rect 5626 9392 5632 9404
rect 5684 9392 5690 9444
rect 5718 9392 5724 9444
rect 5776 9432 5782 9444
rect 6270 9432 6276 9444
rect 5776 9404 6276 9432
rect 5776 9392 5782 9404
rect 6270 9392 6276 9404
rect 6328 9432 6334 9444
rect 7070 9435 7128 9441
rect 7070 9432 7082 9435
rect 6328 9404 7082 9432
rect 6328 9392 6334 9404
rect 7070 9401 7082 9404
rect 7116 9401 7128 9435
rect 7070 9395 7128 9401
rect 7190 9392 7196 9444
rect 7248 9432 7254 9444
rect 8386 9432 8392 9444
rect 7248 9404 8392 9432
rect 7248 9392 7254 9404
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 9048 9432 9076 9472
rect 9125 9469 9137 9503
rect 9171 9500 9183 9503
rect 9674 9500 9680 9512
rect 9171 9472 9680 9500
rect 9171 9469 9183 9472
rect 9125 9463 9183 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 10229 9503 10287 9509
rect 10229 9469 10241 9503
rect 10275 9500 10287 9503
rect 11146 9500 11152 9512
rect 10275 9472 11152 9500
rect 10275 9469 10287 9472
rect 10229 9463 10287 9469
rect 11146 9460 11152 9472
rect 11204 9460 11210 9512
rect 11422 9500 11428 9512
rect 11383 9472 11428 9500
rect 11422 9460 11428 9472
rect 11480 9460 11486 9512
rect 11716 9500 11744 9531
rect 11670 9472 11744 9500
rect 11670 9444 11698 9472
rect 9048 9404 9168 9432
rect 6641 9367 6699 9373
rect 6641 9364 6653 9367
rect 5184 9336 6653 9364
rect 6641 9333 6653 9336
rect 6687 9333 6699 9367
rect 6641 9327 6699 9333
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 7432 9336 8217 9364
rect 7432 9324 7438 9336
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 9030 9364 9036 9376
rect 8991 9336 9036 9364
rect 8205 9327 8263 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9140 9364 9168 9404
rect 9766 9392 9772 9444
rect 9824 9432 9830 9444
rect 10778 9432 10784 9444
rect 9824 9404 10784 9432
rect 9824 9392 9830 9404
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 11670 9432 11704 9444
rect 10980 9404 11704 9432
rect 9674 9364 9680 9376
rect 9140 9336 9680 9364
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 10226 9324 10232 9376
rect 10284 9364 10290 9376
rect 10321 9367 10379 9373
rect 10321 9364 10333 9367
rect 10284 9336 10333 9364
rect 10284 9324 10290 9336
rect 10321 9333 10333 9336
rect 10367 9333 10379 9367
rect 10321 9327 10379 9333
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 10980 9364 11008 9404
rect 11698 9392 11704 9404
rect 11756 9432 11762 9444
rect 11992 9432 12020 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 13906 9568 13912 9580
rect 12989 9531 13047 9537
rect 13096 9540 13912 9568
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9469 12311 9503
rect 13096 9500 13124 9540
rect 13906 9528 13912 9540
rect 13964 9528 13970 9580
rect 14108 9577 14136 9676
rect 14642 9664 14648 9716
rect 14700 9704 14706 9716
rect 15194 9704 15200 9716
rect 14700 9676 15200 9704
rect 14700 9664 14706 9676
rect 15194 9664 15200 9676
rect 15252 9664 15258 9716
rect 14093 9571 14151 9577
rect 14093 9537 14105 9571
rect 14139 9537 14151 9571
rect 14093 9531 14151 9537
rect 14185 9571 14243 9577
rect 14185 9537 14197 9571
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 12253 9463 12311 9469
rect 12452 9472 13124 9500
rect 11756 9404 11803 9432
rect 11900 9404 12020 9432
rect 12268 9432 12296 9463
rect 12452 9432 12480 9472
rect 13170 9460 13176 9512
rect 13228 9500 13234 9512
rect 14200 9500 14228 9531
rect 13228 9472 13676 9500
rect 13228 9460 13234 9472
rect 12268 9404 12480 9432
rect 12805 9435 12863 9441
rect 11756 9392 11762 9404
rect 10560 9336 11008 9364
rect 11057 9367 11115 9373
rect 10560 9324 10566 9336
rect 11057 9333 11069 9367
rect 11103 9364 11115 9367
rect 11330 9364 11336 9376
rect 11103 9336 11336 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 11422 9324 11428 9376
rect 11480 9364 11486 9376
rect 11900 9364 11928 9404
rect 12805 9401 12817 9435
rect 12851 9432 12863 9435
rect 13262 9432 13268 9444
rect 12851 9404 13268 9432
rect 12851 9401 12863 9404
rect 12805 9395 12863 9401
rect 13262 9392 13268 9404
rect 13320 9392 13326 9444
rect 11480 9336 11928 9364
rect 11480 9324 11486 9336
rect 11974 9324 11980 9376
rect 12032 9364 12038 9376
rect 12250 9364 12256 9376
rect 12032 9336 12256 9364
rect 12032 9324 12038 9336
rect 12250 9324 12256 9336
rect 12308 9324 12314 9376
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 13170 9364 13176 9376
rect 12943 9336 13176 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 13648 9373 13676 9472
rect 14108 9472 14228 9500
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 14108 9432 14136 9472
rect 14366 9460 14372 9512
rect 14424 9500 14430 9512
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 14424 9472 14841 9500
rect 14424 9460 14430 9472
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 13780 9404 14136 9432
rect 13780 9392 13786 9404
rect 13633 9367 13691 9373
rect 13633 9333 13645 9367
rect 13679 9333 13691 9367
rect 13633 9327 13691 9333
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14001 9367 14059 9373
rect 14001 9364 14013 9367
rect 13964 9336 14013 9364
rect 13964 9324 13970 9336
rect 14001 9333 14013 9336
rect 14047 9333 14059 9367
rect 15010 9364 15016 9376
rect 14971 9336 15016 9364
rect 14001 9327 14059 9333
rect 15010 9324 15016 9336
rect 15068 9324 15074 9376
rect 1104 9274 15824 9296
rect 1104 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 6104 9274
rect 6156 9222 10843 9274
rect 10895 9222 10907 9274
rect 10959 9222 10971 9274
rect 11023 9222 11035 9274
rect 11087 9222 15824 9274
rect 1104 9200 15824 9222
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 2832 9132 2877 9160
rect 2832 9120 2838 9132
rect 3326 9120 3332 9172
rect 3384 9160 3390 9172
rect 4157 9163 4215 9169
rect 4157 9160 4169 9163
rect 3384 9132 4169 9160
rect 3384 9120 3390 9132
rect 4157 9129 4169 9132
rect 4203 9129 4215 9163
rect 4157 9123 4215 9129
rect 4249 9163 4307 9169
rect 4249 9129 4261 9163
rect 4295 9129 4307 9163
rect 7466 9160 7472 9172
rect 4249 9123 4307 9129
rect 4356 9132 7472 9160
rect 2682 9052 2688 9104
rect 2740 9092 2746 9104
rect 4264 9092 4292 9123
rect 2740 9064 4292 9092
rect 2740 9052 2746 9064
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 9024 2007 9027
rect 2498 9024 2504 9036
rect 1995 8996 2504 9024
rect 1995 8993 2007 8996
rect 1949 8987 2007 8993
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 3145 9027 3203 9033
rect 2832 8996 2912 9024
rect 2832 8984 2838 8996
rect 937 8959 995 8965
rect 937 8925 949 8959
rect 983 8956 995 8959
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 983 8928 2053 8956
rect 983 8925 995 8928
rect 937 8919 995 8925
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8925 2283 8959
rect 2884 8956 2912 8996
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 3694 9024 3700 9036
rect 3191 8996 3700 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 3694 8984 3700 8996
rect 3752 8984 3758 9036
rect 4157 9027 4215 9033
rect 4157 8993 4169 9027
rect 4203 9024 4215 9027
rect 4356 9024 4384 9132
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 7558 9120 7564 9172
rect 7616 9160 7622 9172
rect 7745 9163 7803 9169
rect 7745 9160 7757 9163
rect 7616 9132 7757 9160
rect 7616 9120 7622 9132
rect 7745 9129 7757 9132
rect 7791 9129 7803 9163
rect 7745 9123 7803 9129
rect 8018 9120 8024 9172
rect 8076 9160 8082 9172
rect 10045 9163 10103 9169
rect 8076 9132 9996 9160
rect 8076 9120 8082 9132
rect 4614 9092 4620 9104
rect 4575 9064 4620 9092
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 5166 9052 5172 9104
rect 5224 9092 5230 9104
rect 5224 9064 8616 9092
rect 5224 9052 5230 9064
rect 4203 8996 4384 9024
rect 4203 8993 4215 8996
rect 4157 8987 4215 8993
rect 4430 8984 4436 9036
rect 4488 9024 4494 9036
rect 4709 9027 4767 9033
rect 4709 9024 4721 9027
rect 4488 8996 4721 9024
rect 4488 8984 4494 8996
rect 4709 8993 4721 8996
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 5074 8984 5080 9036
rect 5132 9024 5138 9036
rect 5905 9027 5963 9033
rect 5905 9024 5917 9027
rect 5132 8996 5917 9024
rect 5132 8984 5138 8996
rect 5905 8993 5917 8996
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 7653 9027 7711 9033
rect 7653 8993 7665 9027
rect 7699 9024 7711 9027
rect 7834 9024 7840 9036
rect 7699 8996 7840 9024
rect 7699 8993 7711 8996
rect 7653 8987 7711 8993
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 8110 9024 8116 9036
rect 8071 8996 8116 9024
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 8205 9027 8263 9033
rect 8205 8993 8217 9027
rect 8251 9024 8263 9027
rect 8478 9024 8484 9036
rect 8251 8996 8484 9024
rect 8251 8993 8263 8996
rect 8205 8987 8263 8993
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 2884 8928 3249 8956
rect 2225 8919 2283 8925
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 4893 8959 4951 8965
rect 3467 8928 4752 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 1946 8820 1952 8832
rect 1627 8792 1952 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 2240 8820 2268 8919
rect 3786 8848 3792 8900
rect 3844 8888 3850 8900
rect 4430 8888 4436 8900
rect 3844 8860 4436 8888
rect 3844 8848 3850 8860
rect 4430 8848 4436 8860
rect 4488 8848 4494 8900
rect 4522 8820 4528 8832
rect 2240 8792 4528 8820
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 4724 8820 4752 8928
rect 4893 8925 4905 8959
rect 4939 8956 4951 8959
rect 7006 8956 7012 8968
rect 4939 8928 7012 8956
rect 4939 8925 4951 8928
rect 4893 8919 4951 8925
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 8220 8956 8248 8987
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 8588 9033 8616 9064
rect 8754 9052 8760 9104
rect 8812 9092 8818 9104
rect 9766 9092 9772 9104
rect 8812 9064 9772 9092
rect 8812 9052 8818 9064
rect 9766 9052 9772 9064
rect 9824 9052 9830 9104
rect 8573 9027 8631 9033
rect 8573 8993 8585 9027
rect 8619 8993 8631 9027
rect 9968 9024 9996 9132
rect 10045 9129 10057 9163
rect 10091 9160 10103 9163
rect 10318 9160 10324 9172
rect 10091 9132 10324 9160
rect 10091 9129 10103 9132
rect 10045 9123 10103 9129
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 11330 9160 11336 9172
rect 11291 9132 11336 9160
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 12069 9163 12127 9169
rect 12069 9129 12081 9163
rect 12115 9129 12127 9163
rect 12069 9123 12127 9129
rect 12437 9163 12495 9169
rect 12437 9129 12449 9163
rect 12483 9160 12495 9163
rect 12802 9160 12808 9172
rect 12483 9132 12808 9160
rect 12483 9129 12495 9132
rect 12437 9123 12495 9129
rect 10134 9092 10140 9104
rect 10095 9064 10140 9092
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 10778 9052 10784 9104
rect 10836 9092 10842 9104
rect 12084 9092 12112 9123
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 13170 9120 13176 9172
rect 13228 9160 13234 9172
rect 13265 9163 13323 9169
rect 13265 9160 13277 9163
rect 13228 9132 13277 9160
rect 13228 9120 13234 9132
rect 13265 9129 13277 9132
rect 13311 9129 13323 9163
rect 13265 9123 13323 9129
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 13725 9163 13783 9169
rect 13725 9160 13737 9163
rect 13504 9132 13737 9160
rect 13504 9120 13510 9132
rect 13725 9129 13737 9132
rect 13771 9129 13783 9163
rect 13725 9123 13783 9129
rect 12250 9092 12256 9104
rect 10836 9064 11376 9092
rect 12084 9064 12256 9092
rect 10836 9052 10842 9064
rect 11238 9024 11244 9036
rect 9968 8996 10916 9024
rect 11199 8996 11244 9024
rect 8573 8987 8631 8993
rect 8386 8956 8392 8968
rect 7800 8928 8248 8956
rect 8347 8928 8392 8956
rect 7800 8916 7806 8928
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8925 8815 8959
rect 8757 8919 8815 8925
rect 4798 8848 4804 8900
rect 4856 8888 4862 8900
rect 8772 8888 8800 8919
rect 10042 8916 10048 8968
rect 10100 8956 10106 8968
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 10100 8928 10241 8956
rect 10100 8916 10106 8928
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 10888 8956 10916 8996
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 11348 9024 11376 9064
rect 12250 9052 12256 9064
rect 12308 9052 12314 9104
rect 15194 9092 15200 9104
rect 12360 9064 15200 9092
rect 12360 9024 12388 9064
rect 15194 9052 15200 9064
rect 15252 9052 15258 9104
rect 12526 9024 12532 9036
rect 11348 8996 12388 9024
rect 12487 8996 12532 9024
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 13170 8984 13176 9036
rect 13228 9024 13234 9036
rect 13633 9027 13691 9033
rect 13633 9024 13645 9027
rect 13228 8996 13645 9024
rect 13228 8984 13234 8996
rect 13633 8993 13645 8996
rect 13679 8993 13691 9027
rect 13633 8987 13691 8993
rect 14274 8984 14280 9036
rect 14332 9024 14338 9036
rect 14461 9027 14519 9033
rect 14461 9024 14473 9027
rect 14332 8996 14473 9024
rect 14332 8984 14338 8996
rect 14461 8993 14473 8996
rect 14507 8993 14519 9027
rect 14461 8987 14519 8993
rect 11330 8956 11336 8968
rect 10888 8928 11336 8956
rect 10229 8919 10287 8925
rect 11330 8916 11336 8928
rect 11388 8956 11394 8968
rect 11425 8959 11483 8965
rect 11425 8956 11437 8959
rect 11388 8928 11437 8956
rect 11388 8916 11394 8928
rect 11425 8925 11437 8928
rect 11471 8925 11483 8959
rect 12621 8959 12679 8965
rect 12621 8956 12633 8959
rect 11425 8919 11483 8925
rect 11532 8928 12633 8956
rect 10873 8891 10931 8897
rect 10873 8888 10885 8891
rect 4856 8860 8800 8888
rect 8864 8860 10885 8888
rect 4856 8848 4862 8860
rect 7374 8820 7380 8832
rect 4724 8792 7380 8820
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 7466 8780 7472 8832
rect 7524 8820 7530 8832
rect 8864 8820 8892 8860
rect 10873 8857 10885 8860
rect 10919 8857 10931 8891
rect 10873 8851 10931 8857
rect 10962 8848 10968 8900
rect 11020 8888 11026 8900
rect 11532 8888 11560 8928
rect 12621 8925 12633 8928
rect 12667 8925 12679 8959
rect 12621 8919 12679 8925
rect 13817 8959 13875 8965
rect 13817 8925 13829 8959
rect 13863 8925 13875 8959
rect 13817 8919 13875 8925
rect 13722 8888 13728 8900
rect 11020 8860 11560 8888
rect 12636 8860 13728 8888
rect 11020 8848 11026 8860
rect 12636 8832 12664 8860
rect 13722 8848 13728 8860
rect 13780 8888 13786 8900
rect 13832 8888 13860 8919
rect 13780 8860 13860 8888
rect 13780 8848 13786 8860
rect 9674 8820 9680 8832
rect 7524 8792 8892 8820
rect 9635 8792 9680 8820
rect 7524 8780 7530 8792
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 11054 8820 11060 8832
rect 9824 8792 11060 8820
rect 9824 8780 9830 8792
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 12618 8780 12624 8832
rect 12676 8780 12682 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 14645 8823 14703 8829
rect 14645 8820 14657 8823
rect 13872 8792 14657 8820
rect 13872 8780 13878 8792
rect 14645 8789 14657 8792
rect 14691 8789 14703 8823
rect 14645 8783 14703 8789
rect 1104 8730 15824 8752
rect 1104 8678 3447 8730
rect 3499 8678 3511 8730
rect 3563 8678 3575 8730
rect 3627 8678 3639 8730
rect 3691 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 13308 8730
rect 13360 8678 13372 8730
rect 13424 8678 13436 8730
rect 13488 8678 13500 8730
rect 13552 8678 15824 8730
rect 1104 8656 15824 8678
rect 9582 8616 9588 8628
rect 4080 8588 9588 8616
rect 3697 8551 3755 8557
rect 3697 8548 3709 8551
rect 1596 8520 3709 8548
rect 1596 8421 1624 8520
rect 3697 8517 3709 8520
rect 3743 8517 3755 8551
rect 3697 8511 3755 8517
rect 2958 8480 2964 8492
rect 2919 8452 2964 8480
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 3510 8480 3516 8492
rect 3191 8452 3516 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8381 1639 8415
rect 1581 8375 1639 8381
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 3786 8412 3792 8424
rect 2915 8384 3792 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 3786 8372 3792 8384
rect 3844 8372 3850 8424
rect 1210 8304 1216 8356
rect 1268 8344 1274 8356
rect 1857 8347 1915 8353
rect 1857 8344 1869 8347
rect 1268 8316 1869 8344
rect 1268 8304 1274 8316
rect 1857 8313 1869 8316
rect 1903 8313 1915 8347
rect 3326 8344 3332 8356
rect 1857 8307 1915 8313
rect 2240 8316 3332 8344
rect 1302 8236 1308 8288
rect 1360 8276 1366 8288
rect 2240 8276 2268 8316
rect 3326 8304 3332 8316
rect 3384 8344 3390 8356
rect 3970 8344 3976 8356
rect 3384 8316 3976 8344
rect 3384 8304 3390 8316
rect 3970 8304 3976 8316
rect 4028 8304 4034 8356
rect 4080 8353 4108 8588
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 9858 8576 9864 8628
rect 9916 8616 9922 8628
rect 10318 8616 10324 8628
rect 9916 8588 10324 8616
rect 9916 8576 9922 8588
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 11054 8616 11060 8628
rect 11015 8588 11060 8616
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 12437 8619 12495 8625
rect 12437 8616 12449 8619
rect 11296 8588 12449 8616
rect 11296 8576 11302 8588
rect 12437 8585 12449 8588
rect 12483 8585 12495 8619
rect 12437 8579 12495 8585
rect 13078 8576 13084 8628
rect 13136 8616 13142 8628
rect 13633 8619 13691 8625
rect 13633 8616 13645 8619
rect 13136 8588 13645 8616
rect 13136 8576 13142 8588
rect 13633 8585 13645 8588
rect 13679 8585 13691 8619
rect 13633 8579 13691 8585
rect 6270 8548 6276 8560
rect 6231 8520 6276 8548
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 7834 8508 7840 8560
rect 7892 8548 7898 8560
rect 8202 8548 8208 8560
rect 7892 8520 8208 8548
rect 7892 8508 7898 8520
rect 8202 8508 8208 8520
rect 8260 8548 8266 8560
rect 8938 8548 8944 8560
rect 8260 8520 8944 8548
rect 8260 8508 8266 8520
rect 8938 8508 8944 8520
rect 8996 8508 9002 8560
rect 10962 8548 10968 8560
rect 9232 8520 10968 8548
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4798 8480 4804 8492
rect 4387 8452 4804 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 9232 8489 9260 8520
rect 10962 8508 10968 8520
rect 11020 8508 11026 8560
rect 11606 8508 11612 8560
rect 11664 8548 11670 8560
rect 12894 8548 12900 8560
rect 11664 8520 12900 8548
rect 11664 8508 11670 8520
rect 12894 8508 12900 8520
rect 12952 8548 12958 8560
rect 14458 8548 14464 8560
rect 12952 8520 13032 8548
rect 12952 8508 12958 8520
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 7984 8452 9229 8480
rect 7984 8440 7990 8452
rect 9217 8449 9229 8452
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 9766 8440 9772 8492
rect 9824 8480 9830 8492
rect 10042 8480 10048 8492
rect 9824 8452 10048 8480
rect 9824 8440 9830 8452
rect 10042 8440 10048 8452
rect 10100 8480 10106 8492
rect 10413 8483 10471 8489
rect 10413 8480 10425 8483
rect 10100 8452 10425 8480
rect 10100 8440 10106 8452
rect 10413 8449 10425 8452
rect 10459 8449 10471 8483
rect 10413 8443 10471 8449
rect 11330 8440 11336 8492
rect 11388 8480 11394 8492
rect 13004 8489 13032 8520
rect 13740 8520 14464 8548
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11388 8452 11713 8480
rect 11388 8440 11394 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 12989 8483 13047 8489
rect 12989 8449 13001 8483
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 13740 8424 13768 8520
rect 14458 8508 14464 8520
rect 14516 8508 14522 8560
rect 14277 8483 14335 8489
rect 14277 8480 14289 8483
rect 14200 8452 14289 8480
rect 14200 8424 14228 8452
rect 14277 8449 14289 8452
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 4706 8372 4712 8424
rect 4764 8412 4770 8424
rect 5166 8421 5172 8424
rect 4893 8415 4951 8421
rect 4893 8412 4905 8415
rect 4764 8384 4905 8412
rect 4764 8372 4770 8384
rect 4893 8381 4905 8384
rect 4939 8381 4951 8415
rect 5160 8412 5172 8421
rect 5127 8384 5172 8412
rect 4893 8375 4951 8381
rect 5160 8375 5172 8384
rect 5166 8372 5172 8375
rect 5224 8372 5230 8424
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 11517 8415 11575 8421
rect 11517 8412 11529 8415
rect 6932 8384 11529 8412
rect 4065 8347 4123 8353
rect 4065 8313 4077 8347
rect 4111 8313 4123 8347
rect 4065 8307 4123 8313
rect 4157 8347 4215 8353
rect 4157 8313 4169 8347
rect 4203 8344 4215 8347
rect 6362 8344 6368 8356
rect 4203 8316 6368 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 6362 8304 6368 8316
rect 6420 8304 6426 8356
rect 6932 8344 6960 8384
rect 11517 8381 11529 8384
rect 11563 8381 11575 8415
rect 13722 8412 13728 8424
rect 11517 8375 11575 8381
rect 12820 8384 13728 8412
rect 6840 8316 6960 8344
rect 1360 8248 2268 8276
rect 1360 8236 1366 8248
rect 2314 8236 2320 8288
rect 2372 8276 2378 8288
rect 2501 8279 2559 8285
rect 2501 8276 2513 8279
rect 2372 8248 2513 8276
rect 2372 8236 2378 8248
rect 2501 8245 2513 8248
rect 2547 8245 2559 8279
rect 2501 8239 2559 8245
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 6840 8276 6868 8316
rect 7006 8304 7012 8356
rect 7064 8353 7070 8356
rect 7064 8347 7128 8353
rect 7064 8313 7082 8347
rect 7116 8344 7128 8347
rect 7926 8344 7932 8356
rect 7116 8316 7932 8344
rect 7116 8313 7128 8316
rect 7064 8307 7128 8313
rect 7064 8304 7070 8307
rect 7926 8304 7932 8316
rect 7984 8304 7990 8356
rect 8754 8344 8760 8356
rect 8220 8316 8760 8344
rect 2648 8248 6868 8276
rect 2648 8236 2654 8248
rect 7834 8236 7840 8288
rect 7892 8276 7898 8288
rect 8220 8285 8248 8316
rect 8754 8304 8760 8316
rect 8812 8304 8818 8356
rect 10321 8347 10379 8353
rect 10321 8313 10333 8347
rect 10367 8344 10379 8347
rect 12820 8344 12848 8384
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 13906 8372 13912 8424
rect 13964 8412 13970 8424
rect 14093 8415 14151 8421
rect 14093 8412 14105 8415
rect 13964 8384 14105 8412
rect 13964 8372 13970 8384
rect 14093 8381 14105 8384
rect 14139 8381 14151 8415
rect 14093 8375 14151 8381
rect 14182 8372 14188 8424
rect 14240 8372 14246 8424
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 14829 8415 14887 8421
rect 14829 8412 14841 8415
rect 14608 8384 14841 8412
rect 14608 8372 14614 8384
rect 14829 8381 14841 8384
rect 14875 8381 14887 8415
rect 14829 8375 14887 8381
rect 10367 8316 12848 8344
rect 12897 8347 12955 8353
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 12897 8313 12909 8347
rect 12943 8344 12955 8347
rect 12943 8316 13032 8344
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 7892 8248 8217 8276
rect 7892 8236 7898 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 8205 8239 8263 8245
rect 8294 8236 8300 8288
rect 8352 8276 8358 8288
rect 8665 8279 8723 8285
rect 8665 8276 8677 8279
rect 8352 8248 8677 8276
rect 8352 8236 8358 8248
rect 8665 8245 8677 8248
rect 8711 8245 8723 8279
rect 9030 8276 9036 8288
rect 8991 8248 9036 8276
rect 8665 8239 8723 8245
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 9490 8276 9496 8288
rect 9180 8248 9496 8276
rect 9180 8236 9186 8248
rect 9490 8236 9496 8248
rect 9548 8236 9554 8288
rect 9858 8276 9864 8288
rect 9819 8248 9864 8276
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 10226 8276 10232 8288
rect 10187 8248 10232 8276
rect 10226 8236 10232 8248
rect 10284 8236 10290 8288
rect 11330 8236 11336 8288
rect 11388 8276 11394 8288
rect 11425 8279 11483 8285
rect 11425 8276 11437 8279
rect 11388 8248 11437 8276
rect 11388 8236 11394 8248
rect 11425 8245 11437 8248
rect 11471 8245 11483 8279
rect 11425 8239 11483 8245
rect 11514 8236 11520 8288
rect 11572 8276 11578 8288
rect 11790 8276 11796 8288
rect 11572 8248 11796 8276
rect 11572 8236 11578 8248
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 12802 8276 12808 8288
rect 12763 8248 12808 8276
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 13004 8276 13032 8316
rect 13078 8304 13084 8356
rect 13136 8344 13142 8356
rect 14001 8347 14059 8353
rect 14001 8344 14013 8347
rect 13136 8316 14013 8344
rect 13136 8304 13142 8316
rect 14001 8313 14013 8316
rect 14047 8313 14059 8347
rect 14274 8344 14280 8356
rect 14001 8307 14059 8313
rect 14108 8316 14280 8344
rect 14108 8276 14136 8316
rect 14274 8304 14280 8316
rect 14332 8304 14338 8356
rect 13004 8248 14136 8276
rect 15013 8279 15071 8285
rect 15013 8245 15025 8279
rect 15059 8276 15071 8279
rect 15562 8276 15568 8288
rect 15059 8248 15568 8276
rect 15059 8245 15071 8248
rect 15013 8239 15071 8245
rect 15562 8236 15568 8248
rect 15620 8236 15626 8288
rect 1104 8186 15824 8208
rect 1104 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 6104 8186
rect 6156 8134 10843 8186
rect 10895 8134 10907 8186
rect 10959 8134 10971 8186
rect 11023 8134 11035 8186
rect 11087 8134 15824 8186
rect 1104 8112 15824 8134
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2682 8072 2688 8084
rect 1995 8044 2688 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 5166 8032 5172 8084
rect 5224 8072 5230 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 5224 8044 7297 8072
rect 5224 8032 5230 8044
rect 7285 8041 7297 8044
rect 7331 8072 7343 8075
rect 8018 8072 8024 8084
rect 7331 8044 8024 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 9125 8075 9183 8081
rect 9125 8041 9137 8075
rect 9171 8072 9183 8075
rect 9398 8072 9404 8084
rect 9171 8044 9404 8072
rect 9171 8041 9183 8044
rect 9125 8035 9183 8041
rect 9398 8032 9404 8044
rect 9456 8032 9462 8084
rect 9582 8032 9588 8084
rect 9640 8072 9646 8084
rect 9677 8075 9735 8081
rect 9677 8072 9689 8075
rect 9640 8044 9689 8072
rect 9640 8032 9646 8044
rect 9677 8041 9689 8044
rect 9723 8041 9735 8075
rect 9677 8035 9735 8041
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 9916 8044 10149 8072
rect 9916 8032 9922 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8041 10931 8075
rect 10873 8035 10931 8041
rect 3145 8007 3203 8013
rect 3145 7973 3157 8007
rect 3191 8004 3203 8007
rect 10888 8004 10916 8035
rect 11146 8032 11152 8084
rect 11204 8032 11210 8084
rect 11330 8032 11336 8084
rect 11388 8072 11394 8084
rect 12069 8075 12127 8081
rect 12069 8072 12081 8075
rect 11388 8044 12081 8072
rect 11388 8032 11394 8044
rect 12069 8041 12081 8044
rect 12115 8041 12127 8075
rect 12069 8035 12127 8041
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12492 8044 12537 8072
rect 12492 8032 12498 8044
rect 3191 7976 10916 8004
rect 3191 7973 3203 7976
rect 3145 7967 3203 7973
rect 2682 7896 2688 7948
rect 2740 7936 2746 7948
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 2740 7908 4077 7936
rect 2740 7896 2746 7908
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 4065 7899 4123 7905
rect 4332 7939 4390 7945
rect 4332 7905 4344 7939
rect 4378 7936 4390 7939
rect 5626 7936 5632 7948
rect 4378 7908 5632 7936
rect 4378 7905 4390 7908
rect 4332 7899 4390 7905
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 5994 7896 6000 7948
rect 6052 7936 6058 7948
rect 6161 7939 6219 7945
rect 6161 7936 6173 7939
rect 6052 7908 6173 7936
rect 6052 7896 6058 7908
rect 6161 7905 6173 7908
rect 6207 7936 6219 7939
rect 7834 7936 7840 7948
rect 6207 7908 7840 7936
rect 6207 7905 6219 7908
rect 6161 7899 6219 7905
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 8012 7939 8070 7945
rect 8012 7905 8024 7939
rect 8058 7936 8070 7939
rect 10045 7939 10103 7945
rect 8058 7908 9444 7936
rect 8058 7905 8070 7908
rect 8012 7899 8070 7905
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7837 2099 7871
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2041 7831 2099 7837
rect 2056 7800 2084 7831
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 3234 7868 3240 7880
rect 3195 7840 3240 7868
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7868 3479 7871
rect 3786 7868 3792 7880
rect 3467 7840 3792 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 3970 7800 3976 7812
rect 2056 7772 3976 7800
rect 3970 7760 3976 7772
rect 4028 7760 4034 7812
rect 5368 7772 5948 7800
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 2590 7732 2596 7744
rect 1627 7704 2596 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 2590 7692 2596 7704
rect 2648 7692 2654 7744
rect 2777 7735 2835 7741
rect 2777 7701 2789 7735
rect 2823 7732 2835 7735
rect 5368 7732 5396 7772
rect 2823 7704 5396 7732
rect 2823 7701 2835 7704
rect 2777 7695 2835 7701
rect 5442 7692 5448 7744
rect 5500 7732 5506 7744
rect 5920 7732 5948 7772
rect 7190 7732 7196 7744
rect 5500 7704 5545 7732
rect 5920 7704 7196 7732
rect 5500 7692 5506 7704
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 7760 7732 7788 7831
rect 9214 7800 9220 7812
rect 8680 7772 9220 7800
rect 8680 7744 8708 7772
rect 9214 7760 9220 7772
rect 9272 7760 9278 7812
rect 9416 7800 9444 7908
rect 10045 7905 10057 7939
rect 10091 7936 10103 7939
rect 10778 7936 10784 7948
rect 10091 7908 10784 7936
rect 10091 7905 10103 7908
rect 10045 7899 10103 7905
rect 10778 7896 10784 7908
rect 10836 7896 10842 7948
rect 11164 7936 11192 8032
rect 11241 8007 11299 8013
rect 11241 7973 11253 8007
rect 11287 8004 11299 8007
rect 11790 8004 11796 8016
rect 11287 7976 11796 8004
rect 11287 7973 11299 7976
rect 11241 7967 11299 7973
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 11164 7908 12020 7936
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 9548 7840 10241 7868
rect 9548 7828 9554 7840
rect 10229 7837 10241 7840
rect 10275 7868 10287 7871
rect 11054 7868 11060 7880
rect 10275 7840 11060 7868
rect 10275 7837 10287 7840
rect 10229 7831 10287 7837
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 11204 7840 11345 7868
rect 11204 7828 11210 7840
rect 11333 7837 11345 7840
rect 11379 7837 11391 7871
rect 11514 7868 11520 7880
rect 11475 7840 11520 7868
rect 11333 7831 11391 7837
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 9416 7772 9996 7800
rect 8662 7732 8668 7744
rect 7524 7704 8668 7732
rect 7524 7692 7530 7704
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 9030 7692 9036 7744
rect 9088 7732 9094 7744
rect 9858 7732 9864 7744
rect 9088 7704 9864 7732
rect 9088 7692 9094 7704
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 9968 7732 9996 7772
rect 10042 7760 10048 7812
rect 10100 7800 10106 7812
rect 10962 7800 10968 7812
rect 10100 7772 10968 7800
rect 10100 7760 10106 7772
rect 10962 7760 10968 7772
rect 11020 7760 11026 7812
rect 11992 7800 12020 7908
rect 12250 7896 12256 7948
rect 12308 7936 12314 7948
rect 12308 7908 12388 7936
rect 12308 7896 12314 7908
rect 12360 7868 12388 7908
rect 13170 7896 13176 7948
rect 13228 7936 13234 7948
rect 13633 7939 13691 7945
rect 13633 7936 13645 7939
rect 13228 7908 13645 7936
rect 13228 7896 13234 7908
rect 13633 7905 13645 7908
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 13998 7896 14004 7948
rect 14056 7936 14062 7948
rect 14461 7939 14519 7945
rect 14461 7936 14473 7939
rect 14056 7908 14473 7936
rect 14056 7896 14062 7908
rect 14461 7905 14473 7908
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12360 7840 12541 7868
rect 12529 7837 12541 7840
rect 12575 7837 12587 7871
rect 12529 7831 12587 7837
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7868 12771 7871
rect 12894 7868 12900 7880
rect 12759 7840 12900 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 13909 7871 13967 7877
rect 13909 7837 13921 7871
rect 13955 7868 13967 7871
rect 14182 7868 14188 7880
rect 13955 7840 14188 7868
rect 13955 7837 13967 7840
rect 13909 7831 13967 7837
rect 12250 7800 12256 7812
rect 11992 7772 12256 7800
rect 12250 7760 12256 7772
rect 12308 7760 12314 7812
rect 13262 7800 13268 7812
rect 13223 7772 13268 7800
rect 13262 7760 13268 7772
rect 13320 7760 13326 7812
rect 11238 7732 11244 7744
rect 9968 7704 11244 7732
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 12066 7692 12072 7744
rect 12124 7732 12130 7744
rect 13740 7732 13768 7831
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 13998 7760 14004 7812
rect 14056 7800 14062 7812
rect 14918 7800 14924 7812
rect 14056 7772 14924 7800
rect 14056 7760 14062 7772
rect 14918 7760 14924 7772
rect 14976 7760 14982 7812
rect 14642 7732 14648 7744
rect 12124 7704 13768 7732
rect 14603 7704 14648 7732
rect 12124 7692 12130 7704
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 1104 7642 15824 7664
rect 1104 7590 3447 7642
rect 3499 7590 3511 7642
rect 3563 7590 3575 7642
rect 3627 7590 3639 7642
rect 3691 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 13308 7642
rect 13360 7590 13372 7642
rect 13424 7590 13436 7642
rect 13488 7590 13500 7642
rect 13552 7590 15824 7642
rect 1104 7568 15824 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 1857 7531 1915 7537
rect 1857 7528 1869 7531
rect 1820 7500 1869 7528
rect 1820 7488 1826 7500
rect 1857 7497 1869 7500
rect 1903 7497 1915 7531
rect 1857 7491 1915 7497
rect 2222 7488 2228 7540
rect 2280 7528 2286 7540
rect 5994 7528 6000 7540
rect 2280 7500 6000 7528
rect 2280 7488 2286 7500
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 7190 7488 7196 7540
rect 7248 7528 7254 7540
rect 14182 7528 14188 7540
rect 7248 7500 11008 7528
rect 7248 7488 7254 7500
rect 4154 7420 4160 7472
rect 4212 7460 4218 7472
rect 4433 7463 4491 7469
rect 4433 7460 4445 7463
rect 4212 7432 4445 7460
rect 4212 7420 4218 7432
rect 4433 7429 4445 7432
rect 4479 7460 4491 7463
rect 4890 7460 4896 7472
rect 4479 7432 4896 7460
rect 4479 7429 4491 7432
rect 4433 7423 4491 7429
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 7926 7420 7932 7472
rect 7984 7460 7990 7472
rect 8205 7463 8263 7469
rect 8205 7460 8217 7463
rect 7984 7432 8217 7460
rect 7984 7420 7990 7432
rect 8205 7429 8217 7432
rect 8251 7429 8263 7463
rect 8205 7423 8263 7429
rect 9858 7420 9864 7472
rect 9916 7460 9922 7472
rect 10505 7463 10563 7469
rect 10505 7460 10517 7463
rect 9916 7432 10517 7460
rect 9916 7420 9922 7432
rect 10505 7429 10517 7432
rect 10551 7429 10563 7463
rect 10505 7423 10563 7429
rect 2314 7392 2320 7404
rect 2275 7364 2320 7392
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 2547 7364 3188 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7293 3111 7327
rect 3053 7287 3111 7293
rect 2314 7216 2320 7268
rect 2372 7256 2378 7268
rect 2682 7256 2688 7268
rect 2372 7228 2688 7256
rect 2372 7216 2378 7228
rect 2682 7216 2688 7228
rect 2740 7256 2746 7268
rect 3068 7256 3096 7287
rect 2740 7228 3096 7256
rect 2740 7216 2746 7228
rect 2225 7191 2283 7197
rect 2225 7157 2237 7191
rect 2271 7188 2283 7191
rect 2498 7188 2504 7200
rect 2271 7160 2504 7188
rect 2271 7157 2283 7160
rect 2225 7151 2283 7157
rect 2498 7148 2504 7160
rect 2556 7148 2562 7200
rect 3160 7188 3188 7364
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6328 7364 6960 7392
rect 6328 7352 6334 7364
rect 4706 7284 4712 7336
rect 4764 7324 4770 7336
rect 4893 7327 4951 7333
rect 4893 7324 4905 7327
rect 4764 7296 4905 7324
rect 4764 7284 4770 7296
rect 4893 7293 4905 7296
rect 4939 7293 4951 7327
rect 5718 7324 5724 7336
rect 4893 7287 4951 7293
rect 5092 7296 5724 7324
rect 3320 7259 3378 7265
rect 3320 7225 3332 7259
rect 3366 7256 3378 7259
rect 5092 7256 5120 7296
rect 5718 7284 5724 7296
rect 5776 7284 5782 7336
rect 5902 7284 5908 7336
rect 5960 7324 5966 7336
rect 6822 7324 6828 7336
rect 5960 7296 6828 7324
rect 5960 7284 5966 7296
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 6932 7324 6960 7364
rect 8110 7352 8116 7404
rect 8168 7392 8174 7404
rect 10594 7392 10600 7404
rect 8168 7364 8800 7392
rect 8168 7352 8174 7364
rect 7081 7327 7139 7333
rect 7081 7324 7093 7327
rect 6932 7296 7093 7324
rect 7081 7293 7093 7296
rect 7127 7293 7139 7327
rect 8662 7324 8668 7336
rect 8623 7296 8668 7324
rect 7081 7287 7139 7293
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 8772 7324 8800 7364
rect 10244 7364 10600 7392
rect 8921 7327 8979 7333
rect 8921 7324 8933 7327
rect 8772 7296 8933 7324
rect 8921 7293 8933 7296
rect 8967 7324 8979 7327
rect 10244 7324 10272 7364
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 10980 7401 11008 7500
rect 11164 7500 14188 7528
rect 11164 7472 11192 7500
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 11146 7420 11152 7472
rect 11204 7420 11210 7472
rect 11256 7432 14228 7460
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 11054 7352 11060 7404
rect 11112 7392 11118 7404
rect 11112 7364 11157 7392
rect 11112 7352 11118 7364
rect 10873 7327 10931 7333
rect 10873 7324 10885 7327
rect 8967 7296 10272 7324
rect 10336 7296 10885 7324
rect 8967 7293 8979 7296
rect 8921 7287 8979 7293
rect 3366 7228 5120 7256
rect 5160 7259 5218 7265
rect 3366 7225 3378 7228
rect 3320 7219 3378 7225
rect 5160 7225 5172 7259
rect 5206 7256 5218 7259
rect 8386 7256 8392 7268
rect 5206 7228 8392 7256
rect 5206 7225 5218 7228
rect 5160 7219 5218 7225
rect 8386 7216 8392 7228
rect 8444 7216 8450 7268
rect 9674 7216 9680 7268
rect 9732 7256 9738 7268
rect 10336 7256 10364 7296
rect 10873 7293 10885 7296
rect 10919 7293 10931 7327
rect 10873 7287 10931 7293
rect 9732 7228 10364 7256
rect 9732 7216 9738 7228
rect 10594 7216 10600 7268
rect 10652 7256 10658 7268
rect 11256 7256 11284 7432
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12768 7364 12909 7392
rect 12768 7352 12774 7364
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13630 7392 13636 7404
rect 13127 7364 13636 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 11701 7327 11759 7333
rect 11701 7293 11713 7327
rect 11747 7324 11759 7327
rect 12802 7324 12808 7336
rect 11747 7296 12808 7324
rect 11747 7293 11759 7296
rect 11701 7287 11759 7293
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 13096 7256 13124 7355
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 14200 7401 14228 7432
rect 14185 7395 14243 7401
rect 14185 7361 14197 7395
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 13780 7296 14841 7324
rect 13780 7284 13786 7296
rect 14829 7293 14841 7296
rect 14875 7293 14887 7327
rect 14829 7287 14887 7293
rect 10652 7228 11284 7256
rect 12084 7228 13124 7256
rect 14093 7259 14151 7265
rect 10652 7216 10658 7228
rect 5626 7188 5632 7200
rect 3160 7160 5632 7188
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 5718 7148 5724 7200
rect 5776 7188 5782 7200
rect 6270 7188 6276 7200
rect 5776 7160 6276 7188
rect 5776 7148 5782 7160
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 6822 7148 6828 7200
rect 6880 7188 6886 7200
rect 7466 7188 7472 7200
rect 6880 7160 7472 7188
rect 6880 7148 6886 7160
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 7558 7148 7564 7200
rect 7616 7188 7622 7200
rect 10045 7191 10103 7197
rect 10045 7188 10057 7191
rect 7616 7160 10057 7188
rect 7616 7148 7622 7160
rect 10045 7157 10057 7160
rect 10091 7188 10103 7191
rect 12084 7188 12112 7228
rect 14093 7225 14105 7259
rect 14139 7256 14151 7259
rect 14918 7256 14924 7268
rect 14139 7228 14924 7256
rect 14139 7225 14151 7228
rect 14093 7219 14151 7225
rect 14918 7216 14924 7228
rect 14976 7216 14982 7268
rect 10091 7160 12112 7188
rect 12437 7191 12495 7197
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 12437 7157 12449 7191
rect 12483 7188 12495 7191
rect 12526 7188 12532 7200
rect 12483 7160 12532 7188
rect 12483 7157 12495 7160
rect 12437 7151 12495 7157
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 12802 7188 12808 7200
rect 12763 7160 12808 7188
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 13630 7188 13636 7200
rect 13591 7160 13636 7188
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 14001 7191 14059 7197
rect 14001 7157 14013 7191
rect 14047 7188 14059 7191
rect 14550 7188 14556 7200
rect 14047 7160 14556 7188
rect 14047 7157 14059 7160
rect 14001 7151 14059 7157
rect 14550 7148 14556 7160
rect 14608 7148 14614 7200
rect 15010 7188 15016 7200
rect 14971 7160 15016 7188
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 1104 7098 15824 7120
rect 1104 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 6104 7098
rect 6156 7046 10843 7098
rect 10895 7046 10907 7098
rect 10959 7046 10971 7098
rect 11023 7046 11035 7098
rect 11087 7046 15824 7098
rect 1104 7024 15824 7046
rect 2682 6944 2688 6996
rect 2740 6984 2746 6996
rect 2774 6984 2780 6996
rect 2740 6956 2780 6984
rect 2740 6944 2746 6956
rect 2774 6944 2780 6956
rect 2832 6944 2838 6996
rect 3786 6944 3792 6996
rect 3844 6984 3850 6996
rect 6270 6984 6276 6996
rect 3844 6956 6276 6984
rect 3844 6944 3850 6956
rect 6270 6944 6276 6956
rect 6328 6944 6334 6996
rect 7101 6987 7159 6993
rect 7101 6953 7113 6987
rect 7147 6984 7159 6987
rect 7147 6956 8340 6984
rect 7147 6953 7159 6956
rect 7101 6947 7159 6953
rect 4890 6876 4896 6928
rect 4948 6916 4954 6928
rect 5350 6916 5356 6928
rect 4948 6888 5356 6916
rect 4948 6876 4954 6888
rect 5350 6876 5356 6888
rect 5408 6876 5414 6928
rect 6288 6916 6316 6944
rect 8312 6916 8340 6956
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8444 6956 8953 6984
rect 8444 6944 8450 6956
rect 8941 6953 8953 6956
rect 8987 6984 8999 6987
rect 9490 6984 9496 6996
rect 8987 6956 9496 6984
rect 8987 6953 8999 6956
rect 8941 6947 8999 6953
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 10042 6984 10048 6996
rect 10003 6956 10048 6984
rect 10042 6944 10048 6956
rect 10100 6984 10106 6996
rect 10100 6956 10732 6984
rect 10100 6944 10106 6956
rect 10594 6916 10600 6928
rect 6288 6888 7236 6916
rect 8312 6888 10600 6916
rect 1302 6808 1308 6860
rect 1360 6848 1366 6860
rect 1397 6851 1455 6857
rect 1397 6848 1409 6851
rect 1360 6820 1409 6848
rect 1360 6808 1366 6820
rect 1397 6817 1409 6820
rect 1443 6817 1455 6851
rect 1397 6811 1455 6817
rect 2400 6851 2458 6857
rect 2400 6817 2412 6851
rect 2446 6848 2458 6851
rect 4154 6848 4160 6860
rect 2446 6820 4160 6848
rect 2446 6817 2458 6820
rect 2400 6811 2458 6817
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6817 4307 6851
rect 5074 6848 5080 6860
rect 5035 6820 5080 6848
rect 4249 6811 4307 6817
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 4264 6780 4292 6811
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 5988 6851 6046 6857
rect 5988 6817 6000 6851
rect 6034 6848 6046 6851
rect 6034 6820 7144 6848
rect 6034 6817 6046 6820
rect 5988 6811 6046 6817
rect 4028 6752 4292 6780
rect 4028 6740 4034 6752
rect 4706 6740 4712 6792
rect 4764 6780 4770 6792
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 4764 6752 5733 6780
rect 4764 6740 4770 6752
rect 5721 6749 5733 6752
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 3513 6715 3571 6721
rect 3513 6681 3525 6715
rect 3559 6712 3571 6715
rect 5534 6712 5540 6724
rect 3559 6684 5540 6712
rect 3559 6681 3571 6684
rect 3513 6675 3571 6681
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 1394 6604 1400 6656
rect 1452 6644 1458 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1452 6616 1593 6644
rect 1452 6604 1458 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 2498 6604 2504 6656
rect 2556 6644 2562 6656
rect 5258 6644 5264 6656
rect 2556 6616 5264 6644
rect 2556 6604 2562 6616
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 7116 6644 7144 6820
rect 7208 6780 7236 6888
rect 9140 6860 9168 6888
rect 10594 6876 10600 6888
rect 10652 6876 10658 6928
rect 10704 6916 10732 6956
rect 11146 6944 11152 6996
rect 11204 6984 11210 6996
rect 12069 6987 12127 6993
rect 12069 6984 12081 6987
rect 11204 6956 12081 6984
rect 11204 6944 11210 6956
rect 12069 6953 12081 6956
rect 12115 6953 12127 6987
rect 12069 6947 12127 6953
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 13265 6987 13323 6993
rect 13265 6984 13277 6987
rect 12860 6956 13277 6984
rect 12860 6944 12866 6956
rect 13265 6953 13277 6956
rect 13311 6953 13323 6987
rect 13265 6947 13323 6953
rect 11241 6919 11299 6925
rect 11241 6916 11253 6919
rect 10704 6888 11253 6916
rect 11241 6885 11253 6888
rect 11287 6885 11299 6919
rect 11241 6879 11299 6885
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 7834 6857 7840 6860
rect 7561 6851 7619 6857
rect 7561 6848 7573 6851
rect 7524 6820 7573 6848
rect 7524 6808 7530 6820
rect 7561 6817 7573 6820
rect 7607 6817 7619 6851
rect 7817 6851 7840 6857
rect 7817 6848 7829 6851
rect 7561 6811 7619 6817
rect 7668 6820 7829 6848
rect 7668 6780 7696 6820
rect 7817 6817 7829 6820
rect 7817 6811 7840 6817
rect 7834 6808 7840 6811
rect 7892 6808 7898 6860
rect 9122 6808 9128 6860
rect 9180 6808 9186 6860
rect 11256 6848 11284 6879
rect 11514 6876 11520 6928
rect 11572 6916 11578 6928
rect 12437 6919 12495 6925
rect 12437 6916 12449 6919
rect 11572 6888 12449 6916
rect 11572 6876 11578 6888
rect 12437 6885 12449 6888
rect 12483 6885 12495 6919
rect 13633 6919 13691 6925
rect 12437 6879 12495 6885
rect 12728 6888 13400 6916
rect 11698 6848 11704 6860
rect 10152 6820 10640 6848
rect 11256 6820 11704 6848
rect 7208 6752 7696 6780
rect 10042 6740 10048 6792
rect 10100 6780 10106 6792
rect 10152 6789 10180 6820
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 10100 6752 10149 6780
rect 10100 6740 10106 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10318 6780 10324 6792
rect 10279 6752 10324 6780
rect 10137 6743 10195 6749
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 10612 6780 10640 6820
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 12728 6848 12756 6888
rect 12544 6820 12756 6848
rect 13372 6848 13400 6888
rect 13633 6885 13645 6919
rect 13679 6916 13691 6919
rect 13722 6916 13728 6928
rect 13679 6888 13728 6916
rect 13679 6885 13691 6888
rect 13633 6879 13691 6885
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 14366 6848 14372 6860
rect 13372 6820 14372 6848
rect 11146 6780 11152 6792
rect 10612 6752 11152 6780
rect 11146 6740 11152 6752
rect 11204 6780 11210 6792
rect 11333 6783 11391 6789
rect 11333 6780 11345 6783
rect 11204 6752 11345 6780
rect 11204 6740 11210 6752
rect 11333 6749 11345 6752
rect 11379 6749 11391 6783
rect 11333 6743 11391 6749
rect 11422 6740 11428 6792
rect 11480 6780 11486 6792
rect 12544 6789 12572 6820
rect 14366 6808 14372 6820
rect 14424 6808 14430 6860
rect 14461 6851 14519 6857
rect 14461 6817 14473 6851
rect 14507 6848 14519 6851
rect 14642 6848 14648 6860
rect 14507 6820 14648 6848
rect 14507 6817 14519 6820
rect 14461 6811 14519 6817
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 12529 6783 12587 6789
rect 11480 6752 11573 6780
rect 11480 6740 11486 6752
rect 12529 6749 12541 6783
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 12621 6783 12679 6789
rect 12621 6749 12633 6783
rect 12667 6749 12679 6783
rect 12621 6743 12679 6749
rect 11440 6712 11468 6740
rect 12636 6712 12664 6743
rect 12710 6740 12716 6792
rect 12768 6780 12774 6792
rect 13725 6783 13783 6789
rect 13725 6780 13737 6783
rect 12768 6752 13737 6780
rect 12768 6740 12774 6752
rect 13725 6749 13737 6752
rect 13771 6749 13783 6783
rect 13725 6743 13783 6749
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6749 13967 6783
rect 13909 6743 13967 6749
rect 9508 6684 11468 6712
rect 11532 6684 12664 6712
rect 7926 6644 7932 6656
rect 7116 6616 7932 6644
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8202 6604 8208 6656
rect 8260 6644 8266 6656
rect 9508 6644 9536 6684
rect 9674 6644 9680 6656
rect 8260 6616 9536 6644
rect 9635 6616 9680 6644
rect 8260 6604 8266 6616
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 10873 6647 10931 6653
rect 10873 6644 10885 6647
rect 10192 6616 10885 6644
rect 10192 6604 10198 6616
rect 10873 6613 10885 6616
rect 10919 6613 10931 6647
rect 10873 6607 10931 6613
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 11532 6644 11560 6684
rect 13814 6672 13820 6724
rect 13872 6712 13878 6724
rect 13924 6712 13952 6743
rect 13872 6684 13952 6712
rect 13872 6672 13878 6684
rect 11020 6616 11560 6644
rect 11020 6604 11026 6616
rect 11698 6604 11704 6656
rect 11756 6644 11762 6656
rect 14645 6647 14703 6653
rect 14645 6644 14657 6647
rect 11756 6616 14657 6644
rect 11756 6604 11762 6616
rect 14645 6613 14657 6616
rect 14691 6613 14703 6647
rect 14645 6607 14703 6613
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 1857 6443 1915 6449
rect 1857 6409 1869 6443
rect 1903 6440 1915 6443
rect 3234 6440 3240 6452
rect 1903 6412 3240 6440
rect 1903 6409 1915 6412
rect 1857 6403 1915 6409
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 4433 6443 4491 6449
rect 4433 6409 4445 6443
rect 4479 6440 4491 6443
rect 4614 6440 4620 6452
rect 4479 6412 4620 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 5166 6440 5172 6452
rect 4724 6412 5172 6440
rect 4724 6372 4752 6412
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 5258 6400 5264 6452
rect 5316 6440 5322 6452
rect 10042 6440 10048 6452
rect 5316 6412 10048 6440
rect 5316 6400 5322 6412
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 15013 6443 15071 6449
rect 15013 6440 15025 6443
rect 10192 6412 15025 6440
rect 10192 6400 10198 6412
rect 15013 6409 15025 6412
rect 15059 6409 15071 6443
rect 15013 6403 15071 6409
rect 6270 6372 6276 6384
rect 4632 6344 4752 6372
rect 6231 6344 6276 6372
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6304 2559 6307
rect 2547 6276 3188 6304
rect 2547 6273 2559 6276
rect 2501 6267 2559 6273
rect 2130 6196 2136 6248
rect 2188 6236 2194 6248
rect 3053 6239 3111 6245
rect 3053 6236 3065 6239
rect 2188 6208 3065 6236
rect 2188 6196 2194 6208
rect 3053 6205 3065 6208
rect 3099 6205 3111 6239
rect 3160 6236 3188 6276
rect 4632 6236 4660 6344
rect 6270 6332 6276 6344
rect 6328 6332 6334 6384
rect 7926 6332 7932 6384
rect 7984 6372 7990 6384
rect 8205 6375 8263 6381
rect 8205 6372 8217 6375
rect 7984 6344 8217 6372
rect 7984 6332 7990 6344
rect 8205 6341 8217 6344
rect 8251 6341 8263 6375
rect 8205 6335 8263 6341
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 4893 6307 4951 6313
rect 4893 6304 4905 6307
rect 4764 6276 4905 6304
rect 4764 6264 4770 6276
rect 4893 6273 4905 6276
rect 4939 6273 4951 6307
rect 6822 6304 6828 6316
rect 6783 6276 6828 6304
rect 4893 6267 4951 6273
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 8220 6304 8248 6335
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 11698 6372 11704 6384
rect 9824 6344 11704 6372
rect 9824 6332 9830 6344
rect 11698 6332 11704 6344
rect 11756 6332 11762 6384
rect 13446 6332 13452 6384
rect 13504 6372 13510 6384
rect 13633 6375 13691 6381
rect 13633 6372 13645 6375
rect 13504 6344 13645 6372
rect 13504 6332 13510 6344
rect 13633 6341 13645 6344
rect 13679 6341 13691 6375
rect 13633 6335 13691 6341
rect 8220 6276 8800 6304
rect 7558 6236 7564 6248
rect 3160 6208 4660 6236
rect 5092 6208 7564 6236
rect 3053 6199 3111 6205
rect 2222 6168 2228 6180
rect 2183 6140 2228 6168
rect 2222 6128 2228 6140
rect 2280 6128 2286 6180
rect 2317 6103 2375 6109
rect 2317 6069 2329 6103
rect 2363 6100 2375 6103
rect 2682 6100 2688 6112
rect 2363 6072 2688 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 2682 6060 2688 6072
rect 2740 6060 2746 6112
rect 3068 6100 3096 6199
rect 3320 6171 3378 6177
rect 3320 6137 3332 6171
rect 3366 6168 3378 6171
rect 5092 6168 5120 6208
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 8662 6236 8668 6248
rect 8623 6208 8668 6236
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 8772 6236 8800 6276
rect 9950 6264 9956 6316
rect 10008 6304 10014 6316
rect 10965 6307 11023 6313
rect 10965 6304 10977 6307
rect 10008 6276 10977 6304
rect 10008 6264 10014 6276
rect 10965 6273 10977 6276
rect 11011 6273 11023 6307
rect 11146 6304 11152 6316
rect 11107 6276 11152 6304
rect 10965 6267 11023 6273
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12342 6304 12348 6316
rect 12216 6276 12348 6304
rect 12216 6264 12222 6276
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 12526 6264 12532 6316
rect 12584 6304 12590 6316
rect 12894 6304 12900 6316
rect 12584 6276 12900 6304
rect 12584 6264 12590 6276
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 12989 6307 13047 6313
rect 12989 6273 13001 6307
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 9214 6236 9220 6248
rect 8772 6208 9220 6236
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 10134 6236 10140 6248
rect 9548 6208 10140 6236
rect 9548 6196 9554 6208
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 10744 6208 10885 6236
rect 10744 6196 10750 6208
rect 10873 6205 10885 6208
rect 10919 6205 10931 6239
rect 13004 6236 13032 6267
rect 13998 6264 14004 6316
rect 14056 6304 14062 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 14056 6276 14105 6304
rect 14056 6264 14062 6276
rect 14093 6273 14105 6276
rect 14139 6273 14151 6307
rect 14274 6304 14280 6316
rect 14235 6276 14280 6304
rect 14093 6267 14151 6273
rect 14274 6264 14280 6276
rect 14332 6264 14338 6316
rect 10873 6199 10931 6205
rect 10980 6208 13032 6236
rect 14829 6239 14887 6245
rect 5166 6177 5172 6180
rect 3366 6140 5120 6168
rect 3366 6137 3378 6140
rect 3320 6131 3378 6137
rect 5160 6131 5172 6177
rect 5224 6168 5230 6180
rect 7092 6171 7150 6177
rect 5224 6140 5260 6168
rect 5166 6128 5172 6131
rect 5224 6128 5230 6140
rect 7092 6137 7104 6171
rect 7138 6168 7150 6171
rect 7926 6168 7932 6180
rect 7138 6140 7932 6168
rect 7138 6137 7150 6140
rect 7092 6131 7150 6137
rect 7926 6128 7932 6140
rect 7984 6128 7990 6180
rect 8110 6128 8116 6180
rect 8168 6168 8174 6180
rect 8754 6168 8760 6180
rect 8168 6140 8760 6168
rect 8168 6128 8174 6140
rect 8754 6128 8760 6140
rect 8812 6168 8818 6180
rect 8910 6171 8968 6177
rect 8910 6168 8922 6171
rect 8812 6140 8922 6168
rect 8812 6128 8818 6140
rect 8910 6137 8922 6140
rect 8956 6137 8968 6171
rect 8910 6131 8968 6137
rect 9030 6128 9036 6180
rect 9088 6168 9094 6180
rect 9088 6140 10548 6168
rect 9088 6128 9094 6140
rect 4706 6100 4712 6112
rect 3068 6072 4712 6100
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 5626 6060 5632 6112
rect 5684 6100 5690 6112
rect 10520 6109 10548 6140
rect 10594 6128 10600 6180
rect 10652 6168 10658 6180
rect 10980 6168 11008 6208
rect 14829 6205 14841 6239
rect 14875 6236 14887 6239
rect 15654 6236 15660 6248
rect 14875 6208 15660 6236
rect 14875 6205 14887 6208
rect 14829 6199 14887 6205
rect 15654 6196 15660 6208
rect 15712 6196 15718 6248
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 10652 6140 11008 6168
rect 12728 6140 12817 6168
rect 10652 6128 10658 6140
rect 12728 6112 12756 6140
rect 12805 6137 12817 6140
rect 12851 6137 12863 6171
rect 12805 6131 12863 6137
rect 10045 6103 10103 6109
rect 10045 6100 10057 6103
rect 5684 6072 10057 6100
rect 5684 6060 5690 6072
rect 10045 6069 10057 6072
rect 10091 6069 10103 6103
rect 10045 6063 10103 6069
rect 10505 6103 10563 6109
rect 10505 6069 10517 6103
rect 10551 6069 10563 6103
rect 11698 6100 11704 6112
rect 11659 6072 11704 6100
rect 10505 6063 10563 6069
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12492 6072 12537 6100
rect 12492 6060 12498 6072
rect 12710 6060 12716 6112
rect 12768 6060 12774 6112
rect 12894 6100 12900 6112
rect 12855 6072 12900 6100
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13998 6100 14004 6112
rect 13959 6072 14004 6100
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 2406 5856 2412 5908
rect 2464 5896 2470 5908
rect 3513 5899 3571 5905
rect 3513 5896 3525 5899
rect 2464 5868 3525 5896
rect 2464 5856 2470 5868
rect 3513 5865 3525 5868
rect 3559 5865 3571 5899
rect 3513 5859 3571 5865
rect 4617 5899 4675 5905
rect 4617 5865 4629 5899
rect 4663 5896 4675 5899
rect 8570 5896 8576 5908
rect 4663 5868 8576 5896
rect 4663 5865 4675 5868
rect 4617 5859 4675 5865
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5896 9183 5899
rect 9306 5896 9312 5908
rect 9171 5868 9312 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 10594 5896 10600 5908
rect 9508 5868 10600 5896
rect 2222 5828 2228 5840
rect 1412 5800 2228 5828
rect 1412 5769 1440 5800
rect 2222 5788 2228 5800
rect 2280 5788 2286 5840
rect 4709 5831 4767 5837
rect 4709 5797 4721 5831
rect 4755 5828 4767 5831
rect 7006 5828 7012 5840
rect 4755 5800 7012 5828
rect 4755 5797 4767 5800
rect 4709 5791 4767 5797
rect 7006 5788 7012 5800
rect 7064 5788 7070 5840
rect 7282 5788 7288 5840
rect 7340 5828 7346 5840
rect 9398 5828 9404 5840
rect 7340 5800 9404 5828
rect 7340 5788 7346 5800
rect 9398 5788 9404 5800
rect 9456 5788 9462 5840
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5729 1455 5763
rect 2130 5760 2136 5772
rect 2091 5732 2136 5760
rect 1397 5723 1455 5729
rect 2130 5720 2136 5732
rect 2188 5720 2194 5772
rect 2400 5763 2458 5769
rect 2400 5729 2412 5763
rect 2446 5760 2458 5763
rect 4154 5760 4160 5772
rect 2446 5732 4160 5760
rect 2446 5729 2458 5732
rect 2400 5723 2458 5729
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5760 5503 5763
rect 5534 5760 5540 5772
rect 5491 5732 5540 5760
rect 5491 5729 5503 5732
rect 5445 5723 5503 5729
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 5718 5769 5724 5772
rect 5712 5760 5724 5769
rect 5679 5732 5724 5760
rect 5712 5723 5724 5732
rect 5718 5720 5724 5723
rect 5776 5720 5782 5772
rect 7552 5763 7610 5769
rect 7552 5729 7564 5763
rect 7598 5760 7610 5763
rect 8110 5760 8116 5772
rect 7598 5732 8116 5760
rect 7598 5729 7610 5732
rect 7552 5723 7610 5729
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 8938 5720 8944 5772
rect 8996 5760 9002 5772
rect 9309 5763 9367 5769
rect 9309 5760 9321 5763
rect 8996 5732 9321 5760
rect 8996 5720 9002 5732
rect 9309 5729 9321 5732
rect 9355 5729 9367 5763
rect 9508 5760 9536 5868
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 11057 5899 11115 5905
rect 11057 5865 11069 5899
rect 11103 5896 11115 5899
rect 11238 5896 11244 5908
rect 11103 5868 11244 5896
rect 11103 5865 11115 5868
rect 11057 5859 11115 5865
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 12710 5896 12716 5908
rect 12671 5868 12716 5896
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 13081 5899 13139 5905
rect 13081 5896 13093 5899
rect 13044 5868 13093 5896
rect 13044 5856 13050 5868
rect 13081 5865 13093 5868
rect 13127 5865 13139 5899
rect 13081 5859 13139 5865
rect 13173 5899 13231 5905
rect 13173 5865 13185 5899
rect 13219 5896 13231 5899
rect 14182 5896 14188 5908
rect 13219 5868 14188 5896
rect 13219 5865 13231 5868
rect 13173 5859 13231 5865
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 10042 5788 10048 5840
rect 10100 5828 10106 5840
rect 12434 5828 12440 5840
rect 10100 5800 12440 5828
rect 10100 5788 10106 5800
rect 12434 5788 12440 5800
rect 12492 5788 12498 5840
rect 9309 5723 9367 5729
rect 9416 5732 9536 5760
rect 4062 5692 4068 5704
rect 3160 5664 4068 5692
rect 1578 5556 1584 5568
rect 1539 5528 1584 5556
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 2774 5516 2780 5568
rect 2832 5556 2838 5568
rect 3160 5556 3188 5664
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5692 4951 5695
rect 5166 5692 5172 5704
rect 4939 5664 5172 5692
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 6822 5652 6828 5704
rect 6880 5692 6886 5704
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 6880 5664 7297 5692
rect 6880 5652 6886 5664
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 9416 5692 9444 5732
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 9766 5760 9772 5772
rect 9640 5732 9772 5760
rect 9640 5720 9646 5732
rect 9766 5720 9772 5732
rect 9824 5760 9830 5772
rect 9933 5763 9991 5769
rect 9933 5760 9945 5763
rect 9824 5732 9945 5760
rect 9824 5720 9830 5732
rect 9933 5729 9945 5732
rect 9979 5729 9991 5763
rect 9933 5723 9991 5729
rect 10226 5720 10232 5772
rect 10284 5760 10290 5772
rect 10778 5760 10784 5772
rect 10284 5732 10784 5760
rect 10284 5720 10290 5732
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 11882 5760 11888 5772
rect 11795 5732 11888 5760
rect 11882 5720 11888 5732
rect 11940 5760 11946 5772
rect 13630 5760 13636 5772
rect 11940 5732 13636 5760
rect 11940 5720 11946 5732
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 14182 5720 14188 5772
rect 14240 5760 14246 5772
rect 14277 5763 14335 5769
rect 14277 5760 14289 5763
rect 14240 5732 14289 5760
rect 14240 5720 14246 5732
rect 14277 5729 14289 5732
rect 14323 5729 14335 5763
rect 14277 5723 14335 5729
rect 8812 5664 9444 5692
rect 9677 5695 9735 5701
rect 8812 5652 8818 5664
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 11977 5695 12035 5701
rect 11977 5692 11989 5695
rect 9677 5655 9735 5661
rect 11072 5664 11989 5692
rect 8570 5584 8576 5636
rect 8628 5624 8634 5636
rect 8938 5624 8944 5636
rect 8628 5596 8944 5624
rect 8628 5584 8634 5596
rect 8938 5584 8944 5596
rect 8996 5584 9002 5636
rect 2832 5528 3188 5556
rect 2832 5516 2838 5528
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 4249 5559 4307 5565
rect 4249 5556 4261 5559
rect 4120 5528 4261 5556
rect 4120 5516 4126 5528
rect 4249 5525 4261 5528
rect 4295 5525 4307 5559
rect 4249 5519 4307 5525
rect 4338 5516 4344 5568
rect 4396 5556 4402 5568
rect 4614 5556 4620 5568
rect 4396 5528 4620 5556
rect 4396 5516 4402 5528
rect 4614 5516 4620 5528
rect 4672 5516 4678 5568
rect 5442 5516 5448 5568
rect 5500 5556 5506 5568
rect 6825 5559 6883 5565
rect 6825 5556 6837 5559
rect 5500 5528 6837 5556
rect 5500 5516 5506 5528
rect 6825 5525 6837 5528
rect 6871 5525 6883 5559
rect 8662 5556 8668 5568
rect 8623 5528 8668 5556
rect 6825 5519 6883 5525
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 9692 5556 9720 5655
rect 9858 5556 9864 5568
rect 9692 5528 9864 5556
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 10042 5516 10048 5568
rect 10100 5556 10106 5568
rect 10410 5556 10416 5568
rect 10100 5528 10416 5556
rect 10100 5516 10106 5528
rect 10410 5516 10416 5528
rect 10468 5556 10474 5568
rect 11072 5556 11100 5664
rect 11977 5661 11989 5664
rect 12023 5661 12035 5695
rect 11977 5655 12035 5661
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5661 12127 5695
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 12069 5655 12127 5661
rect 12912 5664 13369 5692
rect 11146 5584 11152 5636
rect 11204 5624 11210 5636
rect 12084 5624 12112 5655
rect 11204 5596 12112 5624
rect 11204 5584 11210 5596
rect 11514 5556 11520 5568
rect 10468 5528 11100 5556
rect 11475 5528 11520 5556
rect 10468 5516 10474 5528
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 12802 5516 12808 5568
rect 12860 5556 12866 5568
rect 12912 5556 12940 5664
rect 13357 5661 13369 5664
rect 13403 5692 13415 5695
rect 13538 5692 13544 5704
rect 13403 5664 13544 5692
rect 13403 5661 13415 5664
rect 13357 5655 13415 5661
rect 13538 5652 13544 5664
rect 13596 5652 13602 5704
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 12986 5584 12992 5636
rect 13044 5624 13050 5636
rect 14384 5624 14412 5655
rect 14458 5652 14464 5704
rect 14516 5692 14522 5704
rect 14516 5664 14561 5692
rect 14516 5652 14522 5664
rect 13044 5596 14412 5624
rect 13044 5584 13050 5596
rect 13906 5556 13912 5568
rect 12860 5528 12940 5556
rect 13867 5528 13912 5556
rect 12860 5516 12866 5528
rect 13906 5516 13912 5528
rect 13964 5516 13970 5568
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 6822 5352 6828 5364
rect 2240 5324 6828 5352
rect 2240 5157 2268 5324
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7926 5312 7932 5364
rect 7984 5352 7990 5364
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 7984 5324 8217 5352
rect 7984 5312 7990 5324
rect 8205 5321 8217 5324
rect 8251 5352 8263 5355
rect 8251 5324 11008 5352
rect 8251 5321 8263 5324
rect 8205 5315 8263 5321
rect 4154 5244 4160 5296
rect 4212 5284 4218 5296
rect 4433 5287 4491 5293
rect 4433 5284 4445 5287
rect 4212 5256 4445 5284
rect 4212 5244 4218 5256
rect 4433 5253 4445 5256
rect 4479 5284 4491 5287
rect 4890 5284 4896 5296
rect 4479 5256 4896 5284
rect 4479 5253 4491 5256
rect 4433 5247 4491 5253
rect 4890 5244 4896 5256
rect 4948 5244 4954 5296
rect 6362 5244 6368 5296
rect 6420 5284 6426 5296
rect 6730 5284 6736 5296
rect 6420 5256 6736 5284
rect 6420 5244 6426 5256
rect 6730 5244 6736 5256
rect 6788 5244 6794 5296
rect 7834 5244 7840 5296
rect 7892 5284 7898 5296
rect 8570 5284 8576 5296
rect 7892 5256 8576 5284
rect 7892 5244 7898 5256
rect 8570 5244 8576 5256
rect 8628 5244 8634 5296
rect 10045 5287 10103 5293
rect 10045 5253 10057 5287
rect 10091 5284 10103 5287
rect 10686 5284 10692 5296
rect 10091 5256 10692 5284
rect 10091 5253 10103 5256
rect 10045 5247 10103 5253
rect 10686 5244 10692 5256
rect 10744 5244 10750 5296
rect 10980 5284 11008 5324
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 12158 5352 12164 5364
rect 12032 5324 12164 5352
rect 12032 5312 12038 5324
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 12894 5352 12900 5364
rect 12483 5324 12900 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 13078 5312 13084 5364
rect 13136 5352 13142 5364
rect 13633 5355 13691 5361
rect 13633 5352 13645 5355
rect 13136 5324 13645 5352
rect 13136 5312 13142 5324
rect 13633 5321 13645 5324
rect 13679 5321 13691 5355
rect 13998 5352 14004 5364
rect 13633 5315 13691 5321
rect 13740 5324 14004 5352
rect 11146 5284 11152 5296
rect 10980 5256 11152 5284
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5185 2559 5219
rect 2501 5179 2559 5185
rect 4071 5188 5028 5216
rect 2225 5151 2283 5157
rect 2225 5117 2237 5151
rect 2271 5117 2283 5151
rect 2225 5111 2283 5117
rect 2406 5108 2412 5160
rect 2464 5148 2470 5160
rect 2516 5148 2544 5179
rect 3053 5151 3111 5157
rect 2464 5120 3004 5148
rect 2464 5108 2470 5120
rect 2976 5080 3004 5120
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 3142 5148 3148 5160
rect 3099 5120 3148 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 3320 5151 3378 5157
rect 3320 5117 3332 5151
rect 3366 5148 3378 5151
rect 3694 5148 3700 5160
rect 3366 5120 3700 5148
rect 3366 5117 3378 5120
rect 3320 5111 3378 5117
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 4071 5080 4099 5188
rect 4890 5148 4896 5160
rect 4851 5120 4896 5148
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 5000 5148 5028 5188
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 11072 5225 11100 5256
rect 11146 5244 11152 5256
rect 11204 5244 11210 5296
rect 13740 5284 13768 5324
rect 13998 5312 14004 5324
rect 14056 5312 14062 5364
rect 14366 5352 14372 5364
rect 14108 5324 14372 5352
rect 14108 5284 14136 5324
rect 14366 5312 14372 5324
rect 14424 5352 14430 5364
rect 14642 5352 14648 5364
rect 14424 5324 14648 5352
rect 14424 5312 14430 5324
rect 14642 5312 14648 5324
rect 14700 5312 14706 5364
rect 15013 5287 15071 5293
rect 15013 5284 15025 5287
rect 11716 5256 13768 5284
rect 14016 5256 14136 5284
rect 14200 5256 15025 5284
rect 11716 5225 11744 5256
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 9732 5188 10977 5216
rect 9732 5176 9738 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 10965 5179 11023 5185
rect 11057 5219 11115 5225
rect 11057 5185 11069 5219
rect 11103 5185 11115 5219
rect 11057 5179 11115 5185
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 12802 5176 12808 5228
rect 12860 5216 12866 5228
rect 12989 5219 13047 5225
rect 12989 5216 13001 5219
rect 12860 5188 13001 5216
rect 12860 5176 12866 5188
rect 12989 5185 13001 5188
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 13078 5176 13084 5228
rect 13136 5216 13142 5228
rect 14016 5216 14044 5256
rect 14200 5216 14228 5256
rect 15013 5253 15025 5256
rect 15059 5253 15071 5287
rect 15013 5247 15071 5253
rect 13136 5188 14044 5216
rect 14108 5188 14228 5216
rect 14277 5219 14335 5225
rect 13136 5176 13142 5188
rect 5160 5151 5218 5157
rect 5160 5148 5172 5151
rect 5000 5120 5172 5148
rect 5160 5117 5172 5120
rect 5206 5148 5218 5151
rect 5442 5148 5448 5160
rect 5206 5120 5448 5148
rect 5206 5117 5218 5120
rect 5160 5111 5218 5117
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 5592 5120 6837 5148
rect 5592 5108 5598 5120
rect 6825 5117 6837 5120
rect 6871 5148 6883 5151
rect 8665 5151 8723 5157
rect 8665 5148 8677 5151
rect 6871 5120 8677 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 8665 5117 8677 5120
rect 8711 5148 8723 5151
rect 9398 5148 9404 5160
rect 8711 5120 9404 5148
rect 8711 5117 8723 5120
rect 8665 5111 8723 5117
rect 9398 5108 9404 5120
rect 9456 5148 9462 5160
rect 9858 5148 9864 5160
rect 9456 5120 9864 5148
rect 9456 5108 9462 5120
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 10410 5108 10416 5160
rect 10468 5148 10474 5160
rect 11790 5148 11796 5160
rect 10468 5120 11796 5148
rect 10468 5108 10474 5120
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 11974 5108 11980 5160
rect 12032 5148 12038 5160
rect 14108 5148 14136 5188
rect 14277 5185 14289 5219
rect 14323 5185 14335 5219
rect 14642 5216 14648 5228
rect 14277 5179 14335 5185
rect 14384 5188 14648 5216
rect 12032 5120 14136 5148
rect 12032 5108 12038 5120
rect 14182 5108 14188 5160
rect 14240 5148 14246 5160
rect 14292 5148 14320 5179
rect 14240 5120 14320 5148
rect 14240 5108 14246 5120
rect 6178 5080 6184 5092
rect 2976 5052 4099 5080
rect 6104 5052 6184 5080
rect 1854 5012 1860 5024
rect 1815 4984 1860 5012
rect 1854 4972 1860 4984
rect 1912 4972 1918 5024
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2372 4984 2417 5012
rect 2372 4972 2378 4984
rect 3326 4972 3332 5024
rect 3384 5012 3390 5024
rect 6104 5012 6132 5052
rect 6178 5040 6184 5052
rect 6236 5040 6242 5092
rect 7098 5089 7104 5092
rect 7092 5080 7104 5089
rect 7011 5052 7104 5080
rect 7092 5043 7104 5052
rect 7156 5080 7162 5092
rect 7834 5080 7840 5092
rect 7156 5052 7840 5080
rect 7098 5040 7104 5043
rect 7156 5040 7162 5052
rect 7834 5040 7840 5052
rect 7892 5040 7898 5092
rect 8570 5040 8576 5092
rect 8628 5080 8634 5092
rect 8754 5080 8760 5092
rect 8628 5052 8760 5080
rect 8628 5040 8634 5052
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 8932 5083 8990 5089
rect 8932 5049 8944 5083
rect 8978 5080 8990 5083
rect 9122 5080 9128 5092
rect 8978 5052 9128 5080
rect 8978 5049 8990 5052
rect 8932 5043 8990 5049
rect 9122 5040 9128 5052
rect 9180 5040 9186 5092
rect 10594 5080 10600 5092
rect 9232 5052 10600 5080
rect 6270 5012 6276 5024
rect 3384 4984 6132 5012
rect 6231 4984 6276 5012
rect 3384 4972 3390 4984
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 9232 5012 9260 5052
rect 10594 5040 10600 5052
rect 10652 5040 10658 5092
rect 10778 5040 10784 5092
rect 10836 5080 10842 5092
rect 11882 5080 11888 5092
rect 10836 5052 11888 5080
rect 10836 5040 10842 5052
rect 11882 5040 11888 5052
rect 11940 5040 11946 5092
rect 12526 5040 12532 5092
rect 12584 5080 12590 5092
rect 13446 5080 13452 5092
rect 12584 5052 13308 5080
rect 13407 5052 13452 5080
rect 12584 5040 12590 5052
rect 6880 4984 9260 5012
rect 6880 4972 6886 4984
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 9950 5012 9956 5024
rect 9732 4984 9956 5012
rect 9732 4972 9738 4984
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 10134 4972 10140 5024
rect 10192 5012 10198 5024
rect 10505 5015 10563 5021
rect 10505 5012 10517 5015
rect 10192 4984 10517 5012
rect 10192 4972 10198 4984
rect 10505 4981 10517 4984
rect 10551 4981 10563 5015
rect 10505 4975 10563 4981
rect 10873 5015 10931 5021
rect 10873 4981 10885 5015
rect 10919 5012 10931 5015
rect 11606 5012 11612 5024
rect 10919 4984 11612 5012
rect 10919 4981 10931 4984
rect 10873 4975 10931 4981
rect 11606 4972 11612 4984
rect 11664 5012 11670 5024
rect 12250 5012 12256 5024
rect 11664 4984 12256 5012
rect 11664 4972 11670 4984
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 12710 4972 12716 5024
rect 12768 5012 12774 5024
rect 12805 5015 12863 5021
rect 12805 5012 12817 5015
rect 12768 4984 12817 5012
rect 12768 4972 12774 4984
rect 12805 4981 12817 4984
rect 12851 4981 12863 5015
rect 12805 4975 12863 4981
rect 12897 5015 12955 5021
rect 12897 4981 12909 5015
rect 12943 5012 12955 5015
rect 13078 5012 13084 5024
rect 12943 4984 13084 5012
rect 12943 4981 12955 4984
rect 12897 4975 12955 4981
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 13280 5012 13308 5052
rect 13446 5040 13452 5052
rect 13504 5080 13510 5092
rect 14001 5083 14059 5089
rect 14001 5080 14013 5083
rect 13504 5052 14013 5080
rect 13504 5040 13510 5052
rect 14001 5049 14013 5052
rect 14047 5049 14059 5083
rect 14001 5043 14059 5049
rect 14093 5083 14151 5089
rect 14093 5049 14105 5083
rect 14139 5080 14151 5083
rect 14384 5080 14412 5188
rect 14642 5176 14648 5188
rect 14700 5216 14706 5228
rect 15286 5216 15292 5228
rect 14700 5188 15292 5216
rect 14700 5176 14706 5188
rect 15286 5176 15292 5188
rect 15344 5176 15350 5228
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5117 14887 5151
rect 14829 5111 14887 5117
rect 14139 5052 14412 5080
rect 14139 5049 14151 5052
rect 14093 5043 14151 5049
rect 14844 5012 14872 5111
rect 13280 4984 14872 5012
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 3326 4808 3332 4820
rect 1412 4780 3332 4808
rect 1412 4681 1440 4780
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 7558 4808 7564 4820
rect 4448 4780 7564 4808
rect 2148 4712 2544 4740
rect 2148 4681 2176 4712
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4641 1455 4675
rect 1397 4635 1455 4641
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4641 2191 4675
rect 2133 4635 2191 4641
rect 2222 4632 2228 4684
rect 2280 4672 2286 4684
rect 2389 4675 2447 4681
rect 2389 4672 2401 4675
rect 2280 4644 2401 4672
rect 2280 4632 2286 4644
rect 2389 4641 2401 4644
rect 2435 4641 2447 4675
rect 2516 4672 2544 4712
rect 2590 4700 2596 4752
rect 2648 4740 2654 4752
rect 4448 4740 4476 4780
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 8941 4811 8999 4817
rect 8941 4777 8953 4811
rect 8987 4808 8999 4811
rect 11241 4811 11299 4817
rect 8987 4780 11100 4808
rect 8987 4777 8999 4780
rect 8941 4771 8999 4777
rect 11072 4752 11100 4780
rect 11241 4777 11253 4811
rect 11287 4808 11299 4811
rect 11790 4808 11796 4820
rect 11287 4780 11796 4808
rect 11287 4777 11299 4780
rect 11241 4771 11299 4777
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 12437 4811 12495 4817
rect 12437 4808 12449 4811
rect 12400 4780 12449 4808
rect 12400 4768 12406 4780
rect 12437 4777 12449 4780
rect 12483 4777 12495 4811
rect 12437 4771 12495 4777
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 12802 4808 12808 4820
rect 12676 4780 12808 4808
rect 12676 4768 12682 4780
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 13170 4768 13176 4820
rect 13228 4808 13234 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 13228 4780 13277 4808
rect 13228 4768 13234 4780
rect 13265 4777 13277 4780
rect 13311 4777 13323 4811
rect 13265 4771 13323 4777
rect 2648 4712 4476 4740
rect 4525 4743 4583 4749
rect 2648 4700 2654 4712
rect 4525 4709 4537 4743
rect 4571 4740 4583 4743
rect 6822 4740 6828 4752
rect 4571 4712 6828 4740
rect 4571 4709 4583 4712
rect 4525 4703 4583 4709
rect 6822 4700 6828 4712
rect 6880 4700 6886 4752
rect 7208 4712 8524 4740
rect 3142 4672 3148 4684
rect 2516 4644 3148 4672
rect 2389 4635 2447 4641
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 5074 4672 5080 4684
rect 4479 4644 5080 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 5074 4632 5080 4644
rect 5132 4632 5138 4684
rect 5534 4681 5540 4684
rect 5528 4672 5540 4681
rect 5495 4644 5540 4672
rect 5528 4635 5540 4644
rect 5534 4632 5540 4635
rect 5592 4632 5598 4684
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 5868 4644 6684 4672
rect 5868 4632 5874 4644
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 3510 4536 3516 4548
rect 3471 4508 3516 4536
rect 3510 4496 3516 4508
rect 3568 4496 3574 4548
rect 3694 4496 3700 4548
rect 3752 4536 3758 4548
rect 4338 4536 4344 4548
rect 3752 4508 4344 4536
rect 3752 4496 3758 4508
rect 4338 4496 4344 4508
rect 4396 4496 4402 4548
rect 4724 4536 4752 4567
rect 4890 4564 4896 4616
rect 4948 4604 4954 4616
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 4948 4576 5273 4604
rect 4948 4564 4954 4576
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 6656 4604 6684 4644
rect 6730 4632 6736 4684
rect 6788 4672 6794 4684
rect 7101 4675 7159 4681
rect 7101 4672 7113 4675
rect 6788 4644 7113 4672
rect 6788 4632 6794 4644
rect 7101 4641 7113 4644
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 7208 4604 7236 4712
rect 7374 4681 7380 4684
rect 7368 4672 7380 4681
rect 7335 4644 7380 4672
rect 7368 4635 7380 4644
rect 7374 4632 7380 4635
rect 7432 4632 7438 4684
rect 6656 4576 7236 4604
rect 5261 4567 5319 4573
rect 8496 4545 8524 4712
rect 8662 4700 8668 4752
rect 8720 4740 8726 4752
rect 8720 4712 9812 4740
rect 8720 4700 8726 4712
rect 8754 4632 8760 4684
rect 8812 4672 8818 4684
rect 9674 4672 9680 4684
rect 8812 4644 9680 4672
rect 8812 4632 8818 4644
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 8938 4564 8944 4616
rect 8996 4604 9002 4616
rect 9582 4604 9588 4616
rect 8996 4576 9588 4604
rect 8996 4564 9002 4576
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 9784 4604 9812 4712
rect 9950 4700 9956 4752
rect 10008 4740 10014 4752
rect 10045 4743 10103 4749
rect 10045 4740 10057 4743
rect 10008 4712 10057 4740
rect 10008 4700 10014 4712
rect 10045 4709 10057 4712
rect 10091 4709 10103 4743
rect 10045 4703 10103 4709
rect 10137 4743 10195 4749
rect 10137 4709 10149 4743
rect 10183 4740 10195 4743
rect 10410 4740 10416 4752
rect 10183 4712 10416 4740
rect 10183 4709 10195 4712
rect 10137 4703 10195 4709
rect 10410 4700 10416 4712
rect 10468 4740 10474 4752
rect 10870 4740 10876 4752
rect 10468 4712 10876 4740
rect 10468 4700 10474 4712
rect 10870 4700 10876 4712
rect 10928 4700 10934 4752
rect 11054 4700 11060 4752
rect 11112 4700 11118 4752
rect 11146 4700 11152 4752
rect 11204 4740 11210 4752
rect 11204 4712 11468 4740
rect 11204 4700 11210 4712
rect 10778 4632 10784 4684
rect 10836 4672 10842 4684
rect 10836 4644 11284 4672
rect 10836 4632 10842 4644
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 9784 4576 10241 4604
rect 10229 4573 10241 4576
rect 10275 4604 10287 4607
rect 10410 4604 10416 4616
rect 10275 4576 10416 4604
rect 10275 4573 10287 4576
rect 10229 4567 10287 4573
rect 10410 4564 10416 4576
rect 10468 4564 10474 4616
rect 11256 4604 11284 4644
rect 11440 4613 11468 4712
rect 11882 4700 11888 4752
rect 11940 4740 11946 4752
rect 12529 4743 12587 4749
rect 12529 4740 12541 4743
rect 11940 4712 12541 4740
rect 11940 4700 11946 4712
rect 12529 4709 12541 4712
rect 12575 4740 12587 4743
rect 12575 4712 14504 4740
rect 12575 4709 12587 4712
rect 12529 4703 12587 4709
rect 13354 4632 13360 4684
rect 13412 4672 13418 4684
rect 14476 4681 14504 4712
rect 13633 4675 13691 4681
rect 13633 4672 13645 4675
rect 13412 4644 13645 4672
rect 13412 4632 13418 4644
rect 13633 4641 13645 4644
rect 13679 4641 13691 4675
rect 13633 4635 13691 4641
rect 14461 4675 14519 4681
rect 14461 4641 14473 4675
rect 14507 4641 14519 4675
rect 14461 4635 14519 4641
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 11256 4576 11345 4604
rect 11333 4573 11345 4576
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4573 11483 4607
rect 11425 4567 11483 4573
rect 11606 4564 11612 4616
rect 11664 4604 11670 4616
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 11664 4576 12633 4604
rect 11664 4564 11670 4576
rect 12621 4573 12633 4576
rect 12667 4573 12679 4607
rect 12621 4567 12679 4573
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 13725 4607 13783 4613
rect 13725 4604 13737 4607
rect 12768 4576 13737 4604
rect 12768 4564 12774 4576
rect 13725 4573 13737 4576
rect 13771 4573 13783 4607
rect 13725 4567 13783 4573
rect 13817 4607 13875 4613
rect 13817 4573 13829 4607
rect 13863 4604 13875 4607
rect 14182 4604 14188 4616
rect 13863 4576 14188 4604
rect 13863 4573 13875 4576
rect 13817 4567 13875 4573
rect 8481 4539 8539 4545
rect 4724 4508 5304 4536
rect 1581 4471 1639 4477
rect 1581 4437 1593 4471
rect 1627 4468 1639 4471
rect 2498 4468 2504 4480
rect 1627 4440 2504 4468
rect 1627 4437 1639 4440
rect 1581 4431 1639 4437
rect 2498 4428 2504 4440
rect 2556 4428 2562 4480
rect 4065 4471 4123 4477
rect 4065 4437 4077 4471
rect 4111 4468 4123 4471
rect 4154 4468 4160 4480
rect 4111 4440 4160 4468
rect 4111 4437 4123 4440
rect 4065 4431 4123 4437
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 5276 4468 5304 4508
rect 8481 4505 8493 4539
rect 8527 4536 8539 4539
rect 8527 4508 8616 4536
rect 8527 4505 8539 4508
rect 8481 4499 8539 4505
rect 6178 4468 6184 4480
rect 5276 4440 6184 4468
rect 6178 4428 6184 4440
rect 6236 4428 6242 4480
rect 6641 4471 6699 4477
rect 6641 4437 6653 4471
rect 6687 4468 6699 4471
rect 7374 4468 7380 4480
rect 6687 4440 7380 4468
rect 6687 4437 6699 4440
rect 6641 4431 6699 4437
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 8588 4468 8616 4508
rect 8662 4496 8668 4548
rect 8720 4536 8726 4548
rect 12069 4539 12127 4545
rect 12069 4536 12081 4539
rect 8720 4508 12081 4536
rect 8720 4496 8726 4508
rect 12069 4505 12081 4508
rect 12115 4505 12127 4539
rect 12069 4499 12127 4505
rect 13078 4496 13084 4548
rect 13136 4536 13142 4548
rect 13832 4536 13860 4567
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14642 4564 14648 4616
rect 14700 4564 14706 4616
rect 14660 4536 14688 4564
rect 13136 4508 13860 4536
rect 13924 4508 14688 4536
rect 13136 4496 13142 4508
rect 9122 4468 9128 4480
rect 8588 4440 9128 4468
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 9677 4471 9735 4477
rect 9677 4437 9689 4471
rect 9723 4468 9735 4471
rect 9858 4468 9864 4480
rect 9723 4440 9864 4468
rect 9723 4437 9735 4440
rect 9677 4431 9735 4437
rect 9858 4428 9864 4440
rect 9916 4428 9922 4480
rect 10226 4428 10232 4480
rect 10284 4468 10290 4480
rect 10873 4471 10931 4477
rect 10873 4468 10885 4471
rect 10284 4440 10885 4468
rect 10284 4428 10290 4440
rect 10873 4437 10885 4440
rect 10919 4437 10931 4471
rect 10873 4431 10931 4437
rect 11146 4428 11152 4480
rect 11204 4468 11210 4480
rect 13924 4468 13952 4508
rect 11204 4440 13952 4468
rect 11204 4428 11210 4440
rect 13998 4428 14004 4480
rect 14056 4468 14062 4480
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 14056 4440 14657 4468
rect 14056 4428 14062 4440
rect 14645 4437 14657 4440
rect 14691 4437 14703 4471
rect 14645 4431 14703 4437
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 5626 4264 5632 4276
rect 3292 4236 5632 4264
rect 3292 4224 3298 4236
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 8110 4224 8116 4276
rect 8168 4264 8174 4276
rect 8938 4264 8944 4276
rect 8168 4236 8944 4264
rect 8168 4224 8174 4236
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 9861 4267 9919 4273
rect 9861 4264 9873 4267
rect 9824 4236 9873 4264
rect 9824 4224 9830 4236
rect 9861 4233 9873 4236
rect 9907 4233 9919 4267
rect 10318 4264 10324 4276
rect 10231 4236 10324 4264
rect 9861 4227 9919 4233
rect 10318 4224 10324 4236
rect 10376 4264 10382 4276
rect 11057 4267 11115 4273
rect 10376 4236 10640 4264
rect 10376 4224 10382 4236
rect 1857 4199 1915 4205
rect 1857 4165 1869 4199
rect 1903 4196 1915 4199
rect 2866 4196 2872 4208
rect 1903 4168 2872 4196
rect 1903 4165 1915 4168
rect 1857 4159 1915 4165
rect 2866 4156 2872 4168
rect 2924 4156 2930 4208
rect 4433 4199 4491 4205
rect 4433 4165 4445 4199
rect 4479 4196 4491 4199
rect 4706 4196 4712 4208
rect 4479 4168 4712 4196
rect 4479 4165 4491 4168
rect 4433 4159 4491 4165
rect 4706 4156 4712 4168
rect 4764 4156 4770 4208
rect 7834 4156 7840 4208
rect 7892 4196 7898 4208
rect 10336 4196 10364 4224
rect 7892 4168 10364 4196
rect 10612 4196 10640 4236
rect 11057 4233 11069 4267
rect 11103 4264 11115 4267
rect 11790 4264 11796 4276
rect 11103 4236 11796 4264
rect 11103 4233 11115 4236
rect 11057 4227 11115 4233
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 12894 4224 12900 4276
rect 12952 4264 12958 4276
rect 13906 4264 13912 4276
rect 12952 4236 13912 4264
rect 12952 4224 12958 4236
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 14182 4224 14188 4276
rect 14240 4264 14246 4276
rect 14366 4264 14372 4276
rect 14240 4236 14372 4264
rect 14240 4224 14246 4236
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 10612 4168 11652 4196
rect 7892 4156 7898 4168
rect 382 4088 388 4140
rect 440 4128 446 4140
rect 1578 4128 1584 4140
rect 440 4100 1584 4128
rect 440 4088 446 4100
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 2406 4128 2412 4140
rect 2367 4100 2412 4128
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 4890 4128 4896 4140
rect 4264 4100 4896 4128
rect 750 4020 756 4072
rect 808 4060 814 4072
rect 1394 4060 1400 4072
rect 808 4032 1400 4060
rect 808 4020 814 4032
rect 1394 4020 1400 4032
rect 1452 4020 1458 4072
rect 3053 4063 3111 4069
rect 3053 4029 3065 4063
rect 3099 4060 3111 4063
rect 3142 4060 3148 4072
rect 3099 4032 3148 4060
rect 3099 4029 3111 4032
rect 3053 4023 3111 4029
rect 3142 4020 3148 4032
rect 3200 4060 3206 4072
rect 4264 4060 4292 4100
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 6003 4100 6960 4128
rect 6003 4060 6031 4100
rect 3200 4032 4292 4060
rect 4347 4032 6031 4060
rect 3200 4020 3206 4032
rect 3320 3995 3378 4001
rect 3320 3961 3332 3995
rect 3366 3992 3378 3995
rect 4246 3992 4252 4004
rect 3366 3964 4252 3992
rect 3366 3961 3378 3964
rect 3320 3955 3378 3961
rect 4246 3952 4252 3964
rect 4304 3952 4310 4004
rect 2222 3924 2228 3936
rect 2183 3896 2228 3924
rect 2222 3884 2228 3896
rect 2280 3884 2286 3936
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 4347 3924 4375 4032
rect 6178 4020 6184 4072
rect 6236 4060 6242 4072
rect 6236 4032 6684 4060
rect 6236 4020 6242 4032
rect 4982 3952 4988 4004
rect 5040 3992 5046 4004
rect 5166 4001 5172 4004
rect 5160 3992 5172 4001
rect 5040 3964 5172 3992
rect 5040 3952 5046 3964
rect 5160 3955 5172 3964
rect 5224 3992 5230 4004
rect 6656 3992 6684 4032
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6788 4032 6837 4060
rect 6788 4020 6794 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6932 4060 6960 4100
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 9324 4137 9352 4168
rect 9309 4131 9367 4137
rect 8168 4100 9168 4128
rect 8168 4088 8174 4100
rect 8662 4060 8668 4072
rect 6932 4032 8668 4060
rect 6825 4023 6883 4029
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 9140 4069 9168 4100
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 10318 4128 10324 4140
rect 9309 4091 9367 4097
rect 9416 4100 10324 4128
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4060 9183 4063
rect 9416 4060 9444 4100
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 10410 4088 10416 4140
rect 10468 4128 10474 4140
rect 10468 4100 10513 4128
rect 10468 4088 10474 4100
rect 10870 4088 10876 4140
rect 10928 4128 10934 4140
rect 11624 4137 11652 4168
rect 12434 4156 12440 4208
rect 12492 4196 12498 4208
rect 13170 4196 13176 4208
rect 12492 4168 13176 4196
rect 12492 4156 12498 4168
rect 13170 4156 13176 4168
rect 13228 4156 13234 4208
rect 13446 4156 13452 4208
rect 13504 4196 13510 4208
rect 13633 4199 13691 4205
rect 13633 4196 13645 4199
rect 13504 4168 13645 4196
rect 13504 4156 13510 4168
rect 13633 4165 13645 4168
rect 13679 4165 13691 4199
rect 14458 4196 14464 4208
rect 13633 4159 13691 4165
rect 14292 4168 14464 4196
rect 11609 4131 11667 4137
rect 10928 4100 11468 4128
rect 10928 4088 10934 4100
rect 11440 4069 11468 4100
rect 11609 4097 11621 4131
rect 11655 4097 11667 4131
rect 11609 4091 11667 4097
rect 12342 4088 12348 4140
rect 12400 4088 12406 4140
rect 12526 4088 12532 4140
rect 12584 4128 12590 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12584 4100 12909 4128
rect 12584 4088 12590 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 13078 4128 13084 4140
rect 13039 4100 13084 4128
rect 12897 4091 12955 4097
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 13998 4088 14004 4140
rect 14056 4128 14062 4140
rect 14292 4137 14320 4168
rect 14458 4156 14464 4168
rect 14516 4156 14522 4208
rect 15010 4196 15016 4208
rect 14971 4168 15016 4196
rect 15010 4156 15016 4168
rect 15068 4156 15074 4208
rect 14093 4131 14151 4137
rect 14093 4128 14105 4131
rect 14056 4100 14105 4128
rect 14056 4088 14062 4100
rect 14093 4097 14105 4100
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4097 14335 4131
rect 14277 4091 14335 4097
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 15470 4128 15476 4140
rect 14424 4100 15476 4128
rect 14424 4088 14430 4100
rect 15470 4088 15476 4100
rect 15528 4088 15534 4140
rect 9171 4032 9444 4060
rect 10229 4063 10287 4069
rect 9171 4029 9183 4032
rect 9125 4023 9183 4029
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 11425 4063 11483 4069
rect 10275 4032 11008 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 7070 3995 7128 4001
rect 7070 3992 7082 3995
rect 5224 3964 6408 3992
rect 6656 3964 7082 3992
rect 5166 3952 5172 3955
rect 5224 3952 5230 3964
rect 2363 3896 4375 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 5534 3884 5540 3936
rect 5592 3924 5598 3936
rect 6273 3927 6331 3933
rect 6273 3924 6285 3927
rect 5592 3896 6285 3924
rect 5592 3884 5598 3896
rect 6273 3893 6285 3896
rect 6319 3893 6331 3927
rect 6380 3924 6408 3964
rect 7070 3961 7082 3964
rect 7116 3992 7128 3995
rect 7466 3992 7472 4004
rect 7116 3964 7472 3992
rect 7116 3961 7128 3964
rect 7070 3955 7128 3961
rect 7466 3952 7472 3964
rect 7524 3952 7530 4004
rect 7742 3952 7748 4004
rect 7800 3992 7806 4004
rect 8110 3992 8116 4004
rect 7800 3964 8116 3992
rect 7800 3952 7806 3964
rect 8110 3952 8116 3964
rect 8168 3952 8174 4004
rect 10778 3992 10784 4004
rect 8680 3964 10784 3992
rect 8680 3933 8708 3964
rect 10778 3952 10784 3964
rect 10836 3952 10842 4004
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 6380 3896 8217 3924
rect 6273 3887 6331 3893
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 8205 3887 8263 3893
rect 8665 3927 8723 3933
rect 8665 3893 8677 3927
rect 8711 3893 8723 3927
rect 8665 3887 8723 3893
rect 9033 3927 9091 3933
rect 9033 3893 9045 3927
rect 9079 3924 9091 3927
rect 9306 3924 9312 3936
rect 9079 3896 9312 3924
rect 9079 3893 9091 3896
rect 9033 3887 9091 3893
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 10100 3896 10333 3924
rect 10100 3884 10106 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 10321 3887 10379 3893
rect 10410 3884 10416 3936
rect 10468 3924 10474 3936
rect 10686 3924 10692 3936
rect 10468 3896 10692 3924
rect 10468 3884 10474 3896
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 10980 3924 11008 4032
rect 11425 4029 11437 4063
rect 11471 4060 11483 4063
rect 11790 4060 11796 4072
rect 11471 4032 11796 4060
rect 11471 4029 11483 4032
rect 11425 4023 11483 4029
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 11974 4020 11980 4072
rect 12032 4060 12038 4072
rect 12360 4060 12388 4088
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12032 4032 12817 4060
rect 12032 4020 12038 4032
rect 12805 4029 12817 4032
rect 12851 4029 12863 4063
rect 12805 4023 12863 4029
rect 14642 4020 14648 4072
rect 14700 4060 14706 4072
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 14700 4032 14841 4060
rect 14700 4020 14706 4032
rect 14829 4029 14841 4032
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 11330 3952 11336 4004
rect 11388 3992 11394 4004
rect 11517 3995 11575 4001
rect 11517 3992 11529 3995
rect 11388 3964 11529 3992
rect 11388 3952 11394 3964
rect 11517 3961 11529 3964
rect 11563 3961 11575 3995
rect 11517 3955 11575 3961
rect 13262 3952 13268 4004
rect 13320 3992 13326 4004
rect 14001 3995 14059 4001
rect 14001 3992 14013 3995
rect 13320 3964 14013 3992
rect 13320 3952 13326 3964
rect 14001 3961 14013 3964
rect 14047 3961 14059 3995
rect 14001 3955 14059 3961
rect 11698 3924 11704 3936
rect 10980 3896 11704 3924
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 13814 3924 13820 3936
rect 12483 3896 13820 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 1670 3720 1676 3732
rect 1627 3692 1676 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 1670 3680 1676 3692
rect 1728 3680 1734 3732
rect 1946 3720 1952 3732
rect 1907 3692 1952 3720
rect 1946 3680 1952 3692
rect 2004 3680 2010 3732
rect 2041 3723 2099 3729
rect 2041 3689 2053 3723
rect 2087 3720 2099 3723
rect 2590 3720 2596 3732
rect 2087 3692 2596 3720
rect 2087 3689 2099 3692
rect 2041 3683 2099 3689
rect 2590 3680 2596 3692
rect 2648 3680 2654 3732
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 3878 3720 3884 3732
rect 2823 3692 3884 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 5718 3720 5724 3732
rect 4816 3692 5724 3720
rect 2866 3612 2872 3664
rect 2924 3652 2930 3664
rect 3145 3655 3203 3661
rect 3145 3652 3157 3655
rect 2924 3624 3157 3652
rect 2924 3612 2930 3624
rect 3145 3621 3157 3624
rect 3191 3621 3203 3655
rect 3145 3615 3203 3621
rect 3326 3612 3332 3664
rect 3384 3652 3390 3664
rect 4816 3652 4844 3692
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 5920 3692 6776 3720
rect 3384 3624 4844 3652
rect 4893 3655 4951 3661
rect 3384 3612 3390 3624
rect 4893 3621 4905 3655
rect 4939 3652 4951 3655
rect 5920 3652 5948 3692
rect 4939 3624 5948 3652
rect 5988 3655 6046 3661
rect 4939 3621 4951 3624
rect 4893 3615 4951 3621
rect 5988 3621 6000 3655
rect 6034 3652 6046 3655
rect 6270 3652 6276 3664
rect 6034 3624 6276 3652
rect 6034 3621 6046 3624
rect 5988 3615 6046 3621
rect 1854 3544 1860 3596
rect 1912 3584 1918 3596
rect 3237 3587 3295 3593
rect 3237 3584 3249 3587
rect 1912 3556 3249 3584
rect 1912 3544 1918 3556
rect 3237 3553 3249 3556
rect 3283 3553 3295 3587
rect 3237 3547 3295 3553
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 4212 3556 4997 3584
rect 4212 3544 4218 3556
rect 4985 3553 4997 3556
rect 5031 3553 5043 3587
rect 6003 3584 6031 3615
rect 6270 3612 6276 3624
rect 6328 3612 6334 3664
rect 6748 3652 6776 3692
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 8570 3720 8576 3732
rect 6880 3692 8576 3720
rect 6880 3680 6886 3692
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 8938 3720 8944 3732
rect 8899 3692 8944 3720
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 9306 3680 9312 3732
rect 9364 3720 9370 3732
rect 9364 3692 9904 3720
rect 9364 3680 9370 3692
rect 9674 3652 9680 3664
rect 6748 3624 9680 3652
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 4985 3547 5043 3553
rect 5245 3556 6031 3584
rect 1946 3476 1952 3528
rect 2004 3516 2010 3528
rect 2133 3519 2191 3525
rect 2133 3516 2145 3519
rect 2004 3488 2145 3516
rect 2004 3476 2010 3488
rect 2133 3485 2145 3488
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 5123 3519 5181 3525
rect 3467 3488 4936 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 4525 3383 4583 3389
rect 4525 3380 4537 3383
rect 4212 3352 4537 3380
rect 4212 3340 4218 3352
rect 4525 3349 4537 3352
rect 4571 3349 4583 3383
rect 4908 3380 4936 3488
rect 5123 3485 5135 3519
rect 5169 3516 5181 3519
rect 5169 3485 5192 3516
rect 5123 3479 5192 3485
rect 4982 3408 4988 3460
rect 5040 3448 5046 3460
rect 5164 3448 5192 3479
rect 5040 3420 5192 3448
rect 5040 3408 5046 3420
rect 5245 3380 5273 3556
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 7558 3584 7564 3596
rect 6788 3556 7564 3584
rect 6788 3544 6794 3556
rect 7558 3544 7564 3556
rect 7616 3544 7622 3596
rect 7828 3587 7886 3593
rect 7828 3553 7840 3587
rect 7874 3584 7886 3587
rect 9766 3584 9772 3596
rect 7874 3556 9772 3584
rect 7874 3553 7886 3556
rect 7828 3547 7886 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 9876 3584 9904 3692
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 12342 3720 12348 3732
rect 10100 3692 12348 3720
rect 10100 3680 10106 3692
rect 12342 3680 12348 3692
rect 12400 3680 12406 3732
rect 12437 3723 12495 3729
rect 12437 3689 12449 3723
rect 12483 3720 12495 3723
rect 13446 3720 13452 3732
rect 12483 3692 13452 3720
rect 12483 3689 12495 3692
rect 12437 3683 12495 3689
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 10008 3624 11560 3652
rect 10008 3612 10014 3624
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 9876 3556 10057 3584
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3584 10195 3587
rect 10318 3584 10324 3596
rect 10183 3556 10324 3584
rect 10183 3553 10195 3556
rect 10137 3547 10195 3553
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 11241 3587 11299 3593
rect 11241 3553 11253 3587
rect 11287 3584 11299 3587
rect 11422 3584 11428 3596
rect 11287 3556 11428 3584
rect 11287 3553 11299 3556
rect 11241 3547 11299 3553
rect 11422 3544 11428 3556
rect 11480 3544 11486 3596
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5500 3488 5733 3516
rect 5500 3476 5506 3488
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 8570 3476 8576 3528
rect 8628 3516 8634 3528
rect 10229 3519 10287 3525
rect 8628 3488 9352 3516
rect 8628 3476 8634 3488
rect 9324 3448 9352 3488
rect 10229 3485 10241 3519
rect 10275 3485 10287 3519
rect 11330 3516 11336 3528
rect 11291 3488 11336 3516
rect 10229 3479 10287 3485
rect 9677 3451 9735 3457
rect 9677 3448 9689 3451
rect 8680 3420 9260 3448
rect 9324 3420 9689 3448
rect 7098 3380 7104 3392
rect 4908 3352 5273 3380
rect 7059 3352 7104 3380
rect 4525 3343 4583 3349
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 8202 3340 8208 3392
rect 8260 3380 8266 3392
rect 8680 3380 8708 3420
rect 8260 3352 8708 3380
rect 9232 3380 9260 3420
rect 9677 3417 9689 3420
rect 9723 3417 9735 3451
rect 9677 3411 9735 3417
rect 10244 3380 10272 3479
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 11532 3525 11560 3624
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 11974 3652 11980 3664
rect 11756 3624 11980 3652
rect 11756 3612 11762 3624
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 12529 3655 12587 3661
rect 12529 3621 12541 3655
rect 12575 3652 12587 3655
rect 12894 3652 12900 3664
rect 12575 3624 12900 3652
rect 12575 3621 12587 3624
rect 12529 3615 12587 3621
rect 12894 3612 12900 3624
rect 12952 3612 12958 3664
rect 13170 3612 13176 3664
rect 13228 3652 13234 3664
rect 13633 3655 13691 3661
rect 13633 3652 13645 3655
rect 13228 3624 13645 3652
rect 13228 3612 13234 3624
rect 13633 3621 13645 3624
rect 13679 3652 13691 3655
rect 13679 3624 14504 3652
rect 13679 3621 13691 3624
rect 13633 3615 13691 3621
rect 11882 3544 11888 3596
rect 11940 3584 11946 3596
rect 14476 3593 14504 3624
rect 13725 3587 13783 3593
rect 13725 3584 13737 3587
rect 11940 3556 13737 3584
rect 11940 3544 11946 3556
rect 13725 3553 13737 3556
rect 13771 3553 13783 3587
rect 13725 3547 13783 3553
rect 14461 3587 14519 3593
rect 14461 3553 14473 3587
rect 14507 3553 14519 3587
rect 14461 3547 14519 3553
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3516 11575 3519
rect 11606 3516 11612 3528
rect 11563 3488 11612 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 12621 3519 12679 3525
rect 12621 3516 12633 3519
rect 12492 3488 12633 3516
rect 12492 3476 12498 3488
rect 12621 3485 12633 3488
rect 12667 3516 12679 3519
rect 13078 3516 13084 3528
rect 12667 3488 13084 3516
rect 12667 3485 12679 3488
rect 12621 3479 12679 3485
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3485 13967 3519
rect 13909 3479 13967 3485
rect 10410 3408 10416 3460
rect 10468 3448 10474 3460
rect 13354 3448 13360 3460
rect 10468 3420 13360 3448
rect 10468 3408 10474 3420
rect 13354 3408 13360 3420
rect 13412 3408 13418 3460
rect 13814 3408 13820 3460
rect 13872 3448 13878 3460
rect 13924 3448 13952 3479
rect 14642 3448 14648 3460
rect 13872 3420 13952 3448
rect 14603 3420 14648 3448
rect 13872 3408 13878 3420
rect 14642 3408 14648 3420
rect 14700 3408 14706 3460
rect 9232 3352 10272 3380
rect 8260 3340 8266 3352
rect 10594 3340 10600 3392
rect 10652 3380 10658 3392
rect 10873 3383 10931 3389
rect 10873 3380 10885 3383
rect 10652 3352 10885 3380
rect 10652 3340 10658 3352
rect 10873 3349 10885 3352
rect 10919 3349 10931 3383
rect 12066 3380 12072 3392
rect 12027 3352 12072 3380
rect 10873 3343 10931 3349
rect 12066 3340 12072 3352
rect 12124 3340 12130 3392
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 12894 3380 12900 3392
rect 12676 3352 12900 3380
rect 12676 3340 12682 3352
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13265 3383 13323 3389
rect 13265 3349 13277 3383
rect 13311 3380 13323 3383
rect 14090 3380 14096 3392
rect 13311 3352 14096 3380
rect 13311 3349 13323 3352
rect 13265 3343 13323 3349
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 2314 3136 2320 3188
rect 2372 3176 2378 3188
rect 2501 3179 2559 3185
rect 2501 3176 2513 3179
rect 2372 3148 2513 3176
rect 2372 3136 2378 3148
rect 2501 3145 2513 3148
rect 2547 3145 2559 3179
rect 2501 3139 2559 3145
rect 3697 3179 3755 3185
rect 3697 3145 3709 3179
rect 3743 3176 3755 3179
rect 4246 3176 4252 3188
rect 3743 3148 4252 3176
rect 3743 3145 3755 3148
rect 3697 3139 3755 3145
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 5534 3176 5540 3188
rect 4356 3148 5540 3176
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 2004 3080 4292 3108
rect 2004 3068 2010 3080
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3040 3203 3043
rect 3326 3040 3332 3052
rect 3191 3012 3332 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 4154 3040 4160 3052
rect 4115 3012 4160 3040
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2972 1639 2975
rect 1670 2972 1676 2984
rect 1627 2944 1676 2972
rect 1627 2941 1639 2944
rect 1581 2935 1639 2941
rect 1670 2932 1676 2944
rect 1728 2932 1734 2984
rect 4062 2972 4068 2984
rect 4023 2944 4068 2972
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 4264 2972 4292 3080
rect 4356 3049 4384 3148
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 5626 3136 5632 3188
rect 5684 3176 5690 3188
rect 9861 3179 9919 3185
rect 9861 3176 9873 3179
rect 5684 3148 9873 3176
rect 5684 3136 5690 3148
rect 9861 3145 9873 3148
rect 9907 3145 9919 3179
rect 11514 3176 11520 3188
rect 9861 3139 9919 3145
rect 9968 3148 11520 3176
rect 5902 3068 5908 3120
rect 5960 3108 5966 3120
rect 6546 3108 6552 3120
rect 5960 3080 6552 3108
rect 5960 3068 5966 3080
rect 6546 3068 6552 3080
rect 6604 3068 6610 3120
rect 7834 3068 7840 3120
rect 7892 3108 7898 3120
rect 8205 3111 8263 3117
rect 8205 3108 8217 3111
rect 7892 3080 8217 3108
rect 7892 3068 7898 3080
rect 8205 3077 8217 3080
rect 8251 3077 8263 3111
rect 9968 3108 9996 3148
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 11606 3136 11612 3188
rect 11664 3176 11670 3188
rect 13170 3176 13176 3188
rect 11664 3148 13176 3176
rect 11664 3136 11670 3148
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 13633 3179 13691 3185
rect 13633 3145 13645 3179
rect 13679 3176 13691 3179
rect 13722 3176 13728 3188
rect 13679 3148 13728 3176
rect 13679 3145 13691 3148
rect 13633 3139 13691 3145
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 8205 3071 8263 3077
rect 9140 3080 9996 3108
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 4724 3012 5028 3040
rect 4724 2972 4752 3012
rect 4890 2972 4896 2984
rect 4264 2944 4752 2972
rect 4851 2944 4896 2972
rect 4890 2932 4896 2944
rect 4948 2932 4954 2984
rect 5000 2972 5028 3012
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 9140 3049 9168 3080
rect 10318 3068 10324 3120
rect 10376 3108 10382 3120
rect 14458 3108 14464 3120
rect 10376 3080 14464 3108
rect 10376 3068 10382 3080
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 15010 3108 15016 3120
rect 14971 3080 15016 3108
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6788 3012 6837 3040
rect 6788 3000 6794 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3009 9183 3043
rect 9306 3040 9312 3052
rect 9267 3012 9312 3040
rect 9125 3003 9183 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 9950 3000 9956 3052
rect 10008 3040 10014 3052
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 10008 3012 10425 3040
rect 10008 3000 10014 3012
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 11609 3043 11667 3049
rect 11609 3040 11621 3043
rect 10413 3003 10471 3009
rect 10520 3012 11621 3040
rect 5149 2975 5207 2981
rect 5149 2972 5161 2975
rect 5000 2944 5161 2972
rect 5149 2941 5161 2944
rect 5195 2972 5207 2975
rect 6362 2972 6368 2984
rect 5195 2944 6368 2972
rect 5195 2941 5207 2944
rect 5149 2935 5207 2941
rect 6362 2932 6368 2944
rect 6420 2932 6426 2984
rect 10520 2972 10548 3012
rect 11609 3009 11621 3012
rect 11655 3040 11667 3043
rect 13081 3043 13139 3049
rect 13081 3040 13093 3043
rect 11655 3012 13093 3040
rect 11655 3009 11667 3012
rect 11609 3003 11667 3009
rect 13081 3009 13093 3012
rect 13127 3040 13139 3043
rect 13722 3040 13728 3052
rect 13127 3012 13728 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 14090 3040 14096 3052
rect 14051 3012 14096 3040
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14274 3040 14280 3052
rect 14187 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3040 14338 3052
rect 14550 3040 14556 3052
rect 14332 3012 14556 3040
rect 14332 3000 14338 3012
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 11146 2972 11152 2984
rect 7085 2944 10548 2972
rect 10980 2944 11152 2972
rect 1854 2904 1860 2916
rect 1815 2876 1860 2904
rect 1854 2864 1860 2876
rect 1912 2864 1918 2916
rect 2961 2907 3019 2913
rect 2961 2873 2973 2907
rect 3007 2904 3019 2907
rect 3007 2876 5273 2904
rect 3007 2873 3019 2876
rect 2961 2867 3019 2873
rect 2869 2839 2927 2845
rect 2869 2805 2881 2839
rect 2915 2836 2927 2839
rect 5074 2836 5080 2848
rect 2915 2808 5080 2836
rect 2915 2805 2927 2808
rect 2869 2799 2927 2805
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 5245 2836 5273 2876
rect 5810 2864 5816 2916
rect 5868 2904 5874 2916
rect 6454 2904 6460 2916
rect 5868 2876 6460 2904
rect 5868 2864 5874 2876
rect 6454 2864 6460 2876
rect 6512 2864 6518 2916
rect 6730 2864 6736 2916
rect 6788 2904 6794 2916
rect 7085 2913 7113 2944
rect 7070 2907 7128 2913
rect 7070 2904 7082 2907
rect 6788 2876 7082 2904
rect 6788 2864 6794 2876
rect 7070 2873 7082 2876
rect 7116 2873 7128 2907
rect 7070 2867 7128 2873
rect 7190 2864 7196 2916
rect 7248 2904 7254 2916
rect 7742 2904 7748 2916
rect 7248 2876 7748 2904
rect 7248 2864 7254 2876
rect 7742 2864 7748 2876
rect 7800 2864 7806 2916
rect 10042 2904 10048 2916
rect 8680 2876 10048 2904
rect 5534 2836 5540 2848
rect 5245 2808 5540 2836
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 6273 2839 6331 2845
rect 6273 2805 6285 2839
rect 6319 2836 6331 2839
rect 8202 2836 8208 2848
rect 6319 2808 8208 2836
rect 6319 2805 6331 2808
rect 6273 2799 6331 2805
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 8680 2845 8708 2876
rect 10042 2864 10048 2876
rect 10100 2864 10106 2916
rect 10321 2907 10379 2913
rect 10321 2873 10333 2907
rect 10367 2904 10379 2907
rect 10980 2904 11008 2944
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 11514 2972 11520 2984
rect 11475 2944 11520 2972
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 11790 2932 11796 2984
rect 11848 2972 11854 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 11848 2944 14841 2972
rect 11848 2932 11854 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 12526 2904 12532 2916
rect 10367 2876 11008 2904
rect 11072 2876 12532 2904
rect 10367 2873 10379 2876
rect 10321 2867 10379 2873
rect 8665 2839 8723 2845
rect 8665 2805 8677 2839
rect 8711 2805 8723 2839
rect 9030 2836 9036 2848
rect 8991 2808 9036 2836
rect 8665 2799 8723 2805
rect 9030 2796 9036 2808
rect 9088 2796 9094 2848
rect 9769 2839 9827 2845
rect 9769 2805 9781 2839
rect 9815 2836 9827 2839
rect 10229 2839 10287 2845
rect 10229 2836 10241 2839
rect 9815 2808 10241 2836
rect 9815 2805 9827 2808
rect 9769 2799 9827 2805
rect 10229 2805 10241 2808
rect 10275 2836 10287 2839
rect 10410 2836 10416 2848
rect 10275 2808 10416 2836
rect 10275 2805 10287 2808
rect 10229 2799 10287 2805
rect 10410 2796 10416 2808
rect 10468 2796 10474 2848
rect 11072 2845 11100 2876
rect 12526 2864 12532 2876
rect 12584 2864 12590 2916
rect 12805 2907 12863 2913
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 13262 2904 13268 2916
rect 12851 2876 13268 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 13262 2864 13268 2876
rect 13320 2864 13326 2916
rect 13446 2864 13452 2916
rect 13504 2904 13510 2916
rect 13504 2876 14872 2904
rect 13504 2864 13510 2876
rect 14844 2848 14872 2876
rect 11057 2839 11115 2845
rect 11057 2805 11069 2839
rect 11103 2805 11115 2839
rect 11057 2799 11115 2805
rect 11238 2796 11244 2848
rect 11296 2836 11302 2848
rect 11425 2839 11483 2845
rect 11425 2836 11437 2839
rect 11296 2808 11437 2836
rect 11296 2796 11302 2808
rect 11425 2805 11437 2808
rect 11471 2805 11483 2839
rect 11425 2799 11483 2805
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12897 2839 12955 2845
rect 12492 2808 12537 2836
rect 12492 2796 12498 2808
rect 12897 2805 12909 2839
rect 12943 2836 12955 2839
rect 12986 2836 12992 2848
rect 12943 2808 12992 2836
rect 12943 2805 12955 2808
rect 12897 2799 12955 2805
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 13170 2796 13176 2848
rect 13228 2836 13234 2848
rect 13630 2836 13636 2848
rect 13228 2808 13636 2836
rect 13228 2796 13234 2808
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 14001 2839 14059 2845
rect 14001 2805 14013 2839
rect 14047 2836 14059 2839
rect 14458 2836 14464 2848
rect 14047 2808 14464 2836
rect 14047 2805 14059 2808
rect 14001 2799 14059 2805
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 14826 2796 14832 2848
rect 14884 2796 14890 2848
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 4982 2632 4988 2644
rect 2148 2604 4988 2632
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 2038 2496 2044 2508
rect 1443 2468 2044 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 2038 2456 2044 2468
rect 2096 2456 2102 2508
rect 2148 2505 2176 2604
rect 4982 2592 4988 2604
rect 5040 2632 5046 2644
rect 5442 2632 5448 2644
rect 5040 2604 5448 2632
rect 5040 2592 5046 2604
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 6362 2632 6368 2644
rect 6323 2604 6368 2632
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2632 6975 2635
rect 7006 2632 7012 2644
rect 6963 2604 7012 2632
rect 6963 2601 6975 2604
rect 6917 2595 6975 2601
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 7377 2635 7435 2641
rect 7377 2601 7389 2635
rect 7423 2632 7435 2635
rect 7558 2632 7564 2644
rect 7423 2604 7564 2632
rect 7423 2601 7435 2604
rect 7377 2595 7435 2601
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 8113 2635 8171 2641
rect 8113 2601 8125 2635
rect 8159 2601 8171 2635
rect 10042 2632 10048 2644
rect 8113 2595 8171 2601
rect 8404 2604 10048 2632
rect 4706 2524 4712 2576
rect 4764 2564 4770 2576
rect 5230 2567 5288 2573
rect 5230 2564 5242 2567
rect 4764 2536 5242 2564
rect 4764 2524 4770 2536
rect 5230 2533 5242 2536
rect 5276 2533 5288 2567
rect 5230 2527 5288 2533
rect 5534 2524 5540 2576
rect 5592 2564 5598 2576
rect 8128 2564 8156 2595
rect 5592 2536 8156 2564
rect 5592 2524 5598 2536
rect 2133 2499 2191 2505
rect 2133 2465 2145 2499
rect 2179 2465 2191 2499
rect 2133 2459 2191 2465
rect 2400 2499 2458 2505
rect 2400 2465 2412 2499
rect 2446 2496 2458 2499
rect 2866 2496 2872 2508
rect 2446 2468 2872 2496
rect 2446 2465 2458 2468
rect 2400 2459 2458 2465
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 3970 2456 3976 2508
rect 4028 2496 4034 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 4028 2468 4077 2496
rect 4028 2456 4034 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 8404 2496 8432 2604
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 10226 2632 10232 2644
rect 10187 2604 10232 2632
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 10965 2635 11023 2641
rect 10965 2601 10977 2635
rect 11011 2601 11023 2635
rect 11330 2632 11336 2644
rect 11291 2604 11336 2632
rect 10965 2595 11023 2601
rect 9582 2564 9588 2576
rect 8772 2536 9588 2564
rect 8772 2508 8800 2536
rect 9582 2524 9588 2536
rect 9640 2524 9646 2576
rect 10134 2564 10140 2576
rect 10095 2536 10140 2564
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 10980 2564 11008 2595
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 11422 2592 11428 2644
rect 11480 2632 11486 2644
rect 12161 2635 12219 2641
rect 12161 2632 12173 2635
rect 11480 2604 12173 2632
rect 11480 2592 11486 2604
rect 12161 2601 12173 2604
rect 12207 2601 12219 2635
rect 12161 2595 12219 2601
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 13081 2635 13139 2641
rect 13081 2632 13093 2635
rect 12492 2604 13093 2632
rect 12492 2592 12498 2604
rect 13081 2601 13093 2604
rect 13127 2601 13139 2635
rect 13081 2595 13139 2601
rect 14182 2592 14188 2644
rect 14240 2632 14246 2644
rect 14277 2635 14335 2641
rect 14277 2632 14289 2635
rect 14240 2604 14289 2632
rect 14240 2592 14246 2604
rect 14277 2601 14289 2604
rect 14323 2601 14335 2635
rect 14277 2595 14335 2601
rect 12710 2564 12716 2576
rect 10980 2536 12716 2564
rect 12710 2524 12716 2536
rect 12768 2524 12774 2576
rect 12986 2564 12992 2576
rect 12947 2536 12992 2564
rect 12986 2524 12992 2536
rect 13044 2524 13050 2576
rect 7331 2468 8432 2496
rect 8481 2499 8539 2505
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 8481 2465 8493 2499
rect 8527 2496 8539 2499
rect 8754 2496 8760 2508
rect 8527 2468 8760 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 8754 2456 8760 2468
rect 8812 2456 8818 2508
rect 9490 2496 9496 2508
rect 9451 2468 9496 2496
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 10686 2456 10692 2508
rect 10744 2496 10750 2508
rect 10744 2468 11560 2496
rect 10744 2456 10750 2468
rect 4338 2428 4344 2440
rect 4299 2400 4344 2428
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 4982 2428 4988 2440
rect 4943 2400 4988 2428
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 7466 2428 7472 2440
rect 7427 2400 7472 2428
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 8570 2428 8576 2440
rect 8168 2400 8576 2428
rect 8168 2388 8174 2400
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 7374 2320 7380 2372
rect 7432 2360 7438 2372
rect 8680 2360 8708 2391
rect 9306 2388 9312 2440
rect 9364 2428 9370 2440
rect 11532 2437 11560 2468
rect 11790 2456 11796 2508
rect 11848 2496 11854 2508
rect 12345 2499 12403 2505
rect 12345 2496 12357 2499
rect 11848 2468 12357 2496
rect 11848 2456 11854 2468
rect 12345 2465 12357 2468
rect 12391 2465 12403 2499
rect 12345 2459 12403 2465
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 12492 2468 14197 2496
rect 12492 2456 12498 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 15194 2496 15200 2508
rect 15155 2468 15200 2496
rect 14185 2459 14243 2465
rect 15194 2456 15200 2468
rect 15252 2456 15258 2508
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 9364 2400 10333 2428
rect 9364 2388 9370 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 11425 2431 11483 2437
rect 11425 2397 11437 2431
rect 11471 2397 11483 2431
rect 11425 2391 11483 2397
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 9858 2360 9864 2372
rect 7432 2332 8708 2360
rect 9140 2332 9864 2360
rect 7432 2320 7438 2332
rect 106 2252 112 2304
rect 164 2292 170 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 164 2264 1593 2292
rect 164 2252 170 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 6730 2292 6736 2304
rect 3559 2264 6736 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 6730 2252 6736 2264
rect 6788 2252 6794 2304
rect 8202 2252 8208 2304
rect 8260 2292 8266 2304
rect 9140 2292 9168 2332
rect 9858 2320 9864 2332
rect 9916 2360 9922 2372
rect 11440 2360 11468 2391
rect 12526 2388 12532 2440
rect 12584 2428 12590 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 12584 2400 13185 2428
rect 12584 2388 12590 2400
rect 13173 2397 13185 2400
rect 13219 2428 13231 2431
rect 14369 2431 14427 2437
rect 14369 2428 14381 2431
rect 13219 2400 14381 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 14369 2397 14381 2400
rect 14415 2428 14427 2431
rect 14550 2428 14556 2440
rect 14415 2400 14556 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 11882 2360 11888 2372
rect 9916 2332 11888 2360
rect 9916 2320 9922 2332
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 12621 2363 12679 2369
rect 12621 2329 12633 2363
rect 12667 2360 12679 2363
rect 12802 2360 12808 2372
rect 12667 2332 12808 2360
rect 12667 2329 12679 2332
rect 12621 2323 12679 2329
rect 12802 2320 12808 2332
rect 12860 2320 12866 2372
rect 9306 2292 9312 2304
rect 8260 2264 9168 2292
rect 9267 2264 9312 2292
rect 8260 2252 8266 2264
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 9766 2292 9772 2304
rect 9727 2264 9772 2292
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 10042 2252 10048 2304
rect 10100 2292 10106 2304
rect 11330 2292 11336 2304
rect 10100 2264 11336 2292
rect 10100 2252 10106 2264
rect 11330 2252 11336 2264
rect 11388 2292 11394 2304
rect 12250 2292 12256 2304
rect 11388 2264 12256 2292
rect 11388 2252 11394 2264
rect 12250 2252 12256 2264
rect 12308 2252 12314 2304
rect 13814 2292 13820 2304
rect 13775 2264 13820 2292
rect 13814 2252 13820 2264
rect 13872 2252 13878 2304
rect 13906 2252 13912 2304
rect 13964 2292 13970 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 13964 2264 15025 2292
rect 13964 2252 13970 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 4062 2048 4068 2100
rect 4120 2088 4126 2100
rect 8846 2088 8852 2100
rect 4120 2060 8852 2088
rect 4120 2048 4126 2060
rect 8846 2048 8852 2060
rect 8904 2048 8910 2100
rect 9306 2048 9312 2100
rect 9364 2088 9370 2100
rect 11790 2088 11796 2100
rect 9364 2060 11796 2088
rect 9364 2048 9370 2060
rect 11790 2048 11796 2060
rect 11848 2048 11854 2100
rect 937 2023 995 2029
rect 937 1989 949 2023
rect 983 2020 995 2023
rect 13814 2020 13820 2032
rect 983 1992 13820 2020
rect 983 1989 995 1992
rect 937 1983 995 1989
rect 13814 1980 13820 1992
rect 13872 1980 13878 2032
rect 4338 1912 4344 1964
rect 4396 1952 4402 1964
rect 16022 1952 16028 1964
rect 4396 1924 16028 1952
rect 4396 1912 4402 1924
rect 16022 1912 16028 1924
rect 16080 1912 16086 1964
rect 2038 1844 2044 1896
rect 2096 1884 2102 1896
rect 8754 1884 8760 1896
rect 2096 1856 8760 1884
rect 2096 1844 2102 1856
rect 8754 1844 8760 1856
rect 8812 1844 8818 1896
rect 3510 1776 3516 1828
rect 3568 1816 3574 1828
rect 6914 1816 6920 1828
rect 3568 1788 6920 1816
rect 3568 1776 3574 1788
rect 6914 1776 6920 1788
rect 6972 1776 6978 1828
rect 9582 1776 9588 1828
rect 9640 1816 9646 1828
rect 13906 1816 13912 1828
rect 9640 1788 13912 1816
rect 9640 1776 9646 1788
rect 13906 1776 13912 1788
rect 13964 1776 13970 1828
rect 3050 1708 3056 1760
rect 3108 1748 3114 1760
rect 9306 1748 9312 1760
rect 3108 1720 9312 1748
rect 3108 1708 3114 1720
rect 9306 1708 9312 1720
rect 9364 1708 9370 1760
rect 9766 1708 9772 1760
rect 9824 1748 9830 1760
rect 14918 1748 14924 1760
rect 9824 1720 14924 1748
rect 9824 1708 9830 1720
rect 14918 1708 14924 1720
rect 14976 1708 14982 1760
rect 7558 1640 7564 1692
rect 7616 1680 7622 1692
rect 11514 1680 11520 1692
rect 7616 1652 11520 1680
rect 7616 1640 7622 1652
rect 11514 1640 11520 1652
rect 11572 1640 11578 1692
rect 4982 1572 4988 1624
rect 5040 1612 5046 1624
rect 11422 1612 11428 1624
rect 5040 1584 11428 1612
rect 5040 1572 5046 1584
rect 11422 1572 11428 1584
rect 11480 1572 11486 1624
rect 6914 1504 6920 1556
rect 6972 1544 6978 1556
rect 13078 1544 13084 1556
rect 6972 1516 13084 1544
rect 6972 1504 6978 1516
rect 8128 1488 8156 1516
rect 13078 1504 13084 1516
rect 13136 1504 13142 1556
rect 8110 1436 8116 1488
rect 8168 1436 8174 1488
rect 1394 1232 1400 1284
rect 1452 1272 1458 1284
rect 6822 1272 6828 1284
rect 1452 1244 6828 1272
rect 1452 1232 1458 1244
rect 6822 1232 6828 1244
rect 6880 1232 6886 1284
<< via1 >>
rect 9772 18028 9824 18080
rect 12348 18028 12400 18080
rect 4068 17892 4120 17944
rect 8944 17892 8996 17944
rect 10508 17960 10560 18012
rect 13360 17960 13412 18012
rect 3516 17824 3568 17876
rect 9496 17824 9548 17876
rect 12808 17892 12860 17944
rect 7840 17756 7892 17808
rect 5540 17688 5592 17740
rect 11244 17688 11296 17740
rect 14556 17756 14608 17808
rect 13176 17688 13228 17740
rect 6920 17620 6972 17672
rect 14280 17620 14332 17672
rect 5448 17552 5500 17604
rect 12716 17552 12768 17604
rect 3148 17484 3200 17536
rect 4252 17484 4304 17536
rect 7196 17484 7248 17536
rect 12900 17484 12952 17536
rect 3447 17382 3499 17434
rect 3511 17382 3563 17434
rect 3575 17382 3627 17434
rect 3639 17382 3691 17434
rect 8378 17382 8430 17434
rect 8442 17382 8494 17434
rect 8506 17382 8558 17434
rect 8570 17382 8622 17434
rect 13308 17382 13360 17434
rect 13372 17382 13424 17434
rect 13436 17382 13488 17434
rect 13500 17382 13552 17434
rect 7564 17280 7616 17332
rect 12900 17280 12952 17332
rect 2412 17212 2464 17264
rect 756 17144 808 17196
rect 1492 17119 1544 17128
rect 1492 17085 1501 17119
rect 1501 17085 1535 17119
rect 1535 17085 1544 17119
rect 1492 17076 1544 17085
rect 2136 17144 2188 17196
rect 4068 17212 4120 17264
rect 6184 17212 6236 17264
rect 10232 17212 10284 17264
rect 2412 17119 2464 17128
rect 2412 17085 2421 17119
rect 2421 17085 2455 17119
rect 2455 17085 2464 17119
rect 2412 17076 2464 17085
rect 3700 17076 3752 17128
rect 4252 17187 4304 17196
rect 4252 17153 4261 17187
rect 4261 17153 4295 17187
rect 4295 17153 4304 17187
rect 4252 17144 4304 17153
rect 7288 17144 7340 17196
rect 7472 17187 7524 17196
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 7472 17144 7524 17153
rect 10140 17144 10192 17196
rect 9496 17119 9548 17128
rect 9496 17085 9505 17119
rect 9505 17085 9539 17119
rect 9539 17085 9548 17119
rect 9496 17076 9548 17085
rect 10048 17076 10100 17128
rect 10416 17076 10468 17128
rect 3148 17008 3200 17060
rect 6276 17008 6328 17060
rect 9128 17008 9180 17060
rect 9680 17008 9732 17060
rect 12440 17076 12492 17128
rect 12900 17076 12952 17128
rect 13360 17119 13412 17128
rect 13360 17085 13369 17119
rect 13369 17085 13403 17119
rect 13403 17085 13412 17119
rect 13360 17076 13412 17085
rect 3332 16983 3384 16992
rect 3332 16949 3341 16983
rect 3341 16949 3375 16983
rect 3375 16949 3384 16983
rect 3332 16940 3384 16949
rect 4988 16983 5040 16992
rect 4988 16949 4997 16983
rect 4997 16949 5031 16983
rect 5031 16949 5040 16983
rect 4988 16940 5040 16949
rect 5632 16983 5684 16992
rect 5632 16949 5641 16983
rect 5641 16949 5675 16983
rect 5675 16949 5684 16983
rect 5632 16940 5684 16949
rect 5724 16940 5776 16992
rect 7656 16940 7708 16992
rect 8116 16983 8168 16992
rect 8116 16949 8125 16983
rect 8125 16949 8159 16983
rect 8159 16949 8168 16983
rect 8116 16940 8168 16949
rect 8576 16983 8628 16992
rect 8576 16949 8585 16983
rect 8585 16949 8619 16983
rect 8619 16949 8628 16983
rect 8576 16940 8628 16949
rect 9312 16983 9364 16992
rect 9312 16949 9321 16983
rect 9321 16949 9355 16983
rect 9355 16949 9364 16983
rect 9312 16940 9364 16949
rect 9404 16940 9456 16992
rect 10232 16940 10284 16992
rect 5912 16838 5964 16890
rect 5976 16838 6028 16890
rect 6040 16838 6092 16890
rect 6104 16838 6156 16890
rect 10843 16838 10895 16890
rect 10907 16838 10959 16890
rect 10971 16838 11023 16890
rect 11035 16838 11087 16890
rect 1676 16711 1728 16720
rect 1676 16677 1685 16711
rect 1685 16677 1719 16711
rect 1719 16677 1728 16711
rect 1676 16668 1728 16677
rect 2780 16736 2832 16788
rect 4896 16736 4948 16788
rect 2688 16643 2740 16652
rect 2688 16609 2697 16643
rect 2697 16609 2731 16643
rect 2731 16609 2740 16643
rect 2688 16600 2740 16609
rect 2780 16643 2832 16652
rect 2780 16609 2789 16643
rect 2789 16609 2823 16643
rect 2823 16609 2832 16643
rect 3884 16643 3936 16652
rect 2780 16600 2832 16609
rect 3884 16609 3893 16643
rect 3893 16609 3927 16643
rect 3927 16609 3936 16643
rect 3884 16600 3936 16609
rect 3976 16600 4028 16652
rect 3332 16532 3384 16584
rect 3700 16532 3752 16584
rect 4436 16668 4488 16720
rect 5356 16736 5408 16788
rect 6276 16779 6328 16788
rect 6276 16745 6285 16779
rect 6285 16745 6319 16779
rect 6319 16745 6328 16779
rect 6276 16736 6328 16745
rect 7840 16779 7892 16788
rect 7840 16745 7849 16779
rect 7849 16745 7883 16779
rect 7883 16745 7892 16779
rect 7840 16736 7892 16745
rect 8944 16736 8996 16788
rect 9588 16736 9640 16788
rect 4252 16600 4304 16652
rect 4528 16600 4580 16652
rect 5448 16600 5500 16652
rect 8116 16668 8168 16720
rect 12164 16736 12216 16788
rect 14280 16779 14332 16788
rect 14280 16745 14289 16779
rect 14289 16745 14323 16779
rect 14323 16745 14332 16779
rect 14280 16736 14332 16745
rect 12072 16668 12124 16720
rect 8668 16643 8720 16652
rect 8668 16609 8677 16643
rect 8677 16609 8711 16643
rect 8711 16609 8720 16643
rect 8668 16600 8720 16609
rect 8852 16600 8904 16652
rect 4712 16532 4764 16584
rect 5080 16532 5132 16584
rect 6092 16532 6144 16584
rect 7288 16532 7340 16584
rect 7748 16532 7800 16584
rect 8116 16532 8168 16584
rect 9036 16532 9088 16584
rect 1492 16464 1544 16516
rect 3792 16464 3844 16516
rect 4344 16464 4396 16516
rect 9404 16464 9456 16516
rect 2320 16396 2372 16448
rect 4436 16396 4488 16448
rect 4804 16396 4856 16448
rect 9588 16396 9640 16448
rect 10508 16600 10560 16652
rect 10968 16600 11020 16652
rect 9864 16532 9916 16584
rect 10784 16532 10836 16584
rect 12532 16600 12584 16652
rect 11428 16532 11480 16584
rect 11152 16464 11204 16516
rect 11244 16464 11296 16516
rect 11888 16464 11940 16516
rect 12808 16507 12860 16516
rect 12808 16473 12817 16507
rect 12817 16473 12851 16507
rect 12851 16473 12860 16507
rect 12808 16464 12860 16473
rect 10232 16396 10284 16448
rect 10324 16396 10376 16448
rect 14372 16396 14424 16448
rect 3447 16294 3499 16346
rect 3511 16294 3563 16346
rect 3575 16294 3627 16346
rect 3639 16294 3691 16346
rect 8378 16294 8430 16346
rect 8442 16294 8494 16346
rect 8506 16294 8558 16346
rect 8570 16294 8622 16346
rect 13308 16294 13360 16346
rect 13372 16294 13424 16346
rect 13436 16294 13488 16346
rect 13500 16294 13552 16346
rect 1124 16192 1176 16244
rect 2504 16192 2556 16244
rect 2780 16192 2832 16244
rect 3424 16124 3476 16176
rect 6644 16192 6696 16244
rect 8760 16192 8812 16244
rect 7012 16124 7064 16176
rect 1400 16056 1452 16108
rect 1768 16056 1820 16108
rect 4068 16056 4120 16108
rect 112 15988 164 16040
rect 1308 15988 1360 16040
rect 388 15920 440 15972
rect 3240 15988 3292 16040
rect 4436 15988 4488 16040
rect 3608 15963 3660 15972
rect 3608 15929 3617 15963
rect 3617 15929 3651 15963
rect 3651 15929 3660 15963
rect 3608 15920 3660 15929
rect 4252 15920 4304 15972
rect 5540 16056 5592 16108
rect 5632 16056 5684 16108
rect 6092 16099 6144 16108
rect 6092 16065 6101 16099
rect 6101 16065 6135 16099
rect 6135 16065 6144 16099
rect 7380 16099 7432 16108
rect 6092 16056 6144 16065
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 9404 16056 9456 16108
rect 9956 16192 10008 16244
rect 10784 16192 10836 16244
rect 14188 16192 14240 16244
rect 15108 16192 15160 16244
rect 16396 16192 16448 16244
rect 10508 16124 10560 16176
rect 10968 16124 11020 16176
rect 4804 16031 4856 16040
rect 4804 15997 4813 16031
rect 4813 15997 4847 16031
rect 4847 15997 4856 16031
rect 4804 15988 4856 15997
rect 4896 15988 4948 16040
rect 7288 16031 7340 16040
rect 4344 15895 4396 15904
rect 4344 15861 4353 15895
rect 4353 15861 4387 15895
rect 4387 15861 4396 15895
rect 4344 15852 4396 15861
rect 6736 15852 6788 15904
rect 7288 15997 7297 16031
rect 7297 15997 7331 16031
rect 7331 15997 7340 16031
rect 7288 15988 7340 15997
rect 9588 16031 9640 16040
rect 7840 15852 7892 15904
rect 8760 15920 8812 15972
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 10324 15988 10376 16040
rect 9772 15920 9824 15972
rect 11796 15988 11848 16040
rect 12716 15988 12768 16040
rect 13176 16031 13228 16040
rect 13176 15997 13185 16031
rect 13185 15997 13219 16031
rect 13219 15997 13228 16031
rect 13176 15988 13228 15997
rect 12348 15920 12400 15972
rect 8944 15852 8996 15904
rect 9036 15852 9088 15904
rect 11152 15852 11204 15904
rect 5912 15750 5964 15802
rect 5976 15750 6028 15802
rect 6040 15750 6092 15802
rect 6104 15750 6156 15802
rect 10843 15750 10895 15802
rect 10907 15750 10959 15802
rect 10971 15750 11023 15802
rect 11035 15750 11087 15802
rect 2964 15648 3016 15700
rect 5172 15648 5224 15700
rect 7380 15648 7432 15700
rect 8116 15691 8168 15700
rect 8116 15657 8125 15691
rect 8125 15657 8159 15691
rect 8159 15657 8168 15691
rect 8116 15648 8168 15657
rect 1308 15580 1360 15632
rect 4620 15580 4672 15632
rect 6828 15580 6880 15632
rect 6920 15580 6972 15632
rect 9220 15648 9272 15700
rect 8300 15580 8352 15632
rect 12164 15648 12216 15700
rect 1308 15444 1360 15496
rect 1492 15512 1544 15564
rect 3332 15512 3384 15564
rect 4712 15512 4764 15564
rect 2044 15444 2096 15496
rect 2596 15444 2648 15496
rect 5448 15444 5500 15496
rect 8116 15512 8168 15564
rect 9128 15512 9180 15564
rect 9680 15512 9732 15564
rect 10508 15512 10560 15564
rect 10692 15512 10744 15564
rect 10876 15555 10928 15564
rect 10876 15521 10885 15555
rect 10885 15521 10919 15555
rect 10919 15521 10928 15555
rect 10876 15512 10928 15521
rect 11520 15512 11572 15564
rect 11704 15512 11756 15564
rect 9220 15444 9272 15496
rect 2228 15376 2280 15428
rect 3240 15376 3292 15428
rect 5724 15376 5776 15428
rect 9772 15444 9824 15496
rect 4160 15308 4212 15360
rect 5264 15308 5316 15360
rect 9956 15376 10008 15428
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 7748 15308 7800 15360
rect 9404 15308 9456 15360
rect 12532 15376 12584 15428
rect 10600 15308 10652 15360
rect 13176 15444 13228 15496
rect 3447 15206 3499 15258
rect 3511 15206 3563 15258
rect 3575 15206 3627 15258
rect 3639 15206 3691 15258
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 13308 15206 13360 15258
rect 13372 15206 13424 15258
rect 13436 15206 13488 15258
rect 13500 15206 13552 15258
rect 4804 15104 4856 15156
rect 5908 15104 5960 15156
rect 8116 15104 8168 15156
rect 8944 15104 8996 15156
rect 9404 15104 9456 15156
rect 10508 15104 10560 15156
rect 12256 15104 12308 15156
rect 7840 15036 7892 15088
rect 3240 14968 3292 15020
rect 4160 15011 4212 15020
rect 4160 14977 4169 15011
rect 4169 14977 4203 15011
rect 4203 14977 4212 15011
rect 4160 14968 4212 14977
rect 4528 14968 4580 15020
rect 6736 14968 6788 15020
rect 9220 15011 9272 15020
rect 9220 14977 9229 15011
rect 9229 14977 9263 15011
rect 9263 14977 9272 15011
rect 9220 14968 9272 14977
rect 9404 14968 9456 15020
rect 10508 14968 10560 15020
rect 11336 14968 11388 15020
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 1860 14900 1912 14952
rect 4804 14900 4856 14952
rect 2964 14875 3016 14884
rect 2964 14841 2973 14875
rect 2973 14841 3007 14875
rect 3007 14841 3016 14875
rect 2964 14832 3016 14841
rect 4344 14832 4396 14884
rect 4712 14832 4764 14884
rect 6920 14832 6972 14884
rect 11428 14900 11480 14952
rect 5264 14764 5316 14816
rect 7932 14764 7984 14816
rect 9680 14832 9732 14884
rect 10784 14832 10836 14884
rect 9588 14764 9640 14816
rect 9864 14807 9916 14816
rect 9864 14773 9873 14807
rect 9873 14773 9907 14807
rect 9907 14773 9916 14807
rect 9864 14764 9916 14773
rect 10508 14764 10560 14816
rect 11152 14764 11204 14816
rect 11704 14832 11756 14884
rect 12164 14832 12216 14884
rect 14096 14832 14148 14884
rect 11612 14764 11664 14816
rect 12256 14764 12308 14816
rect 13084 14807 13136 14816
rect 13084 14773 13093 14807
rect 13093 14773 13127 14807
rect 13127 14773 13136 14807
rect 13084 14764 13136 14773
rect 13728 14807 13780 14816
rect 13728 14773 13737 14807
rect 13737 14773 13771 14807
rect 13771 14773 13780 14807
rect 13728 14764 13780 14773
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 5912 14662 5964 14714
rect 5976 14662 6028 14714
rect 6040 14662 6092 14714
rect 6104 14662 6156 14714
rect 10843 14662 10895 14714
rect 10907 14662 10959 14714
rect 10971 14662 11023 14714
rect 11035 14662 11087 14714
rect 4252 14560 4304 14612
rect 4436 14603 4488 14612
rect 4436 14569 4445 14603
rect 4445 14569 4479 14603
rect 4479 14569 4488 14603
rect 4436 14560 4488 14569
rect 4896 14603 4948 14612
rect 4896 14569 4905 14603
rect 4905 14569 4939 14603
rect 4939 14569 4948 14603
rect 4896 14560 4948 14569
rect 7472 14560 7524 14612
rect 7564 14560 7616 14612
rect 9036 14560 9088 14612
rect 9128 14560 9180 14612
rect 10140 14560 10192 14612
rect 14096 14603 14148 14612
rect 2872 14492 2924 14544
rect 4804 14467 4856 14476
rect 3056 14288 3108 14340
rect 4804 14433 4813 14467
rect 4813 14433 4847 14467
rect 4847 14433 4856 14467
rect 4804 14424 4856 14433
rect 5540 14492 5592 14544
rect 6276 14492 6328 14544
rect 6828 14492 6880 14544
rect 10784 14492 10836 14544
rect 7564 14424 7616 14476
rect 7748 14467 7800 14476
rect 7748 14433 7782 14467
rect 7782 14433 7800 14467
rect 7748 14424 7800 14433
rect 8116 14424 8168 14476
rect 4528 14356 4580 14408
rect 4620 14356 4672 14408
rect 4252 14288 4304 14340
rect 4712 14288 4764 14340
rect 5540 14356 5592 14408
rect 7380 14356 7432 14408
rect 9036 14424 9088 14476
rect 9588 14424 9640 14476
rect 9772 14424 9824 14476
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 11152 14424 11204 14476
rect 11612 14424 11664 14476
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 13636 14424 13688 14476
rect 8944 14356 8996 14408
rect 9864 14356 9916 14408
rect 10140 14399 10192 14408
rect 10140 14365 10149 14399
rect 10149 14365 10183 14399
rect 10183 14365 10192 14399
rect 10140 14356 10192 14365
rect 9220 14288 9272 14340
rect 10416 14356 10468 14408
rect 11060 14356 11112 14408
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 10784 14288 10836 14340
rect 11336 14288 11388 14340
rect 8116 14220 8168 14272
rect 8944 14220 8996 14272
rect 9128 14220 9180 14272
rect 9864 14220 9916 14272
rect 11704 14220 11756 14272
rect 15476 14220 15528 14272
rect 3447 14118 3499 14170
rect 3511 14118 3563 14170
rect 3575 14118 3627 14170
rect 3639 14118 3691 14170
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 13308 14118 13360 14170
rect 13372 14118 13424 14170
rect 13436 14118 13488 14170
rect 13500 14118 13552 14170
rect 4804 14016 4856 14068
rect 3976 13948 4028 14000
rect 8024 14016 8076 14068
rect 8116 14016 8168 14068
rect 6276 13991 6328 14000
rect 1400 13880 1452 13932
rect 4068 13880 4120 13932
rect 6276 13957 6285 13991
rect 6285 13957 6319 13991
rect 6319 13957 6328 13991
rect 6276 13948 6328 13957
rect 7840 13948 7892 14000
rect 10140 14016 10192 14068
rect 12808 14016 12860 14068
rect 13820 14016 13872 14068
rect 14188 14016 14240 14068
rect 13452 13948 13504 14000
rect 14924 13948 14976 14000
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 3332 13812 3384 13864
rect 7932 13880 7984 13932
rect 4620 13812 4672 13864
rect 6736 13812 6788 13864
rect 4436 13744 4488 13796
rect 4528 13744 4580 13796
rect 5448 13744 5500 13796
rect 7472 13812 7524 13864
rect 8668 13855 8720 13864
rect 7380 13744 7432 13796
rect 8668 13821 8677 13855
rect 8677 13821 8711 13855
rect 8711 13821 8720 13855
rect 8668 13812 8720 13821
rect 8116 13744 8168 13796
rect 9864 13812 9916 13864
rect 10232 13812 10284 13864
rect 10140 13744 10192 13796
rect 10416 13744 10468 13796
rect 10508 13744 10560 13796
rect 10692 13744 10744 13796
rect 13544 13880 13596 13932
rect 12532 13812 12584 13864
rect 13268 13812 13320 13864
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 14556 13787 14608 13796
rect 14556 13753 14565 13787
rect 14565 13753 14599 13787
rect 14599 13753 14608 13787
rect 14556 13744 14608 13753
rect 3148 13676 3200 13728
rect 7656 13676 7708 13728
rect 8668 13676 8720 13728
rect 9312 13676 9364 13728
rect 9956 13676 10008 13728
rect 11428 13676 11480 13728
rect 11612 13676 11664 13728
rect 14096 13676 14148 13728
rect 15752 13676 15804 13728
rect 5912 13574 5964 13626
rect 5976 13574 6028 13626
rect 6040 13574 6092 13626
rect 6104 13574 6156 13626
rect 10843 13574 10895 13626
rect 10907 13574 10959 13626
rect 10971 13574 11023 13626
rect 11035 13574 11087 13626
rect 4344 13472 4396 13524
rect 4436 13472 4488 13524
rect 5172 13472 5224 13524
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 8024 13515 8076 13524
rect 8024 13481 8033 13515
rect 8033 13481 8067 13515
rect 8067 13481 8076 13515
rect 8024 13472 8076 13481
rect 8300 13472 8352 13524
rect 9404 13472 9456 13524
rect 9772 13472 9824 13524
rect 13084 13472 13136 13524
rect 13268 13472 13320 13524
rect 3332 13404 3384 13456
rect 2136 13268 2188 13320
rect 2780 13268 2832 13320
rect 2596 13200 2648 13252
rect 2872 13132 2924 13184
rect 5264 13404 5316 13456
rect 5540 13404 5592 13456
rect 6276 13404 6328 13456
rect 7472 13404 7524 13456
rect 4436 13336 4488 13388
rect 5816 13336 5868 13388
rect 6736 13336 6788 13388
rect 6828 13336 6880 13388
rect 8300 13336 8352 13388
rect 8392 13379 8444 13388
rect 8392 13345 8401 13379
rect 8401 13345 8435 13379
rect 8435 13345 8444 13379
rect 9404 13379 9456 13388
rect 8392 13336 8444 13345
rect 9404 13345 9413 13379
rect 9413 13345 9447 13379
rect 9447 13345 9456 13379
rect 9404 13336 9456 13345
rect 9680 13404 9732 13456
rect 11060 13404 11112 13456
rect 9956 13379 10008 13388
rect 9956 13345 9990 13379
rect 9990 13345 10008 13379
rect 9956 13336 10008 13345
rect 10416 13336 10468 13388
rect 8944 13268 8996 13320
rect 12532 13336 12584 13388
rect 12624 13336 12676 13388
rect 12808 13336 12860 13388
rect 13912 13379 13964 13388
rect 13912 13345 13921 13379
rect 13921 13345 13955 13379
rect 13955 13345 13964 13379
rect 13912 13336 13964 13345
rect 11336 13268 11388 13320
rect 13544 13268 13596 13320
rect 13728 13268 13780 13320
rect 7472 13132 7524 13184
rect 7656 13132 7708 13184
rect 9220 13175 9272 13184
rect 9220 13141 9229 13175
rect 9229 13141 9263 13175
rect 9263 13141 9272 13175
rect 9220 13132 9272 13141
rect 9312 13132 9364 13184
rect 11612 13200 11664 13252
rect 11704 13200 11756 13252
rect 12808 13200 12860 13252
rect 13912 13200 13964 13252
rect 14280 13200 14332 13252
rect 14188 13132 14240 13184
rect 15108 13132 15160 13184
rect 3447 13030 3499 13082
rect 3511 13030 3563 13082
rect 3575 13030 3627 13082
rect 3639 13030 3691 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 13308 13030 13360 13082
rect 13372 13030 13424 13082
rect 13436 13030 13488 13082
rect 13500 13030 13552 13082
rect 3056 12928 3108 12980
rect 6276 12971 6328 12980
rect 2412 12860 2464 12912
rect 6276 12937 6285 12971
rect 6285 12937 6319 12971
rect 6319 12937 6328 12971
rect 6276 12928 6328 12937
rect 2504 12835 2556 12844
rect 2504 12801 2513 12835
rect 2513 12801 2547 12835
rect 2547 12801 2556 12835
rect 2504 12792 2556 12801
rect 6828 12860 6880 12912
rect 8944 12928 8996 12980
rect 9312 12928 9364 12980
rect 8484 12860 8536 12912
rect 9680 12928 9732 12980
rect 9956 12860 10008 12912
rect 10232 12860 10284 12912
rect 11428 12860 11480 12912
rect 12532 12860 12584 12912
rect 14280 12860 14332 12912
rect 15384 12860 15436 12912
rect 2596 12724 2648 12776
rect 4620 12724 4672 12776
rect 3516 12656 3568 12708
rect 5172 12767 5224 12776
rect 5172 12733 5206 12767
rect 5206 12733 5224 12767
rect 5172 12724 5224 12733
rect 7840 12792 7892 12844
rect 8668 12835 8720 12844
rect 5264 12656 5316 12708
rect 5540 12656 5592 12708
rect 6920 12724 6972 12776
rect 8116 12724 8168 12776
rect 8668 12801 8677 12835
rect 8677 12801 8711 12835
rect 8711 12801 8720 12835
rect 8668 12792 8720 12801
rect 10692 12792 10744 12844
rect 12808 12792 12860 12844
rect 13636 12792 13688 12844
rect 9220 12724 9272 12776
rect 9312 12724 9364 12776
rect 11152 12724 11204 12776
rect 14188 12792 14240 12844
rect 15016 12792 15068 12844
rect 14832 12767 14884 12776
rect 14832 12733 14841 12767
rect 14841 12733 14875 12767
rect 14875 12733 14884 12767
rect 14832 12724 14884 12733
rect 7380 12656 7432 12708
rect 7564 12588 7616 12640
rect 8208 12656 8260 12708
rect 9772 12656 9824 12708
rect 9588 12588 9640 12640
rect 9956 12588 10008 12640
rect 11336 12656 11388 12708
rect 15752 12656 15804 12708
rect 11704 12631 11756 12640
rect 11704 12597 11713 12631
rect 11713 12597 11747 12631
rect 11747 12597 11756 12631
rect 11704 12588 11756 12597
rect 12072 12588 12124 12640
rect 12256 12588 12308 12640
rect 12808 12631 12860 12640
rect 12808 12597 12817 12631
rect 12817 12597 12851 12631
rect 12851 12597 12860 12631
rect 12808 12588 12860 12597
rect 14004 12588 14056 12640
rect 14832 12588 14884 12640
rect 15016 12631 15068 12640
rect 15016 12597 15025 12631
rect 15025 12597 15059 12631
rect 15059 12597 15068 12631
rect 15016 12588 15068 12597
rect 5912 12486 5964 12538
rect 5976 12486 6028 12538
rect 6040 12486 6092 12538
rect 6104 12486 6156 12538
rect 10843 12486 10895 12538
rect 10907 12486 10959 12538
rect 10971 12486 11023 12538
rect 11035 12486 11087 12538
rect 2780 12427 2832 12436
rect 2780 12393 2789 12427
rect 2789 12393 2823 12427
rect 2823 12393 2832 12427
rect 2780 12384 2832 12393
rect 3056 12384 3108 12436
rect 6644 12384 6696 12436
rect 6920 12427 6972 12436
rect 6920 12393 6929 12427
rect 6929 12393 6963 12427
rect 6963 12393 6972 12427
rect 6920 12384 6972 12393
rect 2596 12316 2648 12368
rect 4712 12359 4764 12368
rect 4712 12325 4721 12359
rect 4721 12325 4755 12359
rect 4755 12325 4764 12359
rect 4712 12316 4764 12325
rect 3148 12248 3200 12300
rect 4620 12248 4672 12300
rect 5540 12291 5592 12300
rect 5540 12257 5549 12291
rect 5549 12257 5583 12291
rect 5583 12257 5592 12291
rect 5540 12248 5592 12257
rect 5724 12316 5776 12368
rect 6552 12316 6604 12368
rect 7748 12316 7800 12368
rect 9496 12384 9548 12436
rect 11152 12384 11204 12436
rect 11704 12384 11756 12436
rect 12532 12427 12584 12436
rect 12532 12393 12541 12427
rect 12541 12393 12575 12427
rect 12575 12393 12584 12427
rect 12532 12384 12584 12393
rect 9404 12291 9456 12300
rect 4068 12180 4120 12232
rect 3056 12112 3108 12164
rect 3516 12112 3568 12164
rect 4896 12223 4948 12232
rect 4896 12189 4905 12223
rect 4905 12189 4939 12223
rect 4939 12189 4948 12223
rect 7380 12223 7432 12232
rect 4896 12180 4948 12189
rect 7380 12189 7389 12223
rect 7389 12189 7423 12223
rect 7423 12189 7432 12223
rect 7380 12180 7432 12189
rect 9404 12257 9413 12291
rect 9413 12257 9447 12291
rect 9447 12257 9456 12291
rect 9404 12248 9456 12257
rect 9588 12316 9640 12368
rect 10232 12316 10284 12368
rect 10876 12316 10928 12368
rect 10968 12316 11020 12368
rect 11336 12359 11388 12368
rect 11060 12248 11112 12300
rect 11336 12325 11345 12359
rect 11345 12325 11379 12359
rect 11379 12325 11388 12359
rect 11336 12316 11388 12325
rect 12256 12316 12308 12368
rect 12348 12316 12400 12368
rect 9864 12180 9916 12232
rect 10140 12223 10192 12232
rect 10140 12189 10149 12223
rect 10149 12189 10183 12223
rect 10183 12189 10192 12223
rect 10140 12180 10192 12189
rect 10232 12180 10284 12232
rect 11980 12248 12032 12300
rect 13452 12291 13504 12300
rect 13452 12257 13461 12291
rect 13461 12257 13495 12291
rect 13495 12257 13504 12291
rect 13452 12248 13504 12257
rect 13176 12180 13228 12232
rect 14556 12248 14608 12300
rect 14832 12248 14884 12300
rect 15384 12180 15436 12232
rect 5540 12112 5592 12164
rect 8392 12112 8444 12164
rect 14556 12112 14608 12164
rect 14740 12112 14792 12164
rect 2872 12044 2924 12096
rect 4344 12087 4396 12096
rect 4344 12053 4353 12087
rect 4353 12053 4387 12087
rect 4387 12053 4396 12087
rect 4344 12044 4396 12053
rect 5448 12044 5500 12096
rect 8944 12044 8996 12096
rect 9496 12044 9548 12096
rect 9680 12087 9732 12096
rect 9680 12053 9689 12087
rect 9689 12053 9723 12087
rect 9723 12053 9732 12087
rect 9680 12044 9732 12053
rect 9864 12044 9916 12096
rect 10048 12044 10100 12096
rect 10140 12044 10192 12096
rect 11704 12044 11756 12096
rect 12256 12044 12308 12096
rect 12808 12044 12860 12096
rect 14096 12044 14148 12096
rect 3447 11942 3499 11994
rect 3511 11942 3563 11994
rect 3575 11942 3627 11994
rect 3639 11942 3691 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 13308 11942 13360 11994
rect 13372 11942 13424 11994
rect 13436 11942 13488 11994
rect 13500 11942 13552 11994
rect 1768 11840 1820 11892
rect 3332 11840 3384 11892
rect 1308 11772 1360 11824
rect 3976 11772 4028 11824
rect 3056 11704 3108 11756
rect 3332 11704 3384 11756
rect 1768 11636 1820 11688
rect 2872 11679 2924 11688
rect 2872 11645 2881 11679
rect 2881 11645 2915 11679
rect 2915 11645 2924 11679
rect 2872 11636 2924 11645
rect 8668 11840 8720 11892
rect 11060 11840 11112 11892
rect 13176 11840 13228 11892
rect 8944 11772 8996 11824
rect 4252 11747 4304 11756
rect 4252 11713 4261 11747
rect 4261 11713 4295 11747
rect 4295 11713 4304 11747
rect 4252 11704 4304 11713
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 8668 11704 8720 11756
rect 11428 11772 11480 11824
rect 12716 11772 12768 11824
rect 10876 11747 10928 11756
rect 4896 11679 4948 11688
rect 4896 11645 4905 11679
rect 4905 11645 4939 11679
rect 4939 11645 4948 11679
rect 4896 11636 4948 11645
rect 5724 11636 5776 11688
rect 7656 11679 7708 11688
rect 7656 11645 7690 11679
rect 7690 11645 7708 11679
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 11244 11704 11296 11756
rect 7656 11636 7708 11645
rect 10232 11636 10284 11688
rect 10508 11636 10560 11688
rect 4252 11568 4304 11620
rect 5172 11611 5224 11620
rect 5172 11577 5206 11611
rect 5206 11577 5224 11611
rect 5172 11568 5224 11577
rect 3056 11500 3108 11552
rect 8668 11568 8720 11620
rect 9588 11611 9640 11620
rect 9588 11577 9597 11611
rect 9597 11577 9631 11611
rect 9631 11577 9640 11611
rect 9588 11568 9640 11577
rect 6920 11500 6972 11552
rect 8944 11500 8996 11552
rect 9220 11543 9272 11552
rect 9220 11509 9229 11543
rect 9229 11509 9263 11543
rect 9263 11509 9272 11543
rect 9220 11500 9272 11509
rect 9864 11500 9916 11552
rect 10232 11500 10284 11552
rect 13544 11704 13596 11756
rect 14924 11704 14976 11756
rect 13176 11568 13228 11620
rect 13728 11636 13780 11688
rect 13820 11636 13872 11688
rect 14004 11568 14056 11620
rect 16396 11568 16448 11620
rect 12348 11500 12400 11552
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 6104 11398 6156 11450
rect 10843 11398 10895 11450
rect 10907 11398 10959 11450
rect 10971 11398 11023 11450
rect 11035 11398 11087 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 4528 11296 4580 11348
rect 8760 11296 8812 11348
rect 9220 11296 9272 11348
rect 10140 11339 10192 11348
rect 9588 11228 9640 11280
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 11704 11296 11756 11348
rect 13084 11296 13136 11348
rect 1952 11203 2004 11212
rect 1952 11169 1961 11203
rect 1961 11169 1995 11203
rect 1995 11169 2004 11203
rect 1952 11160 2004 11169
rect 2412 11160 2464 11212
rect 2504 11160 2556 11212
rect 5632 11160 5684 11212
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 6920 11160 6972 11212
rect 7748 11160 7800 11212
rect 8944 11160 8996 11212
rect 1676 11092 1728 11144
rect 3240 11135 3292 11144
rect 3240 11101 3249 11135
rect 3249 11101 3283 11135
rect 3283 11101 3292 11135
rect 3240 11092 3292 11101
rect 4436 11092 4488 11144
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 5264 11092 5316 11101
rect 5448 11092 5500 11144
rect 7380 11092 7432 11144
rect 9036 11092 9088 11144
rect 9128 11092 9180 11144
rect 9312 11092 9364 11144
rect 10692 11160 10744 11212
rect 13728 11228 13780 11280
rect 11060 11160 11112 11212
rect 11336 11160 11388 11212
rect 11704 11160 11756 11212
rect 11888 11160 11940 11212
rect 12440 11203 12492 11212
rect 12440 11169 12449 11203
rect 12449 11169 12483 11203
rect 12483 11169 12492 11203
rect 12440 11160 12492 11169
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 4528 11024 4580 11076
rect 9588 11024 9640 11076
rect 9772 11024 9824 11076
rect 9956 11024 10008 11076
rect 10508 11024 10560 11076
rect 10968 11024 11020 11076
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 12716 11024 12768 11076
rect 13544 11024 13596 11076
rect 14832 11024 14884 11076
rect 1584 10956 1636 11008
rect 2688 10956 2740 11008
rect 6736 10956 6788 11008
rect 7196 10999 7248 11008
rect 7196 10965 7205 10999
rect 7205 10965 7239 10999
rect 7239 10965 7248 10999
rect 7196 10956 7248 10965
rect 7656 10956 7708 11008
rect 9036 10999 9088 11008
rect 9036 10965 9045 10999
rect 9045 10965 9079 10999
rect 9079 10965 9088 10999
rect 9036 10956 9088 10965
rect 10784 10956 10836 11008
rect 11888 10956 11940 11008
rect 15292 10956 15344 11008
rect 3447 10854 3499 10906
rect 3511 10854 3563 10906
rect 3575 10854 3627 10906
rect 3639 10854 3691 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 13308 10854 13360 10906
rect 13372 10854 13424 10906
rect 13436 10854 13488 10906
rect 13500 10854 13552 10906
rect 3148 10752 3200 10804
rect 2688 10616 2740 10668
rect 5172 10752 5224 10804
rect 5540 10752 5592 10804
rect 9404 10752 9456 10804
rect 11060 10752 11112 10804
rect 11336 10752 11388 10804
rect 13636 10795 13688 10804
rect 13636 10761 13645 10795
rect 13645 10761 13679 10795
rect 13679 10761 13688 10795
rect 13636 10752 13688 10761
rect 10692 10684 10744 10736
rect 4436 10616 4488 10668
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 7932 10616 7984 10668
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 8208 10591 8260 10600
rect 8208 10557 8217 10591
rect 8217 10557 8251 10591
rect 8251 10557 8260 10591
rect 8208 10548 8260 10557
rect 10140 10616 10192 10668
rect 10508 10616 10560 10668
rect 10600 10616 10652 10668
rect 10968 10684 11020 10736
rect 11520 10684 11572 10736
rect 11060 10616 11112 10668
rect 11336 10616 11388 10668
rect 11888 10684 11940 10736
rect 12532 10616 12584 10668
rect 1860 10523 1912 10532
rect 1860 10489 1869 10523
rect 1869 10489 1903 10523
rect 1903 10489 1912 10523
rect 1860 10480 1912 10489
rect 3332 10480 3384 10532
rect 2780 10412 2832 10464
rect 3148 10412 3200 10464
rect 3884 10412 3936 10464
rect 4620 10480 4672 10532
rect 7012 10480 7064 10532
rect 7380 10480 7432 10532
rect 9036 10480 9088 10532
rect 6368 10412 6420 10464
rect 9772 10412 9824 10464
rect 10416 10480 10468 10532
rect 12440 10548 12492 10600
rect 11888 10480 11940 10532
rect 13636 10616 13688 10668
rect 14372 10548 14424 10600
rect 16764 10548 16816 10600
rect 14648 10480 14700 10532
rect 9956 10412 10008 10464
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 14372 10412 14424 10464
rect 15016 10455 15068 10464
rect 15016 10421 15025 10455
rect 15025 10421 15059 10455
rect 15059 10421 15068 10455
rect 15016 10412 15068 10421
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 6104 10310 6156 10362
rect 10843 10310 10895 10362
rect 10907 10310 10959 10362
rect 10971 10310 11023 10362
rect 11035 10310 11087 10362
rect 2504 10208 2556 10260
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 2780 10208 2832 10217
rect 3792 10208 3844 10260
rect 4068 10208 4120 10260
rect 4252 10251 4304 10260
rect 4252 10217 4261 10251
rect 4261 10217 4295 10251
rect 4295 10217 4304 10251
rect 4252 10208 4304 10217
rect 4344 10208 4396 10260
rect 4528 10140 4580 10192
rect 11336 10251 11388 10260
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 11612 10208 11664 10260
rect 11796 10208 11848 10260
rect 13728 10208 13780 10260
rect 2780 10072 2832 10124
rect 7472 10140 7524 10192
rect 7656 10140 7708 10192
rect 9864 10140 9916 10192
rect 10692 10140 10744 10192
rect 11060 10140 11112 10192
rect 11520 10140 11572 10192
rect 12072 10140 12124 10192
rect 13452 10140 13504 10192
rect 13820 10140 13872 10192
rect 5724 10115 5776 10124
rect 5724 10081 5758 10115
rect 5758 10081 5776 10115
rect 2872 10004 2924 10056
rect 5724 10072 5776 10081
rect 7196 10072 7248 10124
rect 7288 10115 7340 10124
rect 7288 10081 7297 10115
rect 7297 10081 7331 10115
rect 7331 10081 7340 10115
rect 9312 10115 9364 10124
rect 7288 10072 7340 10081
rect 9312 10081 9321 10115
rect 9321 10081 9355 10115
rect 9355 10081 9364 10115
rect 9312 10072 9364 10081
rect 10140 10115 10192 10124
rect 3884 10004 3936 10056
rect 4620 10004 4672 10056
rect 4528 9936 4580 9988
rect 4896 10004 4948 10056
rect 6828 10004 6880 10056
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 9864 10004 9916 10056
rect 10416 10072 10468 10124
rect 10508 10072 10560 10124
rect 12348 10072 12400 10124
rect 13360 10072 13412 10124
rect 13728 10115 13780 10124
rect 13728 10081 13737 10115
rect 13737 10081 13771 10115
rect 13771 10081 13780 10115
rect 15660 10140 15712 10192
rect 13728 10072 13780 10081
rect 14188 10072 14240 10124
rect 2596 9868 2648 9920
rect 3792 9868 3844 9920
rect 4896 9868 4948 9920
rect 8024 9868 8076 9920
rect 10416 9936 10468 9988
rect 11888 10004 11940 10056
rect 13544 10004 13596 10056
rect 13728 9936 13780 9988
rect 14648 9979 14700 9988
rect 14648 9945 14657 9979
rect 14657 9945 14691 9979
rect 14691 9945 14700 9979
rect 14648 9936 14700 9945
rect 9404 9868 9456 9920
rect 9496 9868 9548 9920
rect 9772 9868 9824 9920
rect 14004 9868 14056 9920
rect 14924 9868 14976 9920
rect 3447 9766 3499 9818
rect 3511 9766 3563 9818
rect 3575 9766 3627 9818
rect 3639 9766 3691 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 13308 9766 13360 9818
rect 13372 9766 13424 9818
rect 13436 9766 13488 9818
rect 13500 9766 13552 9818
rect 2872 9664 2924 9716
rect 5172 9707 5224 9716
rect 2688 9596 2740 9648
rect 3700 9596 3752 9648
rect 5172 9673 5181 9707
rect 5181 9673 5215 9707
rect 5215 9673 5224 9707
rect 5172 9664 5224 9673
rect 5264 9664 5316 9716
rect 2320 9528 2372 9580
rect 2596 9571 2648 9580
rect 2596 9537 2605 9571
rect 2605 9537 2639 9571
rect 2639 9537 2648 9571
rect 2596 9528 2648 9537
rect 2872 9460 2924 9512
rect 2964 9460 3016 9512
rect 3240 9460 3292 9512
rect 2504 9435 2556 9444
rect 2504 9401 2513 9435
rect 2513 9401 2547 9435
rect 2547 9401 2556 9435
rect 2504 9392 2556 9401
rect 3792 9503 3844 9512
rect 3792 9469 3801 9503
rect 3801 9469 3835 9503
rect 3835 9469 3844 9503
rect 3792 9460 3844 9469
rect 4988 9528 5040 9580
rect 9128 9596 9180 9648
rect 10232 9596 10284 9648
rect 10692 9596 10744 9648
rect 11704 9664 11756 9716
rect 12532 9664 12584 9716
rect 6828 9571 6880 9580
rect 4528 9460 4580 9512
rect 4804 9460 4856 9512
rect 3884 9392 3936 9444
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 8116 9528 8168 9580
rect 8760 9528 8812 9580
rect 8944 9528 8996 9580
rect 9404 9528 9456 9580
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 10508 9528 10560 9580
rect 11244 9528 11296 9580
rect 13452 9596 13504 9648
rect 5816 9460 5868 9512
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 4988 9324 5040 9376
rect 5632 9392 5684 9444
rect 5724 9392 5776 9444
rect 6276 9392 6328 9444
rect 7196 9392 7248 9444
rect 8392 9392 8444 9444
rect 9680 9460 9732 9512
rect 11152 9460 11204 9512
rect 11428 9503 11480 9512
rect 11428 9469 11437 9503
rect 11437 9469 11471 9503
rect 11471 9469 11480 9503
rect 11428 9460 11480 9469
rect 7380 9324 7432 9376
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 9772 9392 9824 9444
rect 10784 9392 10836 9444
rect 9680 9324 9732 9376
rect 10232 9324 10284 9376
rect 10508 9324 10560 9376
rect 11704 9392 11756 9444
rect 13912 9528 13964 9580
rect 14648 9664 14700 9716
rect 15200 9664 15252 9716
rect 13176 9460 13228 9512
rect 11336 9324 11388 9376
rect 11428 9324 11480 9376
rect 13268 9392 13320 9444
rect 11980 9324 12032 9376
rect 12256 9324 12308 9376
rect 13176 9324 13228 9376
rect 13728 9392 13780 9444
rect 14372 9460 14424 9512
rect 13912 9324 13964 9376
rect 15016 9367 15068 9376
rect 15016 9333 15025 9367
rect 15025 9333 15059 9367
rect 15059 9333 15068 9367
rect 15016 9324 15068 9333
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 6104 9222 6156 9274
rect 10843 9222 10895 9274
rect 10907 9222 10959 9274
rect 10971 9222 11023 9274
rect 11035 9222 11087 9274
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 3332 9120 3384 9172
rect 2688 9052 2740 9104
rect 2504 8984 2556 9036
rect 2780 8984 2832 9036
rect 3700 8984 3752 9036
rect 7472 9120 7524 9172
rect 7564 9120 7616 9172
rect 8024 9120 8076 9172
rect 4620 9095 4672 9104
rect 4620 9061 4629 9095
rect 4629 9061 4663 9095
rect 4663 9061 4672 9095
rect 4620 9052 4672 9061
rect 5172 9052 5224 9104
rect 4436 8984 4488 9036
rect 5080 8984 5132 9036
rect 7840 8984 7892 9036
rect 8116 9027 8168 9036
rect 8116 8993 8125 9027
rect 8125 8993 8159 9027
rect 8159 8993 8168 9027
rect 8116 8984 8168 8993
rect 1952 8780 2004 8832
rect 3792 8848 3844 8900
rect 4436 8848 4488 8900
rect 4528 8780 4580 8832
rect 7012 8916 7064 8968
rect 7748 8916 7800 8968
rect 8484 8984 8536 9036
rect 8760 9052 8812 9104
rect 9772 9052 9824 9104
rect 10324 9120 10376 9172
rect 11336 9163 11388 9172
rect 11336 9129 11345 9163
rect 11345 9129 11379 9163
rect 11379 9129 11388 9163
rect 11336 9120 11388 9129
rect 10140 9095 10192 9104
rect 10140 9061 10149 9095
rect 10149 9061 10183 9095
rect 10183 9061 10192 9095
rect 10140 9052 10192 9061
rect 10784 9052 10836 9104
rect 12808 9120 12860 9172
rect 13176 9120 13228 9172
rect 13452 9120 13504 9172
rect 11244 9027 11296 9036
rect 8392 8959 8444 8968
rect 8392 8925 8401 8959
rect 8401 8925 8435 8959
rect 8435 8925 8444 8959
rect 8392 8916 8444 8925
rect 4804 8848 4856 8900
rect 10048 8916 10100 8968
rect 11244 8993 11253 9027
rect 11253 8993 11287 9027
rect 11287 8993 11296 9027
rect 11244 8984 11296 8993
rect 12256 9052 12308 9104
rect 15200 9052 15252 9104
rect 12532 9027 12584 9036
rect 12532 8993 12541 9027
rect 12541 8993 12575 9027
rect 12575 8993 12584 9027
rect 12532 8984 12584 8993
rect 13176 8984 13228 9036
rect 14280 8984 14332 9036
rect 11336 8916 11388 8968
rect 7380 8780 7432 8832
rect 7472 8780 7524 8832
rect 10968 8848 11020 8900
rect 13728 8848 13780 8900
rect 9680 8823 9732 8832
rect 9680 8789 9689 8823
rect 9689 8789 9723 8823
rect 9723 8789 9732 8823
rect 9680 8780 9732 8789
rect 9772 8780 9824 8832
rect 11060 8780 11112 8832
rect 12624 8780 12676 8832
rect 13820 8780 13872 8832
rect 3447 8678 3499 8730
rect 3511 8678 3563 8730
rect 3575 8678 3627 8730
rect 3639 8678 3691 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 13308 8678 13360 8730
rect 13372 8678 13424 8730
rect 13436 8678 13488 8730
rect 13500 8678 13552 8730
rect 2964 8483 3016 8492
rect 2964 8449 2973 8483
rect 2973 8449 3007 8483
rect 3007 8449 3016 8483
rect 2964 8440 3016 8449
rect 3516 8440 3568 8492
rect 3792 8372 3844 8424
rect 1216 8304 1268 8356
rect 1308 8236 1360 8288
rect 3332 8304 3384 8356
rect 3976 8304 4028 8356
rect 9588 8576 9640 8628
rect 9864 8576 9916 8628
rect 10324 8576 10376 8628
rect 11060 8619 11112 8628
rect 11060 8585 11069 8619
rect 11069 8585 11103 8619
rect 11103 8585 11112 8619
rect 11060 8576 11112 8585
rect 11244 8576 11296 8628
rect 13084 8576 13136 8628
rect 6276 8551 6328 8560
rect 6276 8517 6285 8551
rect 6285 8517 6319 8551
rect 6319 8517 6328 8551
rect 6276 8508 6328 8517
rect 7840 8508 7892 8560
rect 8208 8508 8260 8560
rect 8944 8508 8996 8560
rect 4804 8440 4856 8492
rect 7932 8440 7984 8492
rect 10968 8508 11020 8560
rect 11612 8508 11664 8560
rect 12900 8508 12952 8560
rect 9772 8440 9824 8492
rect 10048 8440 10100 8492
rect 11336 8440 11388 8492
rect 14464 8508 14516 8560
rect 4712 8372 4764 8424
rect 5172 8415 5224 8424
rect 5172 8381 5206 8415
rect 5206 8381 5224 8415
rect 5172 8372 5224 8381
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 6368 8304 6420 8356
rect 2320 8236 2372 8288
rect 2596 8236 2648 8288
rect 7012 8304 7064 8356
rect 7932 8304 7984 8356
rect 7840 8236 7892 8288
rect 8760 8304 8812 8356
rect 13728 8372 13780 8424
rect 13912 8372 13964 8424
rect 14188 8372 14240 8424
rect 14556 8372 14608 8424
rect 8300 8236 8352 8288
rect 9036 8279 9088 8288
rect 9036 8245 9045 8279
rect 9045 8245 9079 8279
rect 9079 8245 9088 8279
rect 9036 8236 9088 8245
rect 9128 8279 9180 8288
rect 9128 8245 9137 8279
rect 9137 8245 9171 8279
rect 9171 8245 9180 8279
rect 9128 8236 9180 8245
rect 9496 8236 9548 8288
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 10232 8279 10284 8288
rect 10232 8245 10241 8279
rect 10241 8245 10275 8279
rect 10275 8245 10284 8279
rect 10232 8236 10284 8245
rect 11336 8236 11388 8288
rect 11520 8236 11572 8288
rect 11796 8236 11848 8288
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 13084 8304 13136 8356
rect 14280 8304 14332 8356
rect 15568 8236 15620 8288
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 6104 8134 6156 8186
rect 10843 8134 10895 8186
rect 10907 8134 10959 8186
rect 10971 8134 11023 8186
rect 11035 8134 11087 8186
rect 2688 8032 2740 8084
rect 5172 8032 5224 8084
rect 8024 8032 8076 8084
rect 9404 8032 9456 8084
rect 9588 8032 9640 8084
rect 9864 8032 9916 8084
rect 11152 8032 11204 8084
rect 11336 8032 11388 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 2688 7896 2740 7948
rect 5632 7896 5684 7948
rect 6000 7896 6052 7948
rect 7840 7896 7892 7948
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 3240 7871 3292 7880
rect 3240 7837 3249 7871
rect 3249 7837 3283 7871
rect 3283 7837 3292 7871
rect 3240 7828 3292 7837
rect 3792 7828 3844 7880
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 3976 7760 4028 7812
rect 2596 7692 2648 7744
rect 5448 7735 5500 7744
rect 5448 7701 5457 7735
rect 5457 7701 5491 7735
rect 5491 7701 5500 7735
rect 5448 7692 5500 7701
rect 7196 7692 7248 7744
rect 7472 7692 7524 7744
rect 9220 7760 9272 7812
rect 10784 7896 10836 7948
rect 11796 7964 11848 8016
rect 9496 7828 9548 7880
rect 11060 7828 11112 7880
rect 11152 7828 11204 7880
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 8668 7692 8720 7744
rect 9036 7692 9088 7744
rect 9864 7692 9916 7744
rect 10048 7760 10100 7812
rect 10968 7760 11020 7812
rect 12256 7896 12308 7948
rect 13176 7896 13228 7948
rect 14004 7896 14056 7948
rect 12900 7828 12952 7880
rect 12256 7760 12308 7812
rect 13268 7803 13320 7812
rect 13268 7769 13277 7803
rect 13277 7769 13311 7803
rect 13311 7769 13320 7803
rect 13268 7760 13320 7769
rect 11244 7692 11296 7744
rect 12072 7692 12124 7744
rect 14188 7828 14240 7880
rect 14004 7760 14056 7812
rect 14924 7760 14976 7812
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 3447 7590 3499 7642
rect 3511 7590 3563 7642
rect 3575 7590 3627 7642
rect 3639 7590 3691 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 13308 7590 13360 7642
rect 13372 7590 13424 7642
rect 13436 7590 13488 7642
rect 13500 7590 13552 7642
rect 1768 7488 1820 7540
rect 2228 7488 2280 7540
rect 6000 7488 6052 7540
rect 7196 7488 7248 7540
rect 4160 7420 4212 7472
rect 4896 7420 4948 7472
rect 7932 7420 7984 7472
rect 9864 7420 9916 7472
rect 2320 7395 2372 7404
rect 2320 7361 2329 7395
rect 2329 7361 2363 7395
rect 2363 7361 2372 7395
rect 2320 7352 2372 7361
rect 2320 7216 2372 7268
rect 2688 7216 2740 7268
rect 2504 7148 2556 7200
rect 6276 7352 6328 7404
rect 4712 7284 4764 7336
rect 5724 7284 5776 7336
rect 5908 7284 5960 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 8116 7352 8168 7404
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 10600 7352 10652 7404
rect 14188 7488 14240 7540
rect 11152 7420 11204 7472
rect 11060 7395 11112 7404
rect 11060 7361 11069 7395
rect 11069 7361 11103 7395
rect 11103 7361 11112 7395
rect 11060 7352 11112 7361
rect 8392 7216 8444 7268
rect 9680 7216 9732 7268
rect 10600 7216 10652 7268
rect 12716 7352 12768 7404
rect 12808 7284 12860 7336
rect 13636 7352 13688 7404
rect 13728 7284 13780 7336
rect 5632 7148 5684 7200
rect 5724 7148 5776 7200
rect 6276 7191 6328 7200
rect 6276 7157 6285 7191
rect 6285 7157 6319 7191
rect 6319 7157 6328 7191
rect 6276 7148 6328 7157
rect 6828 7148 6880 7200
rect 7472 7148 7524 7200
rect 7564 7148 7616 7200
rect 14924 7216 14976 7268
rect 12532 7148 12584 7200
rect 12808 7191 12860 7200
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 12808 7148 12860 7157
rect 13636 7191 13688 7200
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 14556 7148 14608 7200
rect 15016 7191 15068 7200
rect 15016 7157 15025 7191
rect 15025 7157 15059 7191
rect 15059 7157 15068 7191
rect 15016 7148 15068 7157
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 6104 7046 6156 7098
rect 10843 7046 10895 7098
rect 10907 7046 10959 7098
rect 10971 7046 11023 7098
rect 11035 7046 11087 7098
rect 2688 6944 2740 6996
rect 2780 6944 2832 6996
rect 3792 6944 3844 6996
rect 6276 6944 6328 6996
rect 4896 6876 4948 6928
rect 5356 6876 5408 6928
rect 8392 6944 8444 6996
rect 9496 6944 9548 6996
rect 10048 6987 10100 6996
rect 10048 6953 10057 6987
rect 10057 6953 10091 6987
rect 10091 6953 10100 6987
rect 10048 6944 10100 6953
rect 1308 6808 1360 6860
rect 4160 6808 4212 6860
rect 5080 6851 5132 6860
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 3976 6740 4028 6792
rect 5080 6817 5089 6851
rect 5089 6817 5123 6851
rect 5123 6817 5132 6851
rect 5080 6808 5132 6817
rect 4712 6740 4764 6792
rect 5540 6672 5592 6724
rect 1400 6604 1452 6656
rect 2504 6604 2556 6656
rect 5264 6604 5316 6656
rect 10600 6876 10652 6928
rect 11152 6944 11204 6996
rect 12808 6944 12860 6996
rect 7472 6808 7524 6860
rect 7840 6851 7892 6860
rect 7840 6817 7863 6851
rect 7863 6817 7892 6851
rect 7840 6808 7892 6817
rect 9128 6808 9180 6860
rect 11520 6876 11572 6928
rect 10048 6740 10100 6792
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 11704 6808 11756 6860
rect 13728 6876 13780 6928
rect 11152 6740 11204 6792
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 14372 6808 14424 6860
rect 14648 6808 14700 6860
rect 11428 6740 11480 6749
rect 12716 6740 12768 6792
rect 7932 6604 7984 6656
rect 8208 6604 8260 6656
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 10140 6604 10192 6656
rect 10968 6604 11020 6656
rect 13820 6672 13872 6724
rect 11704 6604 11756 6656
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 3240 6400 3292 6452
rect 4620 6400 4672 6452
rect 5172 6400 5224 6452
rect 5264 6400 5316 6452
rect 10048 6400 10100 6452
rect 10140 6400 10192 6452
rect 6276 6375 6328 6384
rect 2136 6196 2188 6248
rect 6276 6341 6285 6375
rect 6285 6341 6319 6375
rect 6319 6341 6328 6375
rect 6276 6332 6328 6341
rect 7932 6332 7984 6384
rect 4712 6264 4764 6316
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 9772 6332 9824 6384
rect 11704 6332 11756 6384
rect 13452 6332 13504 6384
rect 2228 6171 2280 6180
rect 2228 6137 2237 6171
rect 2237 6137 2271 6171
rect 2271 6137 2280 6171
rect 2228 6128 2280 6137
rect 2688 6060 2740 6112
rect 7564 6196 7616 6248
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 8668 6196 8720 6205
rect 9956 6264 10008 6316
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 12164 6264 12216 6316
rect 12348 6264 12400 6316
rect 12532 6264 12584 6316
rect 12900 6264 12952 6316
rect 9220 6196 9272 6248
rect 9496 6196 9548 6248
rect 10140 6196 10192 6248
rect 10692 6196 10744 6248
rect 14004 6264 14056 6316
rect 14280 6307 14332 6316
rect 14280 6273 14289 6307
rect 14289 6273 14323 6307
rect 14323 6273 14332 6307
rect 14280 6264 14332 6273
rect 5172 6171 5224 6180
rect 5172 6137 5206 6171
rect 5206 6137 5224 6171
rect 5172 6128 5224 6137
rect 7932 6128 7984 6180
rect 8116 6128 8168 6180
rect 8760 6128 8812 6180
rect 9036 6128 9088 6180
rect 4712 6060 4764 6112
rect 5632 6060 5684 6112
rect 10600 6128 10652 6180
rect 15660 6196 15712 6248
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12440 6060 12492 6069
rect 12716 6060 12768 6112
rect 12900 6103 12952 6112
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 14004 6103 14056 6112
rect 14004 6069 14013 6103
rect 14013 6069 14047 6103
rect 14047 6069 14056 6103
rect 14004 6060 14056 6069
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 2412 5856 2464 5908
rect 8576 5856 8628 5908
rect 9312 5856 9364 5908
rect 2228 5788 2280 5840
rect 7012 5788 7064 5840
rect 7288 5788 7340 5840
rect 9404 5788 9456 5840
rect 2136 5763 2188 5772
rect 2136 5729 2145 5763
rect 2145 5729 2179 5763
rect 2179 5729 2188 5763
rect 2136 5720 2188 5729
rect 4160 5720 4212 5772
rect 5540 5720 5592 5772
rect 5724 5763 5776 5772
rect 5724 5729 5758 5763
rect 5758 5729 5776 5763
rect 5724 5720 5776 5729
rect 8116 5720 8168 5772
rect 8944 5720 8996 5772
rect 10600 5856 10652 5908
rect 11244 5856 11296 5908
rect 12716 5899 12768 5908
rect 12716 5865 12725 5899
rect 12725 5865 12759 5899
rect 12759 5865 12768 5899
rect 12716 5856 12768 5865
rect 12992 5856 13044 5908
rect 14188 5856 14240 5908
rect 10048 5788 10100 5840
rect 12440 5788 12492 5840
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 2780 5516 2832 5568
rect 4068 5652 4120 5704
rect 5172 5652 5224 5704
rect 6828 5652 6880 5704
rect 8760 5652 8812 5704
rect 9588 5720 9640 5772
rect 9772 5720 9824 5772
rect 10232 5720 10284 5772
rect 10784 5720 10836 5772
rect 11888 5763 11940 5772
rect 11888 5729 11897 5763
rect 11897 5729 11931 5763
rect 11931 5729 11940 5763
rect 11888 5720 11940 5729
rect 13636 5720 13688 5772
rect 14188 5720 14240 5772
rect 8576 5584 8628 5636
rect 8944 5584 8996 5636
rect 4068 5516 4120 5568
rect 4344 5516 4396 5568
rect 4620 5516 4672 5568
rect 5448 5516 5500 5568
rect 8668 5559 8720 5568
rect 8668 5525 8677 5559
rect 8677 5525 8711 5559
rect 8711 5525 8720 5559
rect 8668 5516 8720 5525
rect 9864 5516 9916 5568
rect 10048 5516 10100 5568
rect 10416 5516 10468 5568
rect 11152 5584 11204 5636
rect 11520 5559 11572 5568
rect 11520 5525 11529 5559
rect 11529 5525 11563 5559
rect 11563 5525 11572 5559
rect 11520 5516 11572 5525
rect 12808 5516 12860 5568
rect 13544 5652 13596 5704
rect 12992 5584 13044 5636
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 13912 5559 13964 5568
rect 13912 5525 13921 5559
rect 13921 5525 13955 5559
rect 13955 5525 13964 5559
rect 13912 5516 13964 5525
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 6828 5312 6880 5364
rect 7932 5312 7984 5364
rect 4160 5244 4212 5296
rect 4896 5244 4948 5296
rect 6368 5244 6420 5296
rect 6736 5244 6788 5296
rect 7840 5244 7892 5296
rect 8576 5244 8628 5296
rect 10692 5244 10744 5296
rect 11980 5312 12032 5364
rect 12164 5312 12216 5364
rect 12900 5312 12952 5364
rect 13084 5312 13136 5364
rect 2412 5108 2464 5160
rect 3148 5108 3200 5160
rect 3700 5108 3752 5160
rect 4896 5151 4948 5160
rect 4896 5117 4905 5151
rect 4905 5117 4939 5151
rect 4939 5117 4948 5151
rect 4896 5108 4948 5117
rect 9680 5176 9732 5228
rect 11152 5244 11204 5296
rect 14004 5312 14056 5364
rect 14372 5312 14424 5364
rect 14648 5312 14700 5364
rect 12808 5176 12860 5228
rect 13084 5176 13136 5228
rect 5448 5108 5500 5160
rect 5540 5108 5592 5160
rect 9404 5108 9456 5160
rect 9864 5108 9916 5160
rect 10416 5108 10468 5160
rect 11796 5108 11848 5160
rect 11980 5108 12032 5160
rect 14188 5108 14240 5160
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 2320 5015 2372 5024
rect 2320 4981 2329 5015
rect 2329 4981 2363 5015
rect 2363 4981 2372 5015
rect 2320 4972 2372 4981
rect 3332 4972 3384 5024
rect 6184 5040 6236 5092
rect 7104 5083 7156 5092
rect 7104 5049 7138 5083
rect 7138 5049 7156 5083
rect 7104 5040 7156 5049
rect 7840 5040 7892 5092
rect 8576 5040 8628 5092
rect 8760 5040 8812 5092
rect 9128 5040 9180 5092
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 6828 4972 6880 5024
rect 10600 5040 10652 5092
rect 10784 5040 10836 5092
rect 11888 5040 11940 5092
rect 12532 5040 12584 5092
rect 13452 5083 13504 5092
rect 9680 4972 9732 5024
rect 9956 4972 10008 5024
rect 10140 4972 10192 5024
rect 11612 4972 11664 5024
rect 12256 4972 12308 5024
rect 12716 4972 12768 5024
rect 13084 4972 13136 5024
rect 13452 5049 13461 5083
rect 13461 5049 13495 5083
rect 13495 5049 13504 5083
rect 13452 5040 13504 5049
rect 14648 5176 14700 5228
rect 15292 5176 15344 5228
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 3332 4768 3384 4820
rect 2228 4632 2280 4684
rect 2596 4700 2648 4752
rect 7564 4768 7616 4820
rect 11796 4768 11848 4820
rect 12348 4768 12400 4820
rect 12624 4768 12676 4820
rect 12808 4768 12860 4820
rect 13176 4768 13228 4820
rect 6828 4700 6880 4752
rect 3148 4632 3200 4684
rect 5080 4632 5132 4684
rect 5540 4675 5592 4684
rect 5540 4641 5574 4675
rect 5574 4641 5592 4675
rect 5540 4632 5592 4641
rect 5816 4632 5868 4684
rect 3516 4539 3568 4548
rect 3516 4505 3525 4539
rect 3525 4505 3559 4539
rect 3559 4505 3568 4539
rect 3516 4496 3568 4505
rect 3700 4496 3752 4548
rect 4344 4496 4396 4548
rect 4896 4564 4948 4616
rect 6736 4632 6788 4684
rect 7380 4675 7432 4684
rect 7380 4641 7414 4675
rect 7414 4641 7432 4675
rect 7380 4632 7432 4641
rect 8668 4700 8720 4752
rect 8760 4632 8812 4684
rect 9680 4632 9732 4684
rect 8944 4564 8996 4616
rect 9588 4564 9640 4616
rect 9956 4700 10008 4752
rect 10416 4700 10468 4752
rect 10876 4700 10928 4752
rect 11060 4700 11112 4752
rect 11152 4700 11204 4752
rect 10784 4632 10836 4684
rect 10416 4564 10468 4616
rect 11888 4700 11940 4752
rect 13360 4632 13412 4684
rect 11612 4564 11664 4616
rect 12716 4564 12768 4616
rect 2504 4428 2556 4480
rect 4160 4428 4212 4480
rect 6184 4428 6236 4480
rect 7380 4428 7432 4480
rect 8668 4496 8720 4548
rect 13084 4496 13136 4548
rect 14188 4564 14240 4616
rect 14648 4564 14700 4616
rect 9128 4428 9180 4480
rect 9864 4428 9916 4480
rect 10232 4428 10284 4480
rect 11152 4428 11204 4480
rect 14004 4428 14056 4480
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 3240 4224 3292 4276
rect 5632 4224 5684 4276
rect 8116 4224 8168 4276
rect 8944 4224 8996 4276
rect 9772 4224 9824 4276
rect 10324 4224 10376 4276
rect 2872 4156 2924 4208
rect 4712 4156 4764 4208
rect 7840 4156 7892 4208
rect 11796 4224 11848 4276
rect 12900 4224 12952 4276
rect 13912 4224 13964 4276
rect 14188 4224 14240 4276
rect 14372 4224 14424 4276
rect 388 4088 440 4140
rect 1584 4088 1636 4140
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 4896 4131 4948 4140
rect 756 4020 808 4072
rect 1400 4020 1452 4072
rect 3148 4020 3200 4072
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 4252 3952 4304 4004
rect 2228 3927 2280 3936
rect 2228 3893 2237 3927
rect 2237 3893 2271 3927
rect 2271 3893 2280 3927
rect 2228 3884 2280 3893
rect 6184 4020 6236 4072
rect 4988 3952 5040 4004
rect 5172 3995 5224 4004
rect 5172 3961 5206 3995
rect 5206 3961 5224 3995
rect 6736 4020 6788 4072
rect 8116 4088 8168 4140
rect 8668 4020 8720 4072
rect 10324 4088 10376 4140
rect 10416 4131 10468 4140
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 10876 4088 10928 4140
rect 12440 4156 12492 4208
rect 13176 4156 13228 4208
rect 13452 4156 13504 4208
rect 12348 4088 12400 4140
rect 12532 4088 12584 4140
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 14004 4088 14056 4140
rect 14464 4156 14516 4208
rect 15016 4199 15068 4208
rect 15016 4165 15025 4199
rect 15025 4165 15059 4199
rect 15059 4165 15068 4199
rect 15016 4156 15068 4165
rect 14372 4088 14424 4140
rect 15476 4088 15528 4140
rect 5172 3952 5224 3961
rect 5540 3884 5592 3936
rect 7472 3952 7524 4004
rect 7748 3952 7800 4004
rect 8116 3952 8168 4004
rect 10784 3952 10836 4004
rect 9312 3884 9364 3936
rect 10048 3884 10100 3936
rect 10416 3884 10468 3936
rect 10692 3884 10744 3936
rect 11796 4020 11848 4072
rect 11980 4020 12032 4072
rect 14648 4020 14700 4072
rect 11336 3952 11388 4004
rect 13268 3952 13320 4004
rect 11704 3884 11756 3936
rect 13820 3884 13872 3936
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 1676 3680 1728 3732
rect 1952 3723 2004 3732
rect 1952 3689 1961 3723
rect 1961 3689 1995 3723
rect 1995 3689 2004 3723
rect 1952 3680 2004 3689
rect 2596 3680 2648 3732
rect 3884 3680 3936 3732
rect 2872 3612 2924 3664
rect 3332 3612 3384 3664
rect 5724 3680 5776 3732
rect 1860 3544 1912 3596
rect 4160 3544 4212 3596
rect 6276 3612 6328 3664
rect 6828 3680 6880 3732
rect 8576 3680 8628 3732
rect 8944 3723 8996 3732
rect 8944 3689 8953 3723
rect 8953 3689 8987 3723
rect 8987 3689 8996 3723
rect 8944 3680 8996 3689
rect 9312 3680 9364 3732
rect 9680 3612 9732 3664
rect 1952 3476 2004 3528
rect 4160 3340 4212 3392
rect 4988 3408 5040 3460
rect 6736 3544 6788 3596
rect 7564 3587 7616 3596
rect 7564 3553 7573 3587
rect 7573 3553 7607 3587
rect 7607 3553 7616 3587
rect 7564 3544 7616 3553
rect 9772 3544 9824 3596
rect 10048 3680 10100 3732
rect 12348 3680 12400 3732
rect 13452 3680 13504 3732
rect 9956 3612 10008 3664
rect 10324 3544 10376 3596
rect 11428 3544 11480 3596
rect 5448 3476 5500 3528
rect 8576 3476 8628 3528
rect 11336 3519 11388 3528
rect 7104 3383 7156 3392
rect 7104 3349 7113 3383
rect 7113 3349 7147 3383
rect 7147 3349 7156 3383
rect 7104 3340 7156 3349
rect 8208 3340 8260 3392
rect 11336 3485 11345 3519
rect 11345 3485 11379 3519
rect 11379 3485 11388 3519
rect 11336 3476 11388 3485
rect 11704 3612 11756 3664
rect 11980 3612 12032 3664
rect 12900 3612 12952 3664
rect 13176 3612 13228 3664
rect 11888 3544 11940 3596
rect 11612 3476 11664 3528
rect 12440 3476 12492 3528
rect 13084 3476 13136 3528
rect 10416 3408 10468 3460
rect 13360 3408 13412 3460
rect 13820 3408 13872 3460
rect 14648 3451 14700 3460
rect 14648 3417 14657 3451
rect 14657 3417 14691 3451
rect 14691 3417 14700 3451
rect 14648 3408 14700 3417
rect 10600 3340 10652 3392
rect 12072 3383 12124 3392
rect 12072 3349 12081 3383
rect 12081 3349 12115 3383
rect 12115 3349 12124 3383
rect 12072 3340 12124 3349
rect 12624 3340 12676 3392
rect 12900 3340 12952 3392
rect 14096 3340 14148 3392
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 2320 3136 2372 3188
rect 4252 3136 4304 3188
rect 1952 3068 2004 3120
rect 3332 3000 3384 3052
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 1676 2932 1728 2984
rect 4068 2975 4120 2984
rect 4068 2941 4077 2975
rect 4077 2941 4111 2975
rect 4111 2941 4120 2975
rect 4068 2932 4120 2941
rect 5540 3136 5592 3188
rect 5632 3136 5684 3188
rect 5908 3068 5960 3120
rect 6552 3068 6604 3120
rect 7840 3068 7892 3120
rect 11520 3136 11572 3188
rect 11612 3136 11664 3188
rect 13176 3136 13228 3188
rect 13728 3136 13780 3188
rect 4896 2975 4948 2984
rect 4896 2941 4905 2975
rect 4905 2941 4939 2975
rect 4939 2941 4948 2975
rect 4896 2932 4948 2941
rect 6736 3000 6788 3052
rect 10324 3068 10376 3120
rect 14464 3068 14516 3120
rect 15016 3111 15068 3120
rect 15016 3077 15025 3111
rect 15025 3077 15059 3111
rect 15059 3077 15068 3111
rect 15016 3068 15068 3077
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 9956 3000 10008 3052
rect 6368 2932 6420 2984
rect 13728 3000 13780 3052
rect 14096 3043 14148 3052
rect 14096 3009 14105 3043
rect 14105 3009 14139 3043
rect 14139 3009 14148 3043
rect 14096 3000 14148 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 14556 3000 14608 3052
rect 1860 2907 1912 2916
rect 1860 2873 1869 2907
rect 1869 2873 1903 2907
rect 1903 2873 1912 2907
rect 1860 2864 1912 2873
rect 5080 2796 5132 2848
rect 5816 2864 5868 2916
rect 6460 2864 6512 2916
rect 6736 2864 6788 2916
rect 7196 2864 7248 2916
rect 7748 2864 7800 2916
rect 5540 2796 5592 2848
rect 8208 2796 8260 2848
rect 10048 2864 10100 2916
rect 11152 2932 11204 2984
rect 11520 2975 11572 2984
rect 11520 2941 11529 2975
rect 11529 2941 11563 2975
rect 11563 2941 11572 2975
rect 11520 2932 11572 2941
rect 11796 2932 11848 2984
rect 9036 2839 9088 2848
rect 9036 2805 9045 2839
rect 9045 2805 9079 2839
rect 9079 2805 9088 2839
rect 9036 2796 9088 2805
rect 10416 2796 10468 2848
rect 12532 2864 12584 2916
rect 13268 2864 13320 2916
rect 13452 2864 13504 2916
rect 11244 2796 11296 2848
rect 12440 2839 12492 2848
rect 12440 2805 12449 2839
rect 12449 2805 12483 2839
rect 12483 2805 12492 2839
rect 12440 2796 12492 2805
rect 12992 2796 13044 2848
rect 13176 2796 13228 2848
rect 13636 2796 13688 2848
rect 14464 2796 14516 2848
rect 14832 2796 14884 2848
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 2044 2456 2096 2508
rect 4988 2592 5040 2644
rect 5448 2592 5500 2644
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 7012 2592 7064 2644
rect 7564 2592 7616 2644
rect 4712 2524 4764 2576
rect 5540 2524 5592 2576
rect 2872 2456 2924 2508
rect 3976 2456 4028 2508
rect 10048 2592 10100 2644
rect 10232 2635 10284 2644
rect 10232 2601 10241 2635
rect 10241 2601 10275 2635
rect 10275 2601 10284 2635
rect 10232 2592 10284 2601
rect 11336 2635 11388 2644
rect 9588 2524 9640 2576
rect 10140 2567 10192 2576
rect 10140 2533 10149 2567
rect 10149 2533 10183 2567
rect 10183 2533 10192 2567
rect 10140 2524 10192 2533
rect 11336 2601 11345 2635
rect 11345 2601 11379 2635
rect 11379 2601 11388 2635
rect 11336 2592 11388 2601
rect 11428 2592 11480 2644
rect 12440 2592 12492 2644
rect 14188 2592 14240 2644
rect 12716 2524 12768 2576
rect 12992 2567 13044 2576
rect 12992 2533 13001 2567
rect 13001 2533 13035 2567
rect 13035 2533 13044 2567
rect 12992 2524 13044 2533
rect 8760 2456 8812 2508
rect 9496 2499 9548 2508
rect 9496 2465 9505 2499
rect 9505 2465 9539 2499
rect 9539 2465 9548 2499
rect 9496 2456 9548 2465
rect 10692 2456 10744 2508
rect 4344 2431 4396 2440
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 8116 2388 8168 2440
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 7380 2320 7432 2372
rect 9312 2388 9364 2440
rect 11796 2456 11848 2508
rect 12440 2456 12492 2508
rect 15200 2499 15252 2508
rect 15200 2465 15209 2499
rect 15209 2465 15243 2499
rect 15243 2465 15252 2499
rect 15200 2456 15252 2465
rect 112 2252 164 2304
rect 6736 2252 6788 2304
rect 8208 2252 8260 2304
rect 9864 2320 9916 2372
rect 12532 2388 12584 2440
rect 14556 2388 14608 2440
rect 11888 2320 11940 2372
rect 12808 2320 12860 2372
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 9772 2295 9824 2304
rect 9772 2261 9781 2295
rect 9781 2261 9815 2295
rect 9815 2261 9824 2295
rect 9772 2252 9824 2261
rect 10048 2252 10100 2304
rect 11336 2252 11388 2304
rect 12256 2252 12308 2304
rect 13820 2295 13872 2304
rect 13820 2261 13829 2295
rect 13829 2261 13863 2295
rect 13863 2261 13872 2295
rect 13820 2252 13872 2261
rect 13912 2252 13964 2304
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 4068 2048 4120 2100
rect 8852 2048 8904 2100
rect 9312 2048 9364 2100
rect 11796 2048 11848 2100
rect 13820 1980 13872 2032
rect 4344 1912 4396 1964
rect 16028 1912 16080 1964
rect 2044 1844 2096 1896
rect 8760 1844 8812 1896
rect 3516 1776 3568 1828
rect 6920 1776 6972 1828
rect 9588 1776 9640 1828
rect 13912 1776 13964 1828
rect 3056 1708 3108 1760
rect 9312 1708 9364 1760
rect 9772 1708 9824 1760
rect 14924 1708 14976 1760
rect 7564 1640 7616 1692
rect 11520 1640 11572 1692
rect 4988 1572 5040 1624
rect 11428 1572 11480 1624
rect 6920 1504 6972 1556
rect 13084 1504 13136 1556
rect 8116 1436 8168 1488
rect 1400 1232 1452 1284
rect 6828 1232 6880 1284
<< metal2 >>
rect 110 19520 166 20000
rect 386 19520 442 20000
rect 754 19520 810 20000
rect 1122 19520 1178 20000
rect 1398 19520 1454 20000
rect 1766 19520 1822 20000
rect 2134 19520 2190 20000
rect 2410 19520 2466 20000
rect 2778 19520 2834 20000
rect 3146 19520 3202 20000
rect 3514 19520 3570 20000
rect 3790 19520 3846 20000
rect 4158 19520 4214 20000
rect 4526 19520 4582 20000
rect 4802 19520 4858 20000
rect 5170 19520 5226 20000
rect 5538 19520 5594 20000
rect 5814 19520 5870 20000
rect 6182 19520 6238 20000
rect 6550 19520 6606 20000
rect 6918 19520 6974 20000
rect 7194 19520 7250 20000
rect 7562 19520 7618 20000
rect 7930 19520 7986 20000
rect 8206 19520 8262 20000
rect 8574 19520 8630 20000
rect 8942 19520 8998 20000
rect 9218 19520 9274 20000
rect 9586 19520 9642 20000
rect 9954 19520 10010 20000
rect 10322 19520 10378 20000
rect 10598 19520 10654 20000
rect 10966 19520 11022 20000
rect 11334 19520 11390 20000
rect 11610 19520 11666 20000
rect 11978 19520 12034 20000
rect 12346 19520 12402 20000
rect 12622 19520 12678 20000
rect 12990 19520 13046 20000
rect 13358 19520 13414 20000
rect 13726 19520 13782 20000
rect 14002 19520 14058 20000
rect 14370 19520 14426 20000
rect 14738 19520 14794 20000
rect 15014 19520 15070 20000
rect 15382 19520 15438 20000
rect 15750 19520 15806 20000
rect 16026 19520 16082 20000
rect 16394 19520 16450 20000
rect 16762 19520 16818 20000
rect 124 16046 152 19520
rect 112 16040 164 16046
rect 112 15982 164 15988
rect 400 15978 428 19520
rect 768 17202 796 19520
rect 756 17196 808 17202
rect 756 17138 808 17144
rect 1136 16250 1164 19520
rect 1124 16244 1176 16250
rect 1124 16186 1176 16192
rect 1412 16114 1440 19520
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 1504 17134 1532 19343
rect 1674 18456 1730 18465
rect 1674 18391 1730 18400
rect 1492 17128 1544 17134
rect 1492 17070 1544 17076
rect 1504 16522 1532 17070
rect 1688 16726 1716 18391
rect 1676 16720 1728 16726
rect 1676 16662 1728 16668
rect 1492 16516 1544 16522
rect 1492 16458 1544 16464
rect 1780 16114 1808 19520
rect 2148 17202 2176 19520
rect 2424 17270 2452 19520
rect 2412 17264 2464 17270
rect 2412 17206 2464 17212
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 388 15972 440 15978
rect 388 15914 440 15920
rect 1320 15638 1348 15982
rect 1308 15632 1360 15638
rect 1308 15574 1360 15580
rect 1492 15564 1544 15570
rect 1492 15506 1544 15512
rect 1308 15496 1360 15502
rect 1308 15438 1360 15444
rect 1320 11830 1348 15438
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1308 11824 1360 11830
rect 1308 11766 1360 11772
rect 1214 8392 1270 8401
rect 1214 8327 1216 8336
rect 1268 8327 1270 8336
rect 1216 8298 1268 8304
rect 1308 8288 1360 8294
rect 1308 8230 1360 8236
rect 1320 6866 1348 8230
rect 1308 6860 1360 6866
rect 1308 6802 1360 6808
rect 1412 6746 1440 13874
rect 1504 7290 1532 15506
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1596 11354 1624 13806
rect 1780 11898 1808 14894
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 1596 7426 1624 10950
rect 1688 7993 1716 11086
rect 1674 7984 1730 7993
rect 1674 7919 1730 7928
rect 1780 7546 1808 11630
rect 1872 10690 1900 14894
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 1964 11121 1992 11154
rect 1950 11112 2006 11121
rect 1950 11047 2006 11056
rect 1872 10662 1992 10690
rect 1860 10532 1912 10538
rect 1860 10474 1912 10480
rect 1872 10441 1900 10474
rect 1858 10432 1914 10441
rect 1858 10367 1914 10376
rect 1964 10282 1992 10662
rect 1872 10254 1992 10282
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1596 7398 1808 7426
rect 1504 7262 1716 7290
rect 1412 6718 1532 6746
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 388 4140 440 4146
rect 388 4082 440 4088
rect 112 2304 164 2310
rect 112 2246 164 2252
rect 124 480 152 2246
rect 400 480 428 4082
rect 1412 4078 1440 6598
rect 1504 5409 1532 6718
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1490 5400 1546 5409
rect 1490 5335 1546 5344
rect 1596 4146 1624 5510
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 756 4072 808 4078
rect 756 4014 808 4020
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 768 480 796 4014
rect 1688 3738 1716 7262
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1780 3618 1808 7398
rect 1872 7313 1900 10254
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1858 7304 1914 7313
rect 1858 7239 1914 7248
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1688 3590 1808 3618
rect 1872 3602 1900 4966
rect 1964 3738 1992 8774
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1860 3596 1912 3602
rect 1122 3088 1178 3097
rect 1122 3023 1178 3032
rect 1136 480 1164 3023
rect 1688 2990 1716 3590
rect 1860 3538 1912 3544
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1766 3360 1822 3369
rect 1766 3295 1822 3304
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1400 1284 1452 1290
rect 1400 1226 1452 1232
rect 1412 480 1440 1226
rect 1780 480 1808 3295
rect 1964 3126 1992 3470
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1858 2952 1914 2961
rect 1858 2887 1860 2896
rect 1912 2887 1914 2896
rect 1860 2858 1912 2864
rect 2056 2632 2084 15438
rect 2228 15428 2280 15434
rect 2228 15370 2280 15376
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2148 10713 2176 13262
rect 2134 10704 2190 10713
rect 2134 10639 2190 10648
rect 2240 8106 2268 15370
rect 2332 9586 2360 16390
rect 2424 13977 2452 17070
rect 2792 16794 2820 19520
rect 3160 17542 3188 19520
rect 3528 17882 3556 19520
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3421 17436 3717 17456
rect 3477 17434 3501 17436
rect 3557 17434 3581 17436
rect 3637 17434 3661 17436
rect 3499 17382 3501 17434
rect 3563 17382 3575 17434
rect 3637 17382 3639 17434
rect 3477 17380 3501 17382
rect 3557 17380 3581 17382
rect 3637 17380 3661 17382
rect 2962 17368 3018 17377
rect 3421 17360 3717 17380
rect 2962 17303 3018 17312
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2410 13968 2466 13977
rect 2410 13903 2466 13912
rect 2516 13002 2544 16186
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2608 13258 2636 15438
rect 2700 14600 2728 16594
rect 2792 16250 2820 16594
rect 2870 16416 2926 16425
rect 2870 16351 2926 16360
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2700 14572 2820 14600
rect 2792 14521 2820 14572
rect 2884 14550 2912 16351
rect 2976 15706 3004 17303
rect 3700 17128 3752 17134
rect 3804 17116 3832 19520
rect 4068 17944 4120 17950
rect 4068 17886 4120 17892
rect 4080 17270 4108 17886
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 3804 17088 4108 17116
rect 3700 17070 3752 17076
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2964 14884 3016 14890
rect 2964 14826 3016 14832
rect 2872 14544 2924 14550
rect 2778 14512 2834 14521
rect 2872 14486 2924 14492
rect 2778 14447 2834 14456
rect 2870 13832 2926 13841
rect 2870 13767 2926 13776
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2596 13252 2648 13258
rect 2596 13194 2648 13200
rect 2516 12974 2728 13002
rect 2412 12912 2464 12918
rect 2412 12854 2464 12860
rect 2502 12880 2558 12889
rect 2424 12345 2452 12854
rect 2502 12815 2504 12824
rect 2556 12815 2558 12824
rect 2504 12786 2556 12792
rect 2596 12776 2648 12782
rect 2594 12744 2596 12753
rect 2648 12744 2650 12753
rect 2594 12679 2650 12688
rect 2596 12368 2648 12374
rect 2410 12336 2466 12345
rect 2596 12310 2648 12316
rect 2410 12271 2466 12280
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2148 8078 2268 8106
rect 2148 7041 2176 8078
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2240 7546 2268 7822
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2332 7410 2360 8230
rect 2424 8129 2452 11154
rect 2516 10266 2544 11154
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2608 10169 2636 12310
rect 2700 11014 2728 12974
rect 2792 12442 2820 13262
rect 2884 13190 2912 13767
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11694 2912 12038
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2594 10160 2650 10169
rect 2594 10095 2650 10104
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2502 9616 2558 9625
rect 2608 9586 2636 9862
rect 2700 9654 2728 10610
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 10266 2820 10406
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2502 9551 2558 9560
rect 2596 9580 2648 9586
rect 2516 9450 2544 9551
rect 2596 9522 2648 9528
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2792 9178 2820 10066
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2884 9722 2912 9998
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2976 9518 3004 14826
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 3068 12986 3096 14282
rect 3160 13734 3188 17002
rect 3332 16992 3384 16998
rect 3330 16960 3332 16969
rect 3384 16960 3386 16969
rect 3330 16895 3386 16904
rect 3712 16590 3740 17070
rect 3884 16652 3936 16658
rect 3884 16594 3936 16600
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3252 15434 3280 15982
rect 3344 15570 3372 16526
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 3421 16348 3717 16368
rect 3477 16346 3501 16348
rect 3557 16346 3581 16348
rect 3637 16346 3661 16348
rect 3499 16294 3501 16346
rect 3563 16294 3575 16346
rect 3637 16294 3639 16346
rect 3477 16292 3501 16294
rect 3557 16292 3581 16294
rect 3637 16292 3661 16294
rect 3421 16272 3717 16292
rect 3424 16176 3476 16182
rect 3424 16118 3476 16124
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 3436 15348 3464 16118
rect 3608 15972 3660 15978
rect 3608 15914 3660 15920
rect 3620 15473 3648 15914
rect 3606 15464 3662 15473
rect 3606 15399 3662 15408
rect 3344 15320 3464 15348
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3068 12345 3096 12378
rect 3054 12336 3110 12345
rect 3054 12271 3110 12280
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 3068 11762 3096 12106
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2410 8120 2466 8129
rect 2410 8055 2466 8064
rect 2410 7984 2466 7993
rect 2410 7919 2466 7928
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2134 7032 2190 7041
rect 2134 6967 2190 6976
rect 2136 6792 2188 6798
rect 2332 6780 2360 7210
rect 2188 6752 2360 6780
rect 2136 6734 2188 6740
rect 2148 6254 2176 6734
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 2226 6216 2282 6225
rect 2148 5778 2176 6190
rect 2226 6151 2228 6160
rect 2280 6151 2282 6160
rect 2228 6122 2280 6128
rect 2240 5846 2268 6122
rect 2424 5914 2452 7919
rect 2516 7290 2544 8978
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2608 7750 2636 8230
rect 2700 8090 2728 9046
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2516 7262 2636 7290
rect 2700 7274 2728 7890
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 2516 6662 2544 7142
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2608 6361 2636 7262
rect 2688 7268 2740 7274
rect 2688 7210 2740 7216
rect 2792 7002 2820 8978
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2594 6352 2650 6361
rect 2594 6287 2650 6296
rect 2700 6118 2728 6938
rect 2884 6497 2912 9454
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2976 8401 3004 8434
rect 2962 8392 3018 8401
rect 2962 8327 3018 8336
rect 3068 7449 3096 11494
rect 3160 10810 3188 12242
rect 3252 11393 3280 14962
rect 3344 13870 3372 15320
rect 3421 15260 3717 15280
rect 3477 15258 3501 15260
rect 3557 15258 3581 15260
rect 3637 15258 3661 15260
rect 3499 15206 3501 15258
rect 3563 15206 3575 15258
rect 3637 15206 3639 15258
rect 3477 15204 3501 15206
rect 3557 15204 3581 15206
rect 3637 15204 3661 15206
rect 3421 15184 3717 15204
rect 3421 14172 3717 14192
rect 3477 14170 3501 14172
rect 3557 14170 3581 14172
rect 3637 14170 3661 14172
rect 3499 14118 3501 14170
rect 3563 14118 3575 14170
rect 3637 14118 3639 14170
rect 3477 14116 3501 14118
rect 3557 14116 3581 14118
rect 3637 14116 3661 14118
rect 3421 14096 3717 14116
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3332 13456 3384 13462
rect 3332 13398 3384 13404
rect 3344 11898 3372 13398
rect 3421 13084 3717 13104
rect 3477 13082 3501 13084
rect 3557 13082 3581 13084
rect 3637 13082 3661 13084
rect 3499 13030 3501 13082
rect 3563 13030 3575 13082
rect 3637 13030 3639 13082
rect 3477 13028 3501 13030
rect 3557 13028 3581 13030
rect 3637 13028 3661 13030
rect 3421 13008 3717 13028
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3528 12170 3556 12650
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3421 11996 3717 12016
rect 3477 11994 3501 11996
rect 3557 11994 3581 11996
rect 3637 11994 3661 11996
rect 3499 11942 3501 11994
rect 3563 11942 3575 11994
rect 3637 11942 3639 11994
rect 3477 11940 3501 11942
rect 3557 11940 3581 11942
rect 3637 11940 3661 11942
rect 3421 11920 3717 11940
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3238 11384 3294 11393
rect 3238 11319 3294 11328
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3054 7440 3110 7449
rect 3054 7375 3110 7384
rect 3160 7324 3188 10406
rect 3252 9636 3280 11086
rect 3344 10538 3372 11698
rect 3421 10908 3717 10928
rect 3477 10906 3501 10908
rect 3557 10906 3581 10908
rect 3637 10906 3661 10908
rect 3499 10854 3501 10906
rect 3563 10854 3575 10906
rect 3637 10854 3639 10906
rect 3477 10852 3501 10854
rect 3557 10852 3581 10854
rect 3637 10852 3661 10854
rect 3421 10832 3717 10852
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 3330 10432 3386 10441
rect 3330 10367 3386 10376
rect 3344 9704 3372 10367
rect 3804 10266 3832 16458
rect 3896 10470 3924 16594
rect 3988 14006 4016 16594
rect 4080 16114 4108 17088
rect 4172 16810 4200 19520
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4264 17202 4292 17478
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4172 16782 4384 16810
rect 4252 16652 4304 16658
rect 4172 16612 4252 16640
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4172 15450 4200 16612
rect 4252 16594 4304 16600
rect 4356 16522 4384 16782
rect 4436 16720 4488 16726
rect 4436 16662 4488 16668
rect 4344 16516 4396 16522
rect 4344 16458 4396 16464
rect 4448 16454 4476 16662
rect 4540 16658 4568 19520
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4436 16040 4488 16046
rect 4342 16008 4398 16017
rect 4252 15972 4304 15978
rect 4436 15982 4488 15988
rect 4342 15943 4398 15952
rect 4252 15914 4304 15920
rect 4080 15422 4200 15450
rect 4080 14385 4108 15422
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4172 15026 4200 15302
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4264 14618 4292 15914
rect 4356 15910 4384 15943
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4342 15056 4398 15065
rect 4342 14991 4398 15000
rect 4356 14890 4384 14991
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 4448 14618 4476 15982
rect 4620 15632 4672 15638
rect 4620 15574 4672 15580
rect 4632 15473 4660 15574
rect 4724 15570 4752 16526
rect 4816 16454 4844 19520
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4908 16130 4936 16730
rect 5000 16697 5028 16934
rect 4986 16688 5042 16697
rect 4986 16623 5042 16632
rect 5080 16584 5132 16590
rect 5080 16526 5132 16532
rect 4908 16102 5028 16130
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4618 15464 4674 15473
rect 4618 15399 4674 15408
rect 4724 15042 4752 15506
rect 4816 15162 4844 15982
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4632 15014 4844 15042
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4540 14414 4568 14962
rect 4632 14414 4660 15014
rect 4816 14958 4844 15014
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4712 14884 4764 14890
rect 4712 14826 4764 14832
rect 4528 14408 4580 14414
rect 4066 14376 4122 14385
rect 4528 14350 4580 14356
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4066 14311 4122 14320
rect 4252 14340 4304 14346
rect 4252 14282 4304 14288
rect 3976 14000 4028 14006
rect 3976 13942 4028 13948
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4080 13569 4108 13874
rect 4066 13560 4122 13569
rect 4066 13495 4122 13504
rect 4264 12322 4292 14282
rect 4540 13802 4568 14350
rect 4632 13870 4660 14350
rect 4724 14346 4752 14826
rect 4908 14618 4936 15982
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4712 14340 4764 14346
rect 4712 14282 4764 14288
rect 4816 14074 4844 14418
rect 4894 14376 4950 14385
rect 4894 14311 4950 14320
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4436 13796 4488 13802
rect 4436 13738 4488 13744
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4448 13530 4476 13738
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4356 13161 4384 13466
rect 4632 13410 4660 13806
rect 4448 13394 4660 13410
rect 4436 13388 4660 13394
rect 4488 13382 4660 13388
rect 4436 13330 4488 13336
rect 4342 13152 4398 13161
rect 4342 13087 4398 13096
rect 4632 12782 4660 13382
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4908 12481 4936 14311
rect 4894 12472 4950 12481
rect 4894 12407 4950 12416
rect 4080 12294 4292 12322
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4080 12238 4108 12294
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3421 9820 3717 9840
rect 3477 9818 3501 9820
rect 3557 9818 3581 9820
rect 3637 9818 3661 9820
rect 3499 9766 3501 9818
rect 3563 9766 3575 9818
rect 3637 9766 3639 9818
rect 3477 9764 3501 9766
rect 3557 9764 3581 9766
rect 3637 9764 3661 9766
rect 3421 9744 3717 9764
rect 3344 9676 3648 9704
rect 3252 9608 3464 9636
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3252 7970 3280 9454
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 9178 3372 9318
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3436 9058 3464 9608
rect 3620 9353 3648 9676
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3606 9344 3662 9353
rect 3606 9279 3662 9288
rect 3712 9217 3740 9590
rect 3804 9518 3832 9862
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3896 9450 3924 9998
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3988 9330 4016 11766
rect 4264 11762 4292 12294
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4434 12064 4490 12073
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4066 10840 4122 10849
rect 4066 10775 4122 10784
rect 4080 10606 4108 10775
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4264 10266 4292 11562
rect 4356 10266 4384 12038
rect 4434 11999 4490 12008
rect 4448 11150 4476 11999
rect 4526 11792 4582 11801
rect 4526 11727 4582 11736
rect 4540 11354 4568 11727
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4448 10674 4476 11086
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4448 10441 4476 10610
rect 4434 10432 4490 10441
rect 4434 10367 4490 10376
rect 4434 10296 4490 10305
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4344 10260 4396 10266
rect 4434 10231 4490 10240
rect 4344 10202 4396 10208
rect 3896 9302 4016 9330
rect 3698 9208 3754 9217
rect 3698 9143 3754 9152
rect 3344 9030 3464 9058
rect 3698 9072 3754 9081
rect 3344 8362 3372 9030
rect 3698 9007 3700 9016
rect 3752 9007 3754 9016
rect 3700 8978 3752 8984
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3421 8732 3717 8752
rect 3477 8730 3501 8732
rect 3557 8730 3581 8732
rect 3637 8730 3661 8732
rect 3499 8678 3501 8730
rect 3563 8678 3575 8730
rect 3637 8678 3639 8730
rect 3477 8676 3501 8678
rect 3557 8676 3581 8678
rect 3637 8676 3661 8678
rect 3421 8656 3717 8676
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3528 7993 3556 8434
rect 3804 8430 3832 8842
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3514 7984 3570 7993
rect 3252 7942 3372 7970
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3068 7296 3188 7324
rect 2962 7032 3018 7041
rect 2962 6967 3018 6976
rect 2870 6488 2926 6497
rect 2870 6423 2926 6432
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2228 5840 2280 5846
rect 2228 5782 2280 5788
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2424 5386 2452 5850
rect 2700 5658 2728 6054
rect 2700 5630 2820 5658
rect 2792 5574 2820 5630
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2240 5358 2452 5386
rect 2240 4690 2268 5358
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 2134 4584 2190 4593
rect 2134 4519 2190 4528
rect 1964 2604 2084 2632
rect 1964 1465 1992 2604
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 2056 1902 2084 2450
rect 2044 1896 2096 1902
rect 2044 1838 2096 1844
rect 1950 1456 2006 1465
rect 1950 1391 2006 1400
rect 2148 480 2176 4519
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 3777 2268 3878
rect 2226 3768 2282 3777
rect 2226 3703 2282 3712
rect 2332 3194 2360 4966
rect 2424 4146 2452 5102
rect 2596 4752 2648 4758
rect 2596 4694 2648 4700
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2516 3618 2544 4422
rect 2608 3738 2636 4694
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2778 4040 2834 4049
rect 2778 3975 2834 3984
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2424 3590 2544 3618
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2424 480 2452 3590
rect 2792 480 2820 3975
rect 2884 3670 2912 4150
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2976 3505 3004 6967
rect 2962 3496 3018 3505
rect 2962 3431 3018 3440
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2884 513 2912 2450
rect 3068 1766 3096 7296
rect 3252 6458 3280 7822
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3344 5794 3372 7942
rect 3514 7919 3570 7928
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3421 7644 3717 7664
rect 3477 7642 3501 7644
rect 3557 7642 3581 7644
rect 3637 7642 3661 7644
rect 3499 7590 3501 7642
rect 3563 7590 3575 7642
rect 3637 7590 3639 7642
rect 3477 7588 3501 7590
rect 3557 7588 3581 7590
rect 3637 7588 3661 7590
rect 3421 7568 3717 7588
rect 3804 7002 3832 7822
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 3790 6216 3846 6225
rect 3790 6151 3846 6160
rect 3252 5766 3372 5794
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3160 4690 3188 5102
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3160 4078 3188 4626
rect 3252 4457 3280 5766
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 3700 5160 3752 5166
rect 3514 5128 3570 5137
rect 3700 5102 3752 5108
rect 3514 5063 3570 5072
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3344 4826 3372 4966
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3528 4554 3556 5063
rect 3712 4554 3740 5102
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3238 4448 3294 4457
rect 3238 4383 3294 4392
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3252 3346 3280 4218
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 3160 3318 3280 3346
rect 3056 1760 3108 1766
rect 3056 1702 3108 1708
rect 2870 504 2926 513
rect 110 0 166 480
rect 386 0 442 480
rect 754 0 810 480
rect 1122 0 1178 480
rect 1398 0 1454 480
rect 1766 0 1822 480
rect 2134 0 2190 480
rect 2410 0 2466 480
rect 2778 0 2834 480
rect 3160 480 3188 3318
rect 3344 3058 3372 3606
rect 3421 3292 3717 3312
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3421 2128 3717 2148
rect 3516 1828 3568 1834
rect 3516 1770 3568 1776
rect 3528 480 3556 1770
rect 3804 480 3832 6151
rect 3896 3738 3924 9302
rect 3974 8528 4030 8537
rect 3974 8463 4030 8472
rect 3988 8362 4016 8463
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3988 7721 4016 7754
rect 3974 7712 4030 7721
rect 3974 7647 4030 7656
rect 3976 6792 4028 6798
rect 4080 6780 4108 10202
rect 4250 9344 4306 9353
rect 4250 9279 4306 9288
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4172 6866 4200 7414
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4028 6752 4108 6780
rect 3976 6734 4028 6740
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3988 2514 4016 6734
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4068 5704 4120 5710
rect 4066 5672 4068 5681
rect 4120 5672 4122 5681
rect 4066 5607 4122 5616
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 2990 4108 5510
rect 4172 5302 4200 5714
rect 4160 5296 4212 5302
rect 4264 5273 4292 9279
rect 4448 9042 4476 10231
rect 4540 10198 4568 11018
rect 4632 10538 4660 12242
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4632 10062 4660 10474
rect 4724 10305 4752 12310
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4908 12073 4936 12174
rect 4894 12064 4950 12073
rect 4894 11999 4950 12008
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4908 10674 4936 11630
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4710 10296 4766 10305
rect 4710 10231 4766 10240
rect 4908 10062 4936 10610
rect 4620 10056 4672 10062
rect 4896 10056 4948 10062
rect 4620 9998 4672 10004
rect 4710 10024 4766 10033
rect 4528 9988 4580 9994
rect 4896 9998 4948 10004
rect 4710 9959 4766 9968
rect 4528 9930 4580 9936
rect 4540 9761 4568 9930
rect 4526 9752 4582 9761
rect 4526 9687 4582 9696
rect 4724 9568 4752 9959
rect 4908 9926 4936 9998
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 5000 9586 5028 16102
rect 4632 9540 4752 9568
rect 4988 9580 5040 9586
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4540 9353 4568 9454
rect 4526 9344 4582 9353
rect 4526 9279 4582 9288
rect 4632 9194 4660 9540
rect 4988 9522 5040 9528
rect 4804 9512 4856 9518
rect 4540 9166 4660 9194
rect 4724 9472 4804 9500
rect 4436 9036 4488 9042
rect 4356 8996 4436 9024
rect 4356 5574 4384 8996
rect 4436 8978 4488 8984
rect 4540 8922 4568 9166
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 4448 8906 4568 8922
rect 4436 8900 4568 8906
rect 4488 8894 4568 8900
rect 4436 8842 4488 8848
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4434 7032 4490 7041
rect 4434 6967 4490 6976
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4160 5238 4212 5244
rect 4250 5264 4306 5273
rect 4250 5199 4306 5208
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4160 4480 4212 4486
rect 4356 4457 4384 4490
rect 4160 4422 4212 4428
rect 4342 4448 4398 4457
rect 4172 3602 4200 4422
rect 4342 4383 4398 4392
rect 4252 4004 4304 4010
rect 4304 3964 4384 3992
rect 4252 3946 4304 3952
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4250 3360 4306 3369
rect 4172 3058 4200 3334
rect 4250 3295 4306 3304
rect 4264 3194 4292 3295
rect 4356 3233 4384 3964
rect 4342 3224 4398 3233
rect 4252 3188 4304 3194
rect 4342 3159 4398 3168
rect 4252 3130 4304 3136
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4068 2984 4120 2990
rect 4448 2938 4476 6967
rect 4540 5896 4568 8774
rect 4632 8537 4660 9046
rect 4618 8528 4674 8537
rect 4618 8463 4674 8472
rect 4724 8430 4752 9472
rect 4804 9454 4856 9460
rect 4986 9480 5042 9489
rect 4986 9415 5042 9424
rect 5000 9382 5028 9415
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5092 9194 5120 16526
rect 5184 15994 5212 19520
rect 5552 17746 5580 19520
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5448 17604 5500 17610
rect 5448 17546 5500 17552
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5184 15966 5304 15994
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5184 13530 5212 15642
rect 5276 15366 5304 15966
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5184 12782 5212 13466
rect 5276 13462 5304 14758
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 5184 10810 5212 11562
rect 5276 11150 5304 12650
rect 5368 11665 5396 16730
rect 5460 16658 5488 17546
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5644 16114 5672 16934
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5446 15600 5502 15609
rect 5446 15535 5502 15544
rect 5460 15502 5488 15535
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5552 14550 5580 16050
rect 5736 15994 5764 16934
rect 5828 16561 5856 19520
rect 6196 17270 6224 19520
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 5886 16892 6182 16912
rect 5942 16890 5966 16892
rect 6022 16890 6046 16892
rect 6102 16890 6126 16892
rect 5964 16838 5966 16890
rect 6028 16838 6040 16890
rect 6102 16838 6104 16890
rect 5942 16836 5966 16838
rect 6022 16836 6046 16838
rect 6102 16836 6126 16838
rect 5886 16816 6182 16836
rect 6288 16794 6316 17002
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6092 16584 6144 16590
rect 5814 16552 5870 16561
rect 6092 16526 6144 16532
rect 5814 16487 5870 16496
rect 6104 16114 6132 16526
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6104 15994 6132 16050
rect 5644 15966 5764 15994
rect 5828 15966 6132 15994
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 12102 5488 13738
rect 5552 13462 5580 14350
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5552 12306 5580 12650
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5354 11656 5410 11665
rect 5354 11591 5410 11600
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5184 9722 5212 10746
rect 5354 10568 5410 10577
rect 5354 10503 5410 10512
rect 5262 9752 5318 9761
rect 5172 9716 5224 9722
rect 5262 9687 5264 9696
rect 5172 9658 5224 9664
rect 5316 9687 5318 9696
rect 5264 9658 5316 9664
rect 4908 9166 5120 9194
rect 5170 9208 5226 9217
rect 4802 8936 4858 8945
rect 4802 8871 4804 8880
rect 4856 8871 4858 8880
rect 4804 8842 4856 8848
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4618 7984 4674 7993
rect 4618 7919 4674 7928
rect 4632 6497 4660 7919
rect 4724 7342 4752 8366
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4724 6798 4752 7278
rect 4816 7177 4844 8434
rect 4908 7478 4936 9166
rect 5170 9143 5226 9152
rect 5184 9110 5212 9143
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4986 7440 5042 7449
rect 4986 7375 5042 7384
rect 4802 7168 4858 7177
rect 4802 7103 4858 7112
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4618 6488 4674 6497
rect 4618 6423 4620 6432
rect 4672 6423 4674 6432
rect 4620 6394 4672 6400
rect 4632 6363 4660 6394
rect 4724 6322 4752 6734
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4724 6118 4752 6258
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4908 5930 4936 6870
rect 4816 5902 4936 5930
rect 4540 5868 4752 5896
rect 4526 5808 4582 5817
rect 4526 5743 4582 5752
rect 4068 2926 4120 2932
rect 4172 2910 4476 2938
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4066 2408 4122 2417
rect 4066 2343 4122 2352
rect 4080 2106 4108 2343
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 4172 480 4200 2910
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4356 1970 4384 2382
rect 4344 1964 4396 1970
rect 4344 1906 4396 1912
rect 4540 480 4568 5743
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4632 3505 4660 5510
rect 4724 4729 4752 5868
rect 4710 4720 4766 4729
rect 4710 4655 4766 4664
rect 4724 4214 4752 4655
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4618 3496 4674 3505
rect 4618 3431 4674 3440
rect 4724 2582 4752 4150
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4816 480 4844 5902
rect 5000 5386 5028 7375
rect 5092 6866 5120 8978
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5184 8090 5212 8366
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5368 6934 5396 10503
rect 5460 9761 5488 11086
rect 5552 10810 5580 12106
rect 5644 11257 5672 15966
rect 5724 15428 5776 15434
rect 5724 15370 5776 15376
rect 5736 14929 5764 15370
rect 5828 15144 5856 15966
rect 5886 15804 6182 15824
rect 5942 15802 5966 15804
rect 6022 15802 6046 15804
rect 6102 15802 6126 15804
rect 5964 15750 5966 15802
rect 6028 15750 6040 15802
rect 6102 15750 6104 15802
rect 5942 15748 5966 15750
rect 6022 15748 6046 15750
rect 6102 15748 6126 15750
rect 5886 15728 6182 15748
rect 6564 15609 6592 19520
rect 6932 17678 6960 19520
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 7208 17542 7236 19520
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7576 17338 7604 19520
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7300 16590 7328 17138
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6550 15600 6606 15609
rect 6550 15535 6606 15544
rect 6550 15464 6606 15473
rect 6550 15399 6606 15408
rect 5908 15156 5960 15162
rect 5828 15116 5908 15144
rect 5722 14920 5778 14929
rect 5722 14855 5778 14864
rect 5722 13560 5778 13569
rect 5722 13495 5724 13504
rect 5776 13495 5778 13504
rect 5724 13466 5776 13472
rect 5736 12374 5764 13466
rect 5828 13394 5856 15116
rect 5908 15098 5960 15104
rect 5886 14716 6182 14736
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6126 14716
rect 5964 14662 5966 14714
rect 6028 14662 6040 14714
rect 6102 14662 6104 14714
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6126 14662
rect 5886 14640 6182 14660
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 6288 14006 6316 14486
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 5886 13628 6182 13648
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6126 13628
rect 5964 13574 5966 13626
rect 6028 13574 6040 13626
rect 6102 13574 6104 13626
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6126 13574
rect 5886 13552 6182 13572
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 6288 12986 6316 13398
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6182 12744 6238 12753
rect 6182 12679 6238 12688
rect 6196 12628 6224 12679
rect 6196 12600 6316 12628
rect 6288 12594 6316 12600
rect 6458 12608 6514 12617
rect 6288 12566 6458 12594
rect 5886 12540 6182 12560
rect 6458 12543 6514 12552
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6126 12540
rect 5964 12486 5966 12538
rect 6028 12486 6040 12538
rect 6102 12486 6104 12538
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6126 12486
rect 5886 12464 6182 12484
rect 6564 12374 6592 15399
rect 6656 12442 6684 16186
rect 7012 16176 7064 16182
rect 7012 16118 7064 16124
rect 6736 15904 6788 15910
rect 6788 15852 6960 15858
rect 6736 15846 6960 15852
rect 6748 15830 6960 15846
rect 6932 15638 6960 15830
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6920 15632 6972 15638
rect 6920 15574 6972 15580
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6748 13870 6776 14962
rect 6840 14550 6868 15574
rect 6920 14884 6972 14890
rect 7024 14872 7052 16118
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 6972 14844 7052 14872
rect 6920 14826 6972 14832
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6748 13394 6776 13806
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6840 12918 6868 13330
rect 6932 13025 6960 14826
rect 7300 14793 7328 15982
rect 7392 15706 7420 16050
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7286 14784 7342 14793
rect 7286 14719 7342 14728
rect 7484 14618 7512 17138
rect 7656 16992 7708 16998
rect 7654 16960 7656 16969
rect 7708 16960 7710 16969
rect 7654 16895 7710 16904
rect 7852 16794 7880 17750
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7748 16584 7800 16590
rect 7944 16572 7972 19520
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 8128 16726 8156 16934
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8116 16584 8168 16590
rect 7944 16544 8116 16572
rect 7748 16526 7800 16532
rect 8116 16526 8168 16532
rect 7760 15366 7788 16526
rect 8114 16144 8170 16153
rect 8220 16130 8248 19520
rect 8588 17626 8616 19520
rect 8956 17950 8984 19520
rect 8944 17944 8996 17950
rect 8944 17886 8996 17892
rect 8942 17640 8998 17649
rect 8588 17598 8800 17626
rect 8352 17436 8648 17456
rect 8408 17434 8432 17436
rect 8488 17434 8512 17436
rect 8568 17434 8592 17436
rect 8430 17382 8432 17434
rect 8494 17382 8506 17434
rect 8568 17382 8570 17434
rect 8408 17380 8432 17382
rect 8488 17380 8512 17382
rect 8568 17380 8592 17382
rect 8352 17360 8648 17380
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8588 16833 8616 16934
rect 8574 16824 8630 16833
rect 8574 16759 8630 16768
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8352 16348 8648 16368
rect 8408 16346 8432 16348
rect 8488 16346 8512 16348
rect 8568 16346 8592 16348
rect 8430 16294 8432 16346
rect 8494 16294 8506 16346
rect 8568 16294 8570 16346
rect 8408 16292 8432 16294
rect 8488 16292 8512 16294
rect 8568 16292 8592 16294
rect 8352 16272 8648 16292
rect 8220 16102 8340 16130
rect 8114 16079 8170 16088
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7392 13802 7420 14350
rect 7484 13870 7512 14554
rect 7576 14482 7604 14554
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7668 13734 7696 15302
rect 7760 14482 7788 15302
rect 7852 15094 7880 15846
rect 8128 15706 8156 16079
rect 8116 15700 8168 15706
rect 8116 15642 8168 15648
rect 8312 15638 8340 16102
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8128 15473 8156 15506
rect 8114 15464 8170 15473
rect 8114 15399 8170 15408
rect 8352 15260 8648 15280
rect 8408 15258 8432 15260
rect 8488 15258 8512 15260
rect 8568 15258 8592 15260
rect 8430 15206 8432 15258
rect 8494 15206 8506 15258
rect 8568 15206 8570 15258
rect 8408 15204 8432 15206
rect 8488 15204 8512 15206
rect 8568 15204 8592 15206
rect 8352 15184 8648 15204
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7760 13988 7788 14418
rect 7840 14000 7892 14006
rect 7760 13960 7840 13988
rect 7840 13942 7892 13948
rect 7944 13938 7972 14758
rect 8128 14482 8156 15098
rect 8680 14657 8708 16594
rect 8772 16250 8800 17598
rect 8942 17575 8998 17584
rect 8956 16794 8984 17575
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8666 14648 8722 14657
rect 8666 14583 8722 14592
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8128 14074 8156 14214
rect 8352 14172 8648 14192
rect 8408 14170 8432 14172
rect 8488 14170 8512 14172
rect 8568 14170 8592 14172
rect 8430 14118 8432 14170
rect 8494 14118 8506 14170
rect 8568 14118 8570 14170
rect 8408 14116 8432 14118
rect 8488 14116 8512 14118
rect 8568 14116 8592 14118
rect 8352 14096 8648 14116
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7746 13696 7802 13705
rect 7746 13631 7802 13640
rect 7102 13560 7158 13569
rect 7102 13495 7158 13504
rect 7010 13152 7066 13161
rect 7010 13087 7066 13096
rect 6918 13016 6974 13025
rect 6918 12951 6974 12960
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6920 12776 6972 12782
rect 6734 12744 6790 12753
rect 6920 12718 6972 12724
rect 6734 12679 6790 12688
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 5814 12200 5870 12209
rect 5814 12135 5870 12144
rect 5724 11688 5776 11694
rect 5828 11676 5856 12135
rect 5776 11648 5856 11676
rect 5724 11630 5776 11636
rect 5630 11248 5686 11257
rect 5828 11218 5856 11648
rect 5886 11452 6182 11472
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6126 11452
rect 5964 11398 5966 11450
rect 6028 11398 6040 11450
rect 6102 11398 6104 11450
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6126 11398
rect 5886 11376 6182 11396
rect 6550 11384 6606 11393
rect 6550 11319 6606 11328
rect 5630 11183 5632 11192
rect 5684 11183 5686 11192
rect 5816 11212 5868 11218
rect 5632 11154 5684 11160
rect 5816 11154 5868 11160
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 6368 10464 6420 10470
rect 5722 10432 5778 10441
rect 6368 10406 6420 10412
rect 5722 10367 5778 10376
rect 5736 10130 5764 10367
rect 5886 10364 6182 10384
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6126 10364
rect 5964 10310 5966 10362
rect 6028 10310 6040 10362
rect 6102 10310 6104 10362
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6126 10310
rect 5886 10288 6182 10308
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 6380 10033 6408 10406
rect 6366 10024 6422 10033
rect 6366 9959 6422 9968
rect 5630 9888 5686 9897
rect 5630 9823 5686 9832
rect 5446 9752 5502 9761
rect 5446 9687 5502 9696
rect 5644 9450 5672 9823
rect 5816 9512 5868 9518
rect 5814 9480 5816 9489
rect 5868 9480 5870 9489
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5724 9444 5776 9450
rect 5814 9415 5870 9424
rect 6276 9444 6328 9450
rect 5724 9386 5776 9392
rect 6276 9386 6328 9392
rect 5736 9353 5764 9386
rect 5722 9344 5778 9353
rect 5722 9279 5778 9288
rect 5886 9276 6182 9296
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6126 9276
rect 5964 9222 5966 9274
rect 6028 9222 6040 9274
rect 6102 9222 6104 9274
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6126 9222
rect 5886 9200 6182 9220
rect 6288 8566 6316 9386
rect 6458 8800 6514 8809
rect 6458 8735 6514 8744
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 5886 8188 6182 8208
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6126 8188
rect 5964 8134 5966 8186
rect 6028 8134 6040 8186
rect 6102 8134 6104 8186
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6126 8134
rect 5886 8112 6182 8132
rect 6380 8129 6408 8298
rect 6366 8120 6422 8129
rect 6366 8055 6422 8064
rect 5722 7984 5778 7993
rect 5632 7948 5684 7954
rect 5722 7919 5778 7928
rect 6000 7948 6052 7954
rect 5632 7890 5684 7896
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5354 6760 5410 6769
rect 5354 6695 5410 6704
rect 5264 6656 5316 6662
rect 5170 6624 5226 6633
rect 5264 6598 5316 6604
rect 5170 6559 5226 6568
rect 5184 6458 5212 6559
rect 5276 6458 5304 6598
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5184 6186 5212 6394
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 4908 5358 5028 5386
rect 4908 5302 4936 5358
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4908 4622 4936 5102
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4908 4146 4936 4558
rect 5092 4185 5120 4626
rect 5078 4176 5134 4185
rect 4896 4140 4948 4146
rect 5078 4111 5134 4120
rect 4896 4082 4948 4088
rect 4908 2990 4936 4082
rect 5184 4010 5212 5646
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5000 3466 5028 3946
rect 5078 3496 5134 3505
rect 4988 3460 5040 3466
rect 5078 3431 5134 3440
rect 4988 3402 5040 3408
rect 4896 2984 4948 2990
rect 4948 2944 5028 2972
rect 4896 2926 4948 2932
rect 5000 2650 5028 2944
rect 5092 2854 5120 3431
rect 5368 3380 5396 6695
rect 5460 6633 5488 7686
rect 5538 7576 5594 7585
rect 5538 7511 5594 7520
rect 5552 6730 5580 7511
rect 5644 7206 5672 7890
rect 5736 7342 5764 7919
rect 6000 7890 6052 7896
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5920 7342 5948 7822
rect 6012 7546 6040 7890
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 6288 7206 6316 7346
rect 5632 7200 5684 7206
rect 5724 7200 5776 7206
rect 5632 7142 5684 7148
rect 5722 7168 5724 7177
rect 6276 7200 6328 7206
rect 5776 7168 5778 7177
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5446 6624 5502 6633
rect 5446 6559 5502 6568
rect 5644 6118 5672 7142
rect 6276 7142 6328 7148
rect 6366 7168 6422 7177
rect 5722 7103 5778 7112
rect 5886 7100 6182 7120
rect 6366 7103 6422 7112
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6126 7100
rect 5964 7046 5966 7098
rect 6028 7046 6040 7098
rect 6102 7046 6104 7098
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6126 7046
rect 5886 7024 6182 7044
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6288 6390 6316 6938
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 6380 5896 6408 7103
rect 6196 5868 6408 5896
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5460 5166 5488 5510
rect 5552 5166 5580 5714
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5736 4672 5764 5714
rect 6196 5098 6224 5868
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 5816 4684 5868 4690
rect 5736 4644 5816 4672
rect 5552 3942 5580 4626
rect 5630 4312 5686 4321
rect 5630 4247 5632 4256
rect 5684 4247 5686 4256
rect 5632 4218 5684 4224
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5184 3352 5396 3380
rect 5080 2848 5132 2854
rect 5078 2816 5080 2825
rect 5132 2816 5134 2825
rect 5078 2751 5134 2760
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5000 2446 5028 2586
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5000 1630 5028 2382
rect 4988 1624 5040 1630
rect 4988 1566 5040 1572
rect 5184 480 5212 3352
rect 5460 2650 5488 3470
rect 5552 3194 5580 3878
rect 5630 3768 5686 3777
rect 5736 3738 5764 4644
rect 5816 4626 5868 4632
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6196 4078 6224 4422
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 5886 3836 6182 3856
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 5630 3703 5686 3712
rect 5724 3732 5776 3738
rect 5644 3194 5672 3703
rect 5724 3674 5776 3680
rect 6288 3670 6316 4966
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 6380 3482 6408 5238
rect 6288 3454 6408 3482
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5908 3120 5960 3126
rect 5644 3068 5908 3074
rect 5644 3062 5960 3068
rect 5644 3046 5948 3062
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5552 2582 5580 2790
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 5644 1442 5672 3046
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 5552 1414 5672 1442
rect 5552 480 5580 1414
rect 5828 480 5856 2858
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 6288 1170 6316 3454
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6380 2650 6408 2926
rect 6472 2922 6500 8735
rect 6564 3126 6592 11319
rect 6748 11014 6776 12679
rect 6932 12442 6960 12718
rect 7024 12481 7052 13087
rect 7010 12472 7066 12481
rect 6920 12436 6972 12442
rect 7010 12407 7066 12416
rect 6920 12378 6972 12384
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 11218 6960 11494
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 7024 10538 7052 12407
rect 7116 10849 7144 13495
rect 7472 13456 7524 13462
rect 7472 13398 7524 13404
rect 7484 13190 7512 13398
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 7392 12238 7420 12650
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7392 11762 7420 12174
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7392 11150 7420 11698
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7102 10840 7158 10849
rect 7102 10775 7158 10784
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 7024 10441 7052 10474
rect 7010 10432 7066 10441
rect 7010 10367 7066 10376
rect 6642 10160 6698 10169
rect 7208 10130 7236 10950
rect 7286 10704 7342 10713
rect 7286 10639 7288 10648
rect 7340 10639 7342 10648
rect 7288 10610 7340 10616
rect 7392 10538 7420 11086
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 6642 10095 6698 10104
rect 7196 10124 7248 10130
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6656 2972 6684 10095
rect 7196 10066 7248 10072
rect 7288 10124 7340 10130
rect 7392 10112 7420 10474
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7340 10084 7420 10112
rect 7288 10066 7340 10072
rect 6828 10056 6880 10062
rect 6734 10024 6790 10033
rect 7484 10010 7512 10134
rect 6828 9998 6880 10004
rect 6734 9959 6790 9968
rect 6748 5302 6776 9959
rect 6840 9586 6868 9998
rect 7392 9982 7512 10010
rect 7194 9752 7250 9761
rect 7194 9687 7250 9696
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 7208 9450 7236 9687
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7392 9382 7420 9982
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6840 7342 6868 8366
rect 7024 8362 7052 8910
rect 7392 8838 7420 9318
rect 7576 9178 7604 12582
rect 7668 11694 7696 13126
rect 7760 12374 7788 13631
rect 8036 13530 8064 14010
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 7838 13016 7894 13025
rect 7838 12951 7894 12960
rect 7852 12850 7880 12951
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 8128 12782 8156 13738
rect 8680 13734 8708 13806
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8312 13394 8340 13466
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8312 13240 8340 13330
rect 8404 13297 8432 13330
rect 8220 13212 8340 13240
rect 8390 13288 8446 13297
rect 8390 13223 8446 13232
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8220 12714 8248 13212
rect 8352 13084 8648 13104
rect 8408 13082 8432 13084
rect 8488 13082 8512 13084
rect 8568 13082 8592 13084
rect 8430 13030 8432 13082
rect 8494 13030 8506 13082
rect 8568 13030 8570 13082
rect 8408 13028 8432 13030
rect 8488 13028 8512 13030
rect 8568 13028 8592 13030
rect 8352 13008 8648 13028
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 8496 12424 8524 12854
rect 8680 12850 8708 13670
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8496 12396 8708 12424
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 8390 12200 8446 12209
rect 8390 12135 8392 12144
rect 8444 12135 8446 12144
rect 8392 12106 8444 12112
rect 8352 11996 8648 12016
rect 8408 11994 8432 11996
rect 8488 11994 8512 11996
rect 8568 11994 8592 11996
rect 8430 11942 8432 11994
rect 8494 11942 8506 11994
rect 8568 11942 8570 11994
rect 8408 11940 8432 11942
rect 8488 11940 8512 11942
rect 8568 11940 8592 11942
rect 8352 11920 8648 11940
rect 8680 11898 8708 12396
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 8680 11626 8708 11698
rect 8668 11620 8720 11626
rect 8668 11562 8720 11568
rect 8666 11520 8722 11529
rect 8666 11455 8722 11464
rect 7748 11212 7800 11218
rect 7800 11172 7972 11200
rect 7748 11154 7800 11160
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10198 7696 10950
rect 7944 10674 7972 11172
rect 8352 10908 8648 10928
rect 8408 10906 8432 10908
rect 8488 10906 8512 10908
rect 8568 10906 8592 10908
rect 8430 10854 8432 10906
rect 8494 10854 8506 10906
rect 8568 10854 8570 10906
rect 8408 10852 8432 10854
rect 8488 10852 8512 10854
rect 8568 10852 8592 10854
rect 8352 10832 8648 10852
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 8024 9920 8076 9926
rect 8022 9888 8024 9897
rect 8076 9888 8078 9897
rect 8022 9823 8078 9832
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 7654 9208 7710 9217
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7564 9172 7616 9178
rect 7654 9143 7710 9152
rect 8024 9172 8076 9178
rect 7564 9114 7616 9120
rect 7484 8838 7512 9114
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7208 7546 7236 7686
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6840 7206 6868 7278
rect 7484 7206 7512 7686
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 6840 6322 6868 7142
rect 7484 6866 7512 7142
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6840 5710 6868 6258
rect 7576 6254 7604 7142
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 6918 6080 6974 6089
rect 6918 6015 6974 6024
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6840 5030 6868 5306
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6748 4078 6776 4626
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6748 3602 6776 4014
rect 6840 3738 6868 4694
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6748 3058 6776 3538
rect 6826 3360 6882 3369
rect 6826 3295 6882 3304
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6564 2944 6684 2972
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6196 1142 6316 1170
rect 6196 480 6224 1142
rect 6564 480 6592 2944
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6748 2310 6776 2858
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6840 1290 6868 3295
rect 6932 1834 6960 6015
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7024 2650 7052 5782
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7116 3398 7144 5034
rect 7300 4321 7328 5782
rect 7562 5672 7618 5681
rect 7562 5607 7618 5616
rect 7470 4992 7526 5001
rect 7470 4927 7526 4936
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7392 4486 7420 4626
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7286 4312 7342 4321
rect 7286 4247 7342 4256
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 6920 1828 6972 1834
rect 6920 1770 6972 1776
rect 6920 1556 6972 1562
rect 6920 1498 6972 1504
rect 6828 1284 6880 1290
rect 6828 1226 6880 1232
rect 6932 480 6960 1498
rect 7208 480 7236 2858
rect 7392 2378 7420 4422
rect 7484 4010 7512 4927
rect 7576 4826 7604 5607
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7484 2446 7512 3946
rect 7562 3768 7618 3777
rect 7562 3703 7618 3712
rect 7576 3602 7604 3703
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7668 3505 7696 9143
rect 8024 9114 8076 9120
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 6746 7788 8910
rect 7852 8566 7880 8978
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7944 8362 7972 8434
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7852 7954 7880 8230
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7944 7478 7972 8298
rect 8036 8090 8064 9114
rect 8128 9042 8156 9522
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8128 7698 8156 8978
rect 8220 8566 8248 10542
rect 8352 9820 8648 9840
rect 8408 9818 8432 9820
rect 8488 9818 8512 9820
rect 8568 9818 8592 9820
rect 8430 9766 8432 9818
rect 8494 9766 8506 9818
rect 8568 9766 8570 9818
rect 8408 9764 8432 9766
rect 8488 9764 8512 9766
rect 8568 9764 8592 9766
rect 8352 9744 8648 9764
rect 8482 9480 8538 9489
rect 8392 9444 8444 9450
rect 8482 9415 8538 9424
rect 8392 9386 8444 9392
rect 8404 8974 8432 9386
rect 8496 9042 8524 9415
rect 8680 9217 8708 11455
rect 8772 11354 8800 15914
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8758 9888 8814 9897
rect 8758 9823 8814 9832
rect 8772 9586 8800 9823
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8666 9208 8722 9217
rect 8666 9143 8722 9152
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8352 8732 8648 8752
rect 8408 8730 8432 8732
rect 8488 8730 8512 8732
rect 8568 8730 8592 8732
rect 8430 8678 8432 8730
rect 8494 8678 8506 8730
rect 8568 8678 8570 8730
rect 8408 8676 8432 8678
rect 8488 8676 8512 8678
rect 8568 8676 8592 8678
rect 8352 8656 8648 8676
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8772 8362 8800 9046
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8300 8288 8352 8294
rect 8220 8248 8300 8276
rect 8220 7721 8248 8248
rect 8300 8230 8352 8236
rect 8668 7744 8720 7750
rect 8036 7670 8156 7698
rect 8206 7712 8262 7721
rect 7932 7472 7984 7478
rect 7932 7414 7984 7420
rect 7838 6896 7894 6905
rect 7838 6831 7840 6840
rect 7892 6831 7894 6840
rect 7840 6802 7892 6808
rect 7760 6718 7880 6746
rect 7746 5400 7802 5409
rect 7746 5335 7802 5344
rect 7760 4010 7788 5335
rect 7852 5302 7880 6718
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7944 6390 7972 6598
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 7944 5370 7972 6122
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7852 4214 7880 5034
rect 7840 4208 7892 4214
rect 7840 4150 7892 4156
rect 7930 4176 7986 4185
rect 7930 4111 7986 4120
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 7654 3496 7710 3505
rect 7654 3431 7710 3440
rect 7760 2922 7788 3946
rect 7838 3224 7894 3233
rect 7838 3159 7894 3168
rect 7852 3126 7880 3159
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7562 2816 7618 2825
rect 7562 2751 7618 2760
rect 7576 2650 7604 2751
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7852 2553 7880 3062
rect 7562 2544 7618 2553
rect 7562 2479 7618 2488
rect 7838 2544 7894 2553
rect 7838 2479 7894 2488
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 7576 1698 7604 2479
rect 7564 1692 7616 1698
rect 7564 1634 7616 1640
rect 7576 480 7604 1634
rect 7944 480 7972 4111
rect 8036 3913 8064 7670
rect 8668 7686 8720 7692
rect 8206 7647 8262 7656
rect 8352 7644 8648 7664
rect 8408 7642 8432 7644
rect 8488 7642 8512 7644
rect 8568 7642 8592 7644
rect 8430 7590 8432 7642
rect 8494 7590 8506 7642
rect 8568 7590 8570 7642
rect 8408 7588 8432 7590
rect 8488 7588 8512 7590
rect 8568 7588 8592 7590
rect 8114 7576 8170 7585
rect 8352 7568 8648 7588
rect 8114 7511 8170 7520
rect 8128 7410 8156 7511
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8680 7342 8708 7686
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8404 7002 8432 7210
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8208 6656 8260 6662
rect 8206 6624 8208 6633
rect 8260 6624 8262 6633
rect 8206 6559 8262 6568
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8114 6488 8170 6497
rect 8352 6480 8648 6500
rect 8114 6423 8170 6432
rect 8128 6186 8156 6423
rect 8680 6254 8708 7278
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8116 6180 8168 6186
rect 8116 6122 8168 6128
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8116 5772 8168 5778
rect 8168 5732 8248 5760
rect 8116 5714 8168 5720
rect 8114 4448 8170 4457
rect 8114 4383 8170 4392
rect 8128 4282 8156 4383
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8128 4010 8156 4082
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8022 3904 8078 3913
rect 8022 3839 8078 3848
rect 8036 2825 8064 3839
rect 8220 3398 8248 5732
rect 8588 5642 8616 5850
rect 8772 5710 8800 6122
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8352 5392 8648 5412
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 8588 5098 8616 5238
rect 8576 5092 8628 5098
rect 8576 5034 8628 5040
rect 8680 5001 8708 5510
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8666 4992 8722 5001
rect 8666 4927 8722 4936
rect 8680 4758 8708 4927
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8772 4690 8800 5034
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8352 4380 8648 4400
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 8680 4078 8708 4490
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8772 3924 8800 4626
rect 8680 3896 8800 3924
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8588 3534 8616 3674
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8220 2854 8248 3334
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8352 3216 8648 3236
rect 8208 2848 8260 2854
rect 8022 2816 8078 2825
rect 8208 2790 8260 2796
rect 8574 2816 8630 2825
rect 8022 2751 8078 2760
rect 8574 2751 8630 2760
rect 8588 2446 8616 2751
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8128 1494 8156 2382
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8116 1488 8168 1494
rect 8116 1430 8168 1436
rect 8220 480 8248 2246
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 8680 2088 8708 3896
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8588 2060 8708 2088
rect 8588 480 8616 2060
rect 8772 1902 8800 2450
rect 8864 2106 8892 16594
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9048 16425 9076 16526
rect 9034 16416 9090 16425
rect 9034 16351 9090 16360
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 8956 15162 8984 15846
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8942 15056 8998 15065
rect 8942 14991 8998 15000
rect 8956 14414 8984 14991
rect 9048 14618 9076 15846
rect 9140 15570 9168 17002
rect 9232 15706 9260 19520
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9508 17354 9536 17818
rect 9600 17513 9628 19520
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9586 17504 9642 17513
rect 9586 17439 9642 17448
rect 9508 17326 9628 17354
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 9140 15065 9168 15506
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9126 15056 9182 15065
rect 9232 15026 9260 15438
rect 9126 14991 9182 15000
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9126 14784 9182 14793
rect 9126 14719 9182 14728
rect 9140 14618 9168 14719
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8956 13326 8984 14214
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8956 12986 8984 13262
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8942 12880 8998 12889
rect 8942 12815 8998 12824
rect 8956 12617 8984 12815
rect 8942 12608 8998 12617
rect 8942 12543 8998 12552
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8956 11830 8984 12038
rect 8944 11824 8996 11830
rect 8944 11766 8996 11772
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8956 11218 8984 11494
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8956 9586 8984 11154
rect 9048 11150 9076 14418
rect 9232 14346 9260 14962
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9140 11234 9168 14214
rect 9218 14104 9274 14113
rect 9218 14039 9274 14048
rect 9232 13190 9260 14039
rect 9324 13734 9352 16934
rect 9416 16522 9444 16934
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9416 15745 9444 16050
rect 9402 15736 9458 15745
rect 9402 15671 9458 15680
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9416 15162 9444 15302
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9324 13190 9352 13670
rect 9416 13530 9444 14962
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9312 12980 9364 12986
rect 9232 12940 9312 12968
rect 9232 12782 9260 12940
rect 9312 12922 9364 12928
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 11354 9260 11494
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9140 11206 9260 11234
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 10538 9076 10950
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 9034 10432 9090 10441
rect 9034 10367 9090 10376
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 9048 9466 9076 10367
rect 9140 9654 9168 11086
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9048 9438 9168 9466
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 8673 9076 9318
rect 9034 8664 9090 8673
rect 9034 8599 9090 8608
rect 8944 8560 8996 8566
rect 8944 8502 8996 8508
rect 9034 8528 9090 8537
rect 8956 5778 8984 8502
rect 9140 8514 9168 9438
rect 9090 8486 9168 8514
rect 9034 8463 9090 8472
rect 9048 8294 9076 8463
rect 9036 8288 9088 8294
rect 9128 8288 9180 8294
rect 9036 8230 9088 8236
rect 9126 8256 9128 8265
rect 9180 8256 9182 8265
rect 9126 8191 9182 8200
rect 9034 8120 9090 8129
rect 9034 8055 9090 8064
rect 9048 7750 9076 8055
rect 9232 7818 9260 11206
rect 9324 11150 9352 12718
rect 9416 12306 9444 13330
rect 9508 12442 9536 17070
rect 9600 16794 9628 17326
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9588 16448 9640 16454
rect 9692 16436 9720 17002
rect 9640 16408 9720 16436
rect 9588 16390 9640 16396
rect 9586 16280 9642 16289
rect 9586 16215 9642 16224
rect 9600 16046 9628 16215
rect 9784 16096 9812 18022
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9876 16425 9904 16526
rect 9862 16416 9918 16425
rect 9862 16351 9918 16360
rect 9968 16250 9996 19520
rect 10138 17368 10194 17377
rect 10138 17303 10194 17312
rect 10152 17202 10180 17303
rect 10232 17264 10284 17270
rect 10232 17206 10284 17212
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9692 16068 9812 16096
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9692 15570 9720 16068
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9784 15722 9812 15914
rect 9784 15694 9904 15722
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 15337 9720 15506
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9678 15328 9734 15337
rect 9678 15263 9734 15272
rect 9678 15056 9734 15065
rect 9678 14991 9734 15000
rect 9692 14890 9720 14991
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9600 14482 9628 14758
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9600 13161 9628 14418
rect 9692 13462 9720 14826
rect 9784 14793 9812 15438
rect 9876 14822 9904 15694
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 9864 14816 9916 14822
rect 9770 14784 9826 14793
rect 9864 14758 9916 14764
rect 9770 14719 9826 14728
rect 9770 14648 9826 14657
rect 9770 14583 9826 14592
rect 9784 14482 9812 14583
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9876 14278 9904 14350
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 9586 13152 9642 13161
rect 9586 13087 9642 13096
rect 9600 12986 9720 13002
rect 9600 12980 9732 12986
rect 9600 12974 9680 12980
rect 9600 12646 9628 12974
rect 9680 12922 9732 12928
rect 9784 12866 9812 13466
rect 9692 12838 9812 12866
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9588 12368 9640 12374
rect 9586 12336 9588 12345
rect 9640 12336 9642 12345
rect 9404 12300 9456 12306
rect 9586 12271 9642 12280
rect 9404 12242 9456 12248
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9416 10810 9444 12242
rect 9692 12186 9720 12838
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9508 12158 9720 12186
rect 9508 12102 9536 12158
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9586 11928 9642 11937
rect 9586 11863 9642 11872
rect 9600 11626 9628 11863
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9600 11286 9628 11562
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9494 10296 9550 10305
rect 9494 10231 9550 10240
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9036 6180 9088 6186
rect 9036 6122 9088 6128
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8944 5636 8996 5642
rect 8944 5578 8996 5584
rect 8956 4622 8984 5578
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8956 3738 8984 4218
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 8956 3369 8984 3674
rect 8942 3360 8998 3369
rect 8942 3295 8998 3304
rect 9048 2854 9076 6122
rect 9140 5098 9168 6802
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 4185 9168 4422
rect 9126 4176 9182 4185
rect 9126 4111 9182 4120
rect 9232 3040 9260 6190
rect 9324 5914 9352 10066
rect 9508 9926 9536 10231
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9416 9738 9444 9862
rect 9600 9738 9628 11018
rect 9416 9710 9628 9738
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9416 8090 9444 9522
rect 9494 9344 9550 9353
rect 9494 9279 9550 9288
rect 9508 8294 9536 9279
rect 9600 8809 9628 9710
rect 9692 9518 9720 12038
rect 9784 11082 9812 12650
rect 9876 12322 9904 13806
rect 9968 13734 9996 15370
rect 10060 14482 10088 17070
rect 10244 16998 10272 17206
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10336 16538 10364 19520
rect 10508 18012 10560 18018
rect 10508 17954 10560 17960
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10152 16510 10364 16538
rect 10152 15065 10180 16510
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10138 15056 10194 15065
rect 10138 14991 10194 15000
rect 10138 14920 10194 14929
rect 10138 14855 10194 14864
rect 10152 14618 10180 14855
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9968 13394 9996 13670
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 9968 12646 9996 12854
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9876 12294 9996 12322
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9876 12102 9904 12174
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9876 11257 9904 11494
rect 9862 11248 9918 11257
rect 9862 11183 9918 11192
rect 9968 11082 9996 12294
rect 10060 12102 10088 14418
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10152 14074 10180 14350
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10244 13870 10272 16390
rect 10336 16046 10364 16390
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10322 15328 10378 15337
rect 10322 15263 10378 15272
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10152 12238 10180 13738
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10244 12374 10272 12854
rect 10232 12368 10284 12374
rect 10232 12310 10284 12316
rect 10140 12232 10192 12238
rect 10138 12200 10140 12209
rect 10232 12232 10284 12238
rect 10192 12200 10194 12209
rect 10232 12174 10284 12180
rect 10138 12135 10194 12144
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10046 11520 10102 11529
rect 10046 11455 10102 11464
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9968 10713 9996 11018
rect 9954 10704 10010 10713
rect 9954 10639 10010 10648
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9784 9926 9812 10406
rect 9862 10296 9918 10305
rect 9862 10231 9918 10240
rect 9876 10198 9904 10231
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9770 9752 9826 9761
rect 9770 9687 9826 9696
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9784 9450 9812 9687
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9770 9344 9826 9353
rect 9692 8956 9720 9318
rect 9770 9279 9826 9288
rect 9784 9110 9812 9279
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9692 8928 9812 8956
rect 9784 8838 9812 8928
rect 9680 8832 9732 8838
rect 9586 8800 9642 8809
rect 9680 8774 9732 8780
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9586 8735 9642 8744
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9600 8090 9628 8570
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9416 7993 9444 8026
rect 9402 7984 9458 7993
rect 9402 7919 9458 7928
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9508 7002 9536 7822
rect 9586 7576 9642 7585
rect 9586 7511 9642 7520
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9402 6488 9458 6497
rect 9402 6423 9458 6432
rect 9416 6225 9444 6423
rect 9496 6248 9548 6254
rect 9402 6216 9458 6225
rect 9496 6190 9548 6196
rect 9402 6151 9458 6160
rect 9508 6066 9536 6190
rect 9416 6038 9536 6066
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9324 5692 9352 5850
rect 9416 5846 9444 6038
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 9600 5778 9628 7511
rect 9692 7274 9720 8774
rect 9876 8634 9904 9998
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9784 6905 9812 8434
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9876 8090 9904 8230
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9876 7478 9904 7686
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9770 6896 9826 6905
rect 9770 6831 9826 6840
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9324 5664 9536 5692
rect 9310 5536 9366 5545
rect 9310 5471 9366 5480
rect 9324 3942 9352 5471
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9416 5001 9444 5102
rect 9402 4992 9458 5001
rect 9402 4927 9458 4936
rect 9402 4720 9458 4729
rect 9402 4655 9458 4664
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 3738 9352 3878
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9312 3052 9364 3058
rect 9232 3012 9312 3040
rect 9312 2994 9364 3000
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9218 2816 9274 2825
rect 9218 2751 9274 2760
rect 8942 2680 8998 2689
rect 8942 2615 8998 2624
rect 8852 2100 8904 2106
rect 8852 2042 8904 2048
rect 8760 1896 8812 1902
rect 8760 1838 8812 1844
rect 8956 480 8984 2615
rect 9232 480 9260 2751
rect 9324 2446 9352 2994
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9324 2106 9352 2246
rect 9312 2100 9364 2106
rect 9312 2042 9364 2048
rect 9324 1766 9352 2042
rect 9312 1760 9364 1766
rect 9312 1702 9364 1708
rect 9416 1442 9444 4655
rect 9508 2514 9536 5664
rect 9692 5234 9720 6598
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9784 6089 9812 6326
rect 9968 6322 9996 10406
rect 10060 9432 10088 11455
rect 10152 11354 10180 12038
rect 10244 11694 10272 12174
rect 10336 12152 10364 15263
rect 10428 14521 10456 17070
rect 10520 16833 10548 17954
rect 10612 16969 10640 19520
rect 10690 17368 10746 17377
rect 10690 17303 10746 17312
rect 10598 16960 10654 16969
rect 10598 16895 10654 16904
rect 10506 16824 10562 16833
rect 10506 16759 10562 16768
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10520 16425 10548 16594
rect 10506 16416 10562 16425
rect 10506 16351 10562 16360
rect 10508 16176 10560 16182
rect 10508 16118 10560 16124
rect 10520 15570 10548 16118
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10520 15337 10548 15506
rect 10612 15450 10640 16895
rect 10704 15570 10732 17303
rect 10980 17241 11008 19520
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 10966 17232 11022 17241
rect 10966 17167 11022 17176
rect 10817 16892 11113 16912
rect 10873 16890 10897 16892
rect 10953 16890 10977 16892
rect 11033 16890 11057 16892
rect 10895 16838 10897 16890
rect 10959 16838 10971 16890
rect 11033 16838 11035 16890
rect 10873 16836 10897 16838
rect 10953 16836 10977 16838
rect 11033 16836 11057 16838
rect 10817 16816 11113 16836
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10796 16250 10824 16526
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10980 16182 11008 16594
rect 11256 16522 11284 17682
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11244 16516 11296 16522
rect 11244 16458 11296 16464
rect 11164 16402 11192 16458
rect 11164 16374 11284 16402
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 10817 15804 11113 15824
rect 10873 15802 10897 15804
rect 10953 15802 10977 15804
rect 11033 15802 11057 15804
rect 10895 15750 10897 15802
rect 10959 15750 10971 15802
rect 11033 15750 11035 15802
rect 10873 15748 10897 15750
rect 10953 15748 10977 15750
rect 11033 15748 11057 15750
rect 10817 15728 11113 15748
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10612 15422 10824 15450
rect 10600 15360 10652 15366
rect 10506 15328 10562 15337
rect 10600 15302 10652 15308
rect 10506 15263 10562 15272
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 10520 15026 10548 15098
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10414 14512 10470 14521
rect 10414 14447 10470 14456
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10428 13802 10456 14350
rect 10520 14249 10548 14758
rect 10506 14240 10562 14249
rect 10506 14175 10562 14184
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 10508 13796 10560 13802
rect 10508 13738 10560 13744
rect 10414 13696 10470 13705
rect 10414 13631 10470 13640
rect 10428 13394 10456 13631
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 10520 12900 10548 13738
rect 10416 12872 10548 12900
rect 10416 12696 10444 12872
rect 10416 12668 10456 12696
rect 10428 12481 10456 12668
rect 10414 12472 10470 12481
rect 10414 12407 10470 12416
rect 10336 12124 10456 12152
rect 10322 12064 10378 12073
rect 10322 11999 10378 12008
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10152 10130 10180 10610
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10244 9654 10272 11494
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10060 9404 10180 9432
rect 10152 9217 10180 9404
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10138 9208 10194 9217
rect 10138 9143 10194 9152
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10060 8498 10088 8910
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10060 7449 10088 7754
rect 10046 7440 10102 7449
rect 10046 7375 10102 7384
rect 10046 7168 10102 7177
rect 10046 7103 10102 7112
rect 10060 7002 10088 7103
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6633 10088 6734
rect 10152 6662 10180 9046
rect 10244 8956 10272 9318
rect 10336 9178 10364 11999
rect 10428 10826 10456 12124
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10520 11082 10548 11630
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10428 10798 10548 10826
rect 10414 10704 10470 10713
rect 10520 10674 10548 10798
rect 10612 10674 10640 15302
rect 10690 15056 10746 15065
rect 10690 14991 10746 15000
rect 10704 13802 10732 14991
rect 10796 14890 10824 15422
rect 10888 15065 10916 15506
rect 10874 15056 10930 15065
rect 10874 14991 10930 15000
rect 11164 14929 11192 15846
rect 11150 14920 11206 14929
rect 10784 14884 10836 14890
rect 11150 14855 11206 14864
rect 10784 14826 10836 14832
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 10817 14716 11113 14736
rect 10873 14714 10897 14716
rect 10953 14714 10977 14716
rect 11033 14714 11057 14716
rect 10895 14662 10897 14714
rect 10959 14662 10971 14714
rect 11033 14662 11035 14714
rect 10873 14660 10897 14662
rect 10953 14660 10977 14662
rect 11033 14660 11057 14662
rect 10817 14640 11113 14660
rect 11164 14600 11192 14758
rect 11072 14572 11192 14600
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10796 14346 10824 14486
rect 11072 14414 11100 14572
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10784 14340 10836 14346
rect 10784 14282 10836 14288
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10817 13628 11113 13648
rect 10873 13626 10897 13628
rect 10953 13626 10977 13628
rect 11033 13626 11057 13628
rect 10895 13574 10897 13626
rect 10959 13574 10971 13626
rect 11033 13574 11035 13626
rect 10873 13572 10897 13574
rect 10953 13572 10977 13574
rect 11033 13572 11057 13574
rect 10817 13552 11113 13572
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11072 12968 11100 13398
rect 11164 13161 11192 14418
rect 11256 13297 11284 16374
rect 11348 15026 11376 19520
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 11348 14521 11376 14962
rect 11440 14958 11468 16526
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11428 14952 11480 14958
rect 11428 14894 11480 14900
rect 11440 14657 11468 14894
rect 11426 14648 11482 14657
rect 11426 14583 11482 14592
rect 11334 14512 11390 14521
rect 11334 14447 11390 14456
rect 11428 14408 11480 14414
rect 11334 14376 11390 14385
rect 11428 14350 11480 14356
rect 11334 14311 11336 14320
rect 11388 14311 11390 14320
rect 11336 14282 11388 14288
rect 11440 13734 11468 14350
rect 11428 13728 11480 13734
rect 11428 13670 11480 13676
rect 11336 13320 11388 13326
rect 11242 13288 11298 13297
rect 11336 13262 11388 13268
rect 11242 13223 11298 13232
rect 11150 13152 11206 13161
rect 11150 13087 11206 13096
rect 11072 12940 11284 12968
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10704 11801 10732 12786
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 10817 12540 11113 12560
rect 10873 12538 10897 12540
rect 10953 12538 10977 12540
rect 11033 12538 11057 12540
rect 10895 12486 10897 12538
rect 10959 12486 10971 12538
rect 11033 12486 11035 12538
rect 10873 12484 10897 12486
rect 10953 12484 10977 12486
rect 11033 12484 11057 12486
rect 10817 12464 11113 12484
rect 11164 12442 11192 12718
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10968 12368 11020 12374
rect 11256 12356 11284 12940
rect 11348 12714 11376 13262
rect 11428 12912 11480 12918
rect 11428 12854 11480 12860
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11336 12368 11388 12374
rect 11256 12328 11336 12356
rect 10968 12310 11020 12316
rect 11336 12310 11388 12316
rect 10690 11792 10746 11801
rect 10888 11762 10916 12310
rect 10690 11727 10746 11736
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10980 11540 11008 12310
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 11072 11898 11100 12242
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 11440 11830 11468 12854
rect 11428 11824 11480 11830
rect 11150 11792 11206 11801
rect 11334 11792 11390 11801
rect 11150 11727 11206 11736
rect 11244 11756 11296 11762
rect 10704 11512 11008 11540
rect 10704 11218 10732 11512
rect 10817 11452 11113 11472
rect 10873 11450 10897 11452
rect 10953 11450 10977 11452
rect 11033 11450 11057 11452
rect 10895 11398 10897 11450
rect 10959 11398 10971 11450
rect 11033 11398 11035 11450
rect 10873 11396 10897 11398
rect 10953 11396 10977 11398
rect 11033 11396 11057 11398
rect 10817 11376 11113 11396
rect 11164 11336 11192 11727
rect 11428 11766 11480 11772
rect 11334 11727 11390 11736
rect 11244 11698 11296 11704
rect 10796 11308 11192 11336
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10704 10742 10732 11154
rect 10796 11014 10824 11308
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10968 11076 11020 11082
rect 10888 11036 10968 11064
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10414 10639 10470 10648
rect 10508 10668 10560 10674
rect 10428 10538 10456 10639
rect 10508 10610 10560 10616
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10888 10554 10916 11036
rect 10968 11018 11020 11024
rect 11072 10810 11100 11154
rect 11150 10976 11206 10985
rect 11150 10911 11206 10920
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10416 10532 10468 10538
rect 10704 10526 10916 10554
rect 10704 10520 10732 10526
rect 10468 10492 10548 10520
rect 10416 10474 10468 10480
rect 10414 10296 10470 10305
rect 10414 10231 10470 10240
rect 10428 10130 10456 10231
rect 10520 10130 10548 10492
rect 10612 10492 10732 10520
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10428 9586 10456 9930
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10520 9489 10548 9522
rect 10506 9480 10562 9489
rect 10506 9415 10562 9424
rect 10508 9376 10560 9382
rect 10506 9344 10508 9353
rect 10560 9344 10562 9353
rect 10506 9279 10562 9288
rect 10324 9172 10376 9178
rect 10376 9132 10548 9160
rect 10324 9114 10376 9120
rect 10336 9049 10364 9114
rect 10244 8928 10456 8956
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10244 7721 10272 8230
rect 10230 7712 10286 7721
rect 10230 7647 10286 7656
rect 10336 7562 10364 8570
rect 10428 7993 10456 8928
rect 10414 7984 10470 7993
rect 10414 7919 10470 7928
rect 10244 7534 10364 7562
rect 10140 6656 10192 6662
rect 10046 6624 10102 6633
rect 10140 6598 10192 6604
rect 10046 6559 10102 6568
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9770 6080 9826 6089
rect 9770 6015 9826 6024
rect 10060 5846 10088 6394
rect 10152 6254 10180 6394
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10138 5808 10194 5817
rect 9772 5772 9824 5778
rect 10244 5778 10272 7534
rect 10322 7440 10378 7449
rect 10322 7375 10378 7384
rect 10336 7041 10364 7375
rect 10322 7032 10378 7041
rect 10322 6967 10378 6976
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10138 5743 10194 5752
rect 10232 5772 10284 5778
rect 9772 5714 9824 5720
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9784 5137 9812 5714
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9876 5166 9904 5510
rect 9864 5160 9916 5166
rect 9770 5128 9826 5137
rect 9864 5102 9916 5108
rect 9770 5063 9826 5072
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9692 4690 9720 4966
rect 9968 4758 9996 4966
rect 9956 4752 10008 4758
rect 9956 4694 10008 4700
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9588 4616 9640 4622
rect 9640 4564 9720 4570
rect 9588 4558 9720 4564
rect 9600 4542 9720 4558
rect 9692 4536 9720 4542
rect 9692 4508 9812 4536
rect 9586 4448 9642 4457
rect 9586 4383 9642 4392
rect 9600 2689 9628 4383
rect 9784 4282 9812 4508
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9876 3890 9904 4422
rect 9954 4176 10010 4185
rect 9954 4111 10010 4120
rect 9692 3862 9904 3890
rect 9692 3670 9720 3862
rect 9770 3768 9826 3777
rect 9770 3703 9826 3712
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9784 3602 9812 3703
rect 9968 3670 9996 4111
rect 10060 3942 10088 5510
rect 10152 5114 10180 5743
rect 10232 5714 10284 5720
rect 10152 5086 10272 5114
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9968 3058 9996 3606
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 10060 2922 10088 3674
rect 10048 2916 10100 2922
rect 10048 2858 10100 2864
rect 9954 2816 10010 2825
rect 9954 2751 10010 2760
rect 9586 2680 9642 2689
rect 9586 2615 9642 2624
rect 9862 2680 9918 2689
rect 9862 2615 9918 2624
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9600 2417 9628 2518
rect 9586 2408 9642 2417
rect 9876 2378 9904 2615
rect 9586 2343 9642 2352
rect 9864 2372 9916 2378
rect 9864 2314 9916 2320
rect 9772 2304 9824 2310
rect 9586 2272 9642 2281
rect 9772 2246 9824 2252
rect 9586 2207 9642 2216
rect 9600 1834 9628 2207
rect 9588 1828 9640 1834
rect 9588 1770 9640 1776
rect 9784 1766 9812 2246
rect 9772 1760 9824 1766
rect 9772 1702 9824 1708
rect 9416 1414 9628 1442
rect 9600 480 9628 1414
rect 9968 480 9996 2751
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10060 2310 10088 2586
rect 10152 2582 10180 4966
rect 10244 4865 10272 5086
rect 10230 4856 10286 4865
rect 10230 4791 10286 4800
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10244 2650 10272 4422
rect 10336 4282 10364 6734
rect 10428 5574 10456 7919
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10428 4758 10456 5102
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10322 4176 10378 4185
rect 10428 4146 10456 4558
rect 10322 4111 10324 4120
rect 10376 4111 10378 4120
rect 10416 4140 10468 4146
rect 10324 4082 10376 4088
rect 10416 4082 10468 4088
rect 10336 3602 10364 4082
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10428 3777 10456 3878
rect 10414 3768 10470 3777
rect 10414 3703 10470 3712
rect 10414 3632 10470 3641
rect 10324 3596 10376 3602
rect 10414 3567 10470 3576
rect 10324 3538 10376 3544
rect 10428 3466 10456 3567
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10414 3224 10470 3233
rect 10520 3210 10548 9132
rect 10612 7410 10640 10492
rect 10980 10452 11008 10678
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11072 10577 11100 10610
rect 11058 10568 11114 10577
rect 11058 10503 11114 10512
rect 10704 10424 11008 10452
rect 10704 10198 10732 10424
rect 10817 10364 11113 10384
rect 10873 10362 10897 10364
rect 10953 10362 10977 10364
rect 11033 10362 11057 10364
rect 10895 10310 10897 10362
rect 10959 10310 10971 10362
rect 11033 10310 11035 10362
rect 10873 10308 10897 10310
rect 10953 10308 10977 10310
rect 11033 10308 11057 10310
rect 10817 10288 11113 10308
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10612 6934 10640 7210
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10704 6254 10732 9590
rect 10782 9480 10838 9489
rect 10782 9415 10784 9424
rect 10836 9415 10838 9424
rect 10784 9386 10836 9392
rect 11072 9364 11100 10134
rect 11164 9518 11192 10911
rect 11256 10713 11284 11698
rect 11348 11218 11376 11727
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11242 10704 11298 10713
rect 11348 10674 11376 10746
rect 11532 10742 11560 15506
rect 11624 14822 11652 19520
rect 11886 17504 11942 17513
rect 11886 17439 11942 17448
rect 11900 16522 11928 17439
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11716 14890 11744 15506
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11624 13841 11652 14418
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11610 13832 11666 13841
rect 11610 13767 11666 13776
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11624 13258 11652 13670
rect 11716 13258 11744 14214
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11702 13152 11758 13161
rect 11702 13087 11758 13096
rect 11610 13016 11666 13025
rect 11610 12951 11666 12960
rect 11520 10736 11572 10742
rect 11520 10678 11572 10684
rect 11242 10639 11298 10648
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11242 10568 11298 10577
rect 11242 10503 11298 10512
rect 11256 9586 11284 10503
rect 11624 10266 11652 12951
rect 11716 12764 11744 13087
rect 11808 12889 11836 15982
rect 11992 13025 12020 19520
rect 12360 18086 12388 19520
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 11978 13016 12034 13025
rect 11978 12951 12034 12960
rect 11794 12880 11850 12889
rect 11794 12815 11850 12824
rect 11716 12736 11836 12764
rect 11704 12640 11756 12646
rect 11702 12608 11704 12617
rect 11756 12608 11758 12617
rect 11702 12543 11758 12552
rect 11702 12472 11758 12481
rect 11702 12407 11704 12416
rect 11756 12407 11758 12416
rect 11704 12378 11756 12384
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11716 11354 11744 12038
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11348 9897 11376 10202
rect 11520 10192 11572 10198
rect 11716 10146 11744 11154
rect 11808 10266 11836 12736
rect 12084 12646 12112 16662
rect 12176 16561 12204 16730
rect 12162 16552 12218 16561
rect 12162 16487 12218 16496
rect 12348 15972 12400 15978
rect 12348 15914 12400 15920
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 12176 15609 12204 15642
rect 12162 15600 12218 15609
rect 12162 15535 12218 15544
rect 12162 15464 12218 15473
rect 12162 15399 12218 15408
rect 12176 14890 12204 15399
rect 12254 15192 12310 15201
rect 12254 15127 12256 15136
rect 12308 15127 12310 15136
rect 12256 15098 12308 15104
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12268 12730 12296 14758
rect 12176 12702 12296 12730
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 11886 12472 11942 12481
rect 11886 12407 11942 12416
rect 11900 11218 11928 12407
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11900 10742 11928 10950
rect 11888 10736 11940 10742
rect 11888 10678 11940 10684
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11572 10140 11652 10146
rect 11520 10134 11652 10140
rect 11532 10118 11652 10134
rect 11716 10118 11836 10146
rect 11624 10010 11652 10118
rect 11532 9982 11652 10010
rect 11334 9888 11390 9897
rect 11334 9823 11390 9832
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11152 9512 11204 9518
rect 11428 9512 11480 9518
rect 11152 9454 11204 9460
rect 11426 9480 11428 9489
rect 11480 9480 11482 9489
rect 11426 9415 11482 9424
rect 11336 9376 11388 9382
rect 11072 9336 11192 9364
rect 10817 9276 11113 9296
rect 10873 9274 10897 9276
rect 10953 9274 10977 9276
rect 11033 9274 11057 9276
rect 10895 9222 10897 9274
rect 10959 9222 10971 9274
rect 11033 9222 11035 9274
rect 10873 9220 10897 9222
rect 10953 9220 10977 9222
rect 11033 9220 11057 9222
rect 10817 9200 11113 9220
rect 10784 9104 10836 9110
rect 10784 9046 10836 9052
rect 10796 8809 10824 9046
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10782 8800 10838 8809
rect 10782 8735 10838 8744
rect 10980 8566 11008 8842
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 8634 11100 8774
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10817 8188 11113 8208
rect 10873 8186 10897 8188
rect 10953 8186 10977 8188
rect 11033 8186 11057 8188
rect 10895 8134 10897 8186
rect 10959 8134 10971 8186
rect 11033 8134 11035 8186
rect 10873 8132 10897 8134
rect 10953 8132 10977 8134
rect 11033 8132 11057 8134
rect 10817 8112 11113 8132
rect 11164 8090 11192 9336
rect 11336 9318 11388 9324
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11348 9178 11376 9318
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11256 8634 11284 8978
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11348 8498 11376 8910
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11440 8378 11468 9318
rect 11532 8412 11560 9982
rect 11702 9888 11758 9897
rect 11702 9823 11758 9832
rect 11716 9722 11744 9823
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11612 8560 11664 8566
rect 11716 8548 11744 9386
rect 11664 8520 11744 8548
rect 11612 8502 11664 8508
rect 11532 8384 11652 8412
rect 11256 8350 11468 8378
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11256 7970 11284 8350
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11348 8090 11376 8230
rect 11532 8129 11560 8230
rect 11518 8120 11574 8129
rect 11336 8084 11388 8090
rect 11518 8055 11574 8064
rect 11336 8026 11388 8032
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10888 7942 11284 7970
rect 10796 7188 10824 7890
rect 10888 7585 10916 7942
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10874 7576 10930 7585
rect 10874 7511 10930 7520
rect 10980 7290 11008 7754
rect 11072 7410 11100 7822
rect 11164 7585 11192 7822
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11150 7576 11206 7585
rect 11150 7511 11206 7520
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11164 7290 11192 7414
rect 10980 7262 11192 7290
rect 10796 7160 11192 7188
rect 10817 7100 11113 7120
rect 10873 7098 10897 7100
rect 10953 7098 10977 7100
rect 11033 7098 11057 7100
rect 10895 7046 10897 7098
rect 10959 7046 10971 7098
rect 11033 7046 11035 7098
rect 10873 7044 10897 7046
rect 10953 7044 10977 7046
rect 11033 7044 11057 7046
rect 10817 7024 11113 7044
rect 11164 7002 11192 7160
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 10966 6896 11022 6905
rect 10966 6831 11022 6840
rect 11150 6896 11206 6905
rect 11150 6831 11206 6840
rect 10980 6662 11008 6831
rect 11164 6798 11192 6831
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10600 6180 10652 6186
rect 10600 6122 10652 6128
rect 10612 5914 10640 6122
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10704 5137 10732 5238
rect 10690 5128 10746 5137
rect 10600 5092 10652 5098
rect 10796 5098 10824 5714
rect 11164 5642 11192 6258
rect 11256 5953 11284 7686
rect 11532 7460 11560 7822
rect 11440 7432 11560 7460
rect 11440 6798 11468 7432
rect 11520 6928 11572 6934
rect 11520 6870 11572 6876
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11242 5944 11298 5953
rect 11242 5879 11244 5888
rect 11296 5879 11298 5888
rect 11244 5850 11296 5856
rect 11532 5658 11560 6870
rect 11152 5636 11204 5642
rect 11152 5578 11204 5584
rect 11256 5630 11560 5658
rect 11164 5302 11192 5578
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 10690 5063 10746 5072
rect 10784 5092 10836 5098
rect 10600 5034 10652 5040
rect 10612 3398 10640 5034
rect 10704 3942 10732 5063
rect 10784 5034 10836 5040
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10817 4848 11113 4868
rect 11164 4758 11192 5238
rect 10876 4752 10928 4758
rect 10876 4694 10928 4700
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10796 4010 10824 4626
rect 10888 4146 10916 4694
rect 11072 4604 11100 4694
rect 11256 4604 11284 5630
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11426 5400 11482 5409
rect 11426 5335 11482 5344
rect 11072 4576 11284 4604
rect 11440 4536 11468 5335
rect 11256 4508 11468 4536
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10520 3182 10640 3210
rect 10414 3159 10470 3168
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 10336 480 10364 3062
rect 10428 2854 10456 3159
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10612 480 10640 3182
rect 10704 2514 10732 3878
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 11164 2990 11192 4422
rect 11256 3913 11284 4508
rect 11426 4448 11482 4457
rect 11426 4383 11482 4392
rect 11334 4312 11390 4321
rect 11334 4247 11390 4256
rect 11348 4010 11376 4247
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 11242 3904 11298 3913
rect 11242 3839 11298 3848
rect 11256 3516 11284 3839
rect 11440 3602 11468 4383
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11336 3528 11388 3534
rect 11256 3488 11336 3516
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11256 2854 11284 3488
rect 11336 3470 11388 3476
rect 11532 3194 11560 5510
rect 11624 5030 11652 8384
rect 11808 8294 11836 10118
rect 11900 10062 11928 10474
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11992 9908 12020 12242
rect 12070 11520 12126 11529
rect 12070 11455 12126 11464
rect 12084 10198 12112 11455
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 11900 9880 12020 9908
rect 12070 9888 12126 9897
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11702 8120 11758 8129
rect 11702 8055 11758 8064
rect 11716 6866 11744 8055
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11808 7585 11836 7958
rect 11794 7576 11850 7585
rect 11794 7511 11850 7520
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11716 6390 11744 6598
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11624 3534 11652 4558
rect 11716 3942 11744 6054
rect 11808 5166 11836 7511
rect 11900 5778 11928 9880
rect 12070 9823 12126 9832
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11992 8673 12020 9318
rect 11978 8664 12034 8673
rect 11978 8599 12034 8608
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11992 5370 12020 8599
rect 12084 8129 12112 9823
rect 12070 8120 12126 8129
rect 12070 8055 12126 8064
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11808 4282 11836 4762
rect 11900 4758 11928 5034
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11992 4298 12020 5102
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11900 4270 12020 4298
rect 11796 4072 11848 4078
rect 11900 4049 11928 4270
rect 11980 4072 12032 4078
rect 11796 4014 11848 4020
rect 11886 4040 11942 4049
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11624 3074 11652 3130
rect 11348 3046 11652 3074
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10817 2672 11113 2692
rect 11348 2650 11376 3046
rect 11520 2984 11572 2990
rect 11716 2972 11744 3606
rect 11808 2990 11836 4014
rect 11980 4014 12032 4020
rect 11886 3975 11942 3984
rect 11992 3670 12020 4014
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11520 2926 11572 2932
rect 11624 2944 11744 2972
rect 11796 2984 11848 2990
rect 11532 2825 11560 2926
rect 11518 2816 11574 2825
rect 11518 2751 11574 2760
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 11336 2304 11388 2310
rect 10966 2272 11022 2281
rect 11336 2246 11388 2252
rect 10966 2207 11022 2216
rect 10980 480 11008 2207
rect 11348 480 11376 2246
rect 11440 1630 11468 2586
rect 11532 1698 11560 2751
rect 11520 1692 11572 1698
rect 11520 1634 11572 1640
rect 11428 1624 11480 1630
rect 11428 1566 11480 1572
rect 11624 480 11652 2944
rect 11796 2926 11848 2932
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11808 2106 11836 2450
rect 11900 2378 11928 3538
rect 12084 3398 12112 7686
rect 12176 6322 12204 12702
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12268 12481 12296 12582
rect 12254 12472 12310 12481
rect 12254 12407 12310 12416
rect 12360 12374 12388 15914
rect 12256 12368 12308 12374
rect 12256 12310 12308 12316
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 12268 12186 12296 12310
rect 12268 12158 12388 12186
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12268 9382 12296 12038
rect 12360 11665 12388 12158
rect 12452 11801 12480 17070
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12544 16561 12572 16594
rect 12530 16552 12586 16561
rect 12530 16487 12586 16496
rect 12636 15745 12664 19520
rect 12808 17944 12860 17950
rect 12808 17886 12860 17892
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12728 16402 12756 17546
rect 12820 16522 12848 17886
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12912 17338 12940 17478
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12728 16374 12848 16402
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12622 15736 12678 15745
rect 12622 15671 12678 15680
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12544 13870 12572 15370
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12544 12918 12572 13330
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12544 12442 12572 12854
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12530 12064 12586 12073
rect 12530 11999 12586 12008
rect 12438 11792 12494 11801
rect 12438 11727 12494 11736
rect 12346 11656 12402 11665
rect 12346 11591 12402 11600
rect 12348 11552 12400 11558
rect 12400 11500 12480 11506
rect 12348 11494 12480 11500
rect 12360 11478 12480 11494
rect 12452 11393 12480 11478
rect 12438 11384 12494 11393
rect 12438 11319 12494 11328
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12452 10985 12480 11154
rect 12438 10976 12494 10985
rect 12438 10911 12494 10920
rect 12544 10674 12572 11999
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12440 10600 12492 10606
rect 12438 10568 12440 10577
rect 12492 10568 12494 10577
rect 12438 10503 12494 10512
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12268 7954 12296 9046
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 12176 3210 12204 5306
rect 12268 5114 12296 7754
rect 12360 7154 12388 10066
rect 12452 9625 12480 10406
rect 12544 9722 12572 10610
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12438 9616 12494 9625
rect 12438 9551 12494 9560
rect 12544 9489 12572 9658
rect 12530 9480 12586 9489
rect 12530 9415 12586 9424
rect 12636 9364 12664 13330
rect 12728 12628 12756 15982
rect 12820 14074 12848 16374
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12912 13954 12940 17070
rect 12820 13926 12940 13954
rect 12820 13394 12848 13926
rect 13004 13818 13032 19520
rect 13372 18018 13400 19520
rect 13360 18012 13412 18018
rect 13360 17954 13412 17960
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 13188 16697 13216 17682
rect 13282 17436 13578 17456
rect 13338 17434 13362 17436
rect 13418 17434 13442 17436
rect 13498 17434 13522 17436
rect 13360 17382 13362 17434
rect 13424 17382 13436 17434
rect 13498 17382 13500 17434
rect 13338 17380 13362 17382
rect 13418 17380 13442 17382
rect 13498 17380 13522 17382
rect 13282 17360 13578 17380
rect 13740 17218 13768 19520
rect 13740 17190 13860 17218
rect 13360 17128 13412 17134
rect 13358 17096 13360 17105
rect 13412 17096 13414 17105
rect 13358 17031 13414 17040
rect 13174 16688 13230 16697
rect 13174 16623 13230 16632
rect 13282 16348 13578 16368
rect 13338 16346 13362 16348
rect 13418 16346 13442 16348
rect 13498 16346 13522 16348
rect 13360 16294 13362 16346
rect 13424 16294 13436 16346
rect 13498 16294 13500 16346
rect 13338 16292 13362 16294
rect 13418 16292 13442 16294
rect 13498 16292 13522 16294
rect 13282 16272 13578 16292
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13188 15609 13216 15982
rect 13174 15600 13230 15609
rect 13174 15535 13230 15544
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 12912 13790 13032 13818
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12820 12850 12848 13194
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12808 12640 12860 12646
rect 12728 12600 12808 12628
rect 12808 12582 12860 12588
rect 12820 12102 12848 12582
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12714 11928 12770 11937
rect 12714 11863 12770 11872
rect 12728 11830 12756 11863
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12912 11642 12940 13790
rect 13096 13530 13124 14758
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 13188 13410 13216 15438
rect 13282 15260 13578 15280
rect 13338 15258 13362 15260
rect 13418 15258 13442 15260
rect 13498 15258 13522 15260
rect 13360 15206 13362 15258
rect 13424 15206 13436 15258
rect 13498 15206 13500 15258
rect 13338 15204 13362 15206
rect 13418 15204 13442 15206
rect 13498 15204 13522 15206
rect 13282 15184 13578 15204
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13282 14172 13578 14192
rect 13338 14170 13362 14172
rect 13418 14170 13442 14172
rect 13498 14170 13522 14172
rect 13360 14118 13362 14170
rect 13424 14118 13436 14170
rect 13498 14118 13500 14170
rect 13338 14116 13362 14118
rect 13418 14116 13442 14118
rect 13498 14116 13522 14118
rect 13282 14096 13578 14116
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13280 13530 13308 13806
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 12820 11614 12940 11642
rect 13004 13382 13216 13410
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12452 9336 12664 9364
rect 12452 8090 12480 9336
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12544 8809 12572 8978
rect 12624 8832 12676 8838
rect 12530 8800 12586 8809
rect 12624 8774 12676 8780
rect 12530 8735 12586 8744
rect 12530 8392 12586 8401
rect 12530 8327 12586 8336
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12452 7585 12480 8026
rect 12438 7576 12494 7585
rect 12438 7511 12494 7520
rect 12544 7206 12572 8327
rect 12636 8129 12664 8774
rect 12622 8120 12678 8129
rect 12622 8055 12678 8064
rect 12728 7800 12756 11018
rect 12820 9178 12848 11614
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 9217 12940 11494
rect 12898 9208 12954 9217
rect 12808 9172 12860 9178
rect 12898 9143 12954 9152
rect 12808 9114 12860 9120
rect 12820 8537 12848 9114
rect 12900 8560 12952 8566
rect 12806 8528 12862 8537
rect 12900 8502 12952 8508
rect 12806 8463 12862 8472
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12636 7772 12756 7800
rect 12636 7562 12664 7772
rect 12636 7534 12756 7562
rect 12728 7410 12756 7534
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12820 7342 12848 8230
rect 12912 7886 12940 8502
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12898 7576 12954 7585
rect 12898 7511 12954 7520
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12532 7200 12584 7206
rect 12360 7126 12480 7154
rect 12808 7200 12860 7206
rect 12532 7142 12584 7148
rect 12806 7168 12808 7177
rect 12860 7168 12862 7177
rect 12452 6882 12480 7126
rect 12806 7103 12862 7112
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12360 6854 12480 6882
rect 12360 6610 12388 6854
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12360 6582 12480 6610
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12360 5216 12388 6258
rect 12452 6225 12480 6582
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12438 6216 12494 6225
rect 12438 6151 12494 6160
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12452 5846 12480 6054
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12360 5188 12480 5216
rect 12268 5086 12388 5114
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 11992 3182 12204 3210
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 11992 480 12020 3182
rect 12268 2310 12296 4966
rect 12360 4826 12388 5086
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12360 4146 12388 4762
rect 12452 4214 12480 5188
rect 12544 5098 12572 6258
rect 12728 6202 12756 6734
rect 12636 6174 12756 6202
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 12544 4146 12572 5034
rect 12636 4826 12664 6174
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12728 5914 12756 6054
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12820 5681 12848 6938
rect 12912 6322 12940 7511
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12806 5672 12862 5681
rect 12806 5607 12862 5616
rect 12808 5568 12860 5574
rect 12714 5536 12770 5545
rect 12808 5510 12860 5516
rect 12714 5471 12770 5480
rect 12728 5030 12756 5471
rect 12820 5234 12848 5510
rect 12912 5370 12940 6054
rect 13004 5914 13032 13382
rect 13464 13308 13492 13942
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13556 13326 13584 13874
rect 13096 13280 13492 13308
rect 13544 13320 13596 13326
rect 13096 11354 13124 13280
rect 13544 13262 13596 13268
rect 13282 13084 13578 13104
rect 13338 13082 13362 13084
rect 13418 13082 13442 13084
rect 13498 13082 13522 13084
rect 13360 13030 13362 13082
rect 13424 13030 13436 13082
rect 13498 13030 13500 13082
rect 13338 13028 13362 13030
rect 13418 13028 13442 13030
rect 13498 13028 13522 13030
rect 13282 13008 13578 13028
rect 13450 12880 13506 12889
rect 13648 12850 13676 14418
rect 13740 13569 13768 14758
rect 13832 14074 13860 17190
rect 13910 16008 13966 16017
rect 13910 15943 13966 15952
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13818 13968 13874 13977
rect 13818 13903 13874 13912
rect 13832 13870 13860 13903
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13726 13560 13782 13569
rect 13726 13495 13782 13504
rect 13726 13424 13782 13433
rect 13726 13359 13782 13368
rect 13740 13326 13768 13359
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13726 13152 13782 13161
rect 13726 13087 13782 13096
rect 13450 12815 13506 12824
rect 13636 12844 13688 12850
rect 13464 12306 13492 12815
rect 13636 12786 13688 12792
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13188 11898 13216 12174
rect 13282 11996 13578 12016
rect 13338 11994 13362 11996
rect 13418 11994 13442 11996
rect 13498 11994 13522 11996
rect 13360 11942 13362 11994
rect 13424 11942 13436 11994
rect 13498 11942 13500 11994
rect 13338 11940 13362 11942
rect 13418 11940 13442 11942
rect 13498 11940 13522 11942
rect 13282 11920 13578 11940
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13082 11112 13138 11121
rect 13082 11047 13138 11056
rect 13096 8634 13124 11047
rect 13188 9518 13216 11562
rect 13556 11082 13584 11698
rect 13740 11694 13768 13087
rect 13832 11694 13860 13806
rect 13924 13394 13952 15943
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13740 11286 13768 11630
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13282 10908 13578 10928
rect 13338 10906 13362 10908
rect 13418 10906 13442 10908
rect 13498 10906 13522 10908
rect 13360 10854 13362 10906
rect 13424 10854 13436 10906
rect 13498 10854 13500 10906
rect 13338 10852 13362 10854
rect 13418 10852 13442 10854
rect 13498 10852 13522 10854
rect 13282 10832 13578 10852
rect 13648 10810 13676 11154
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13450 10432 13506 10441
rect 13450 10367 13506 10376
rect 13464 10198 13492 10367
rect 13452 10192 13504 10198
rect 13358 10160 13414 10169
rect 13452 10134 13504 10140
rect 13358 10095 13360 10104
rect 13412 10095 13414 10104
rect 13360 10066 13412 10072
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13556 9908 13584 9998
rect 13648 9976 13676 10610
rect 13740 10266 13768 11086
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13820 10192 13872 10198
rect 13726 10160 13782 10169
rect 13820 10134 13872 10140
rect 13726 10095 13728 10104
rect 13780 10095 13782 10104
rect 13728 10066 13780 10072
rect 13728 9988 13780 9994
rect 13648 9948 13728 9976
rect 13728 9930 13780 9936
rect 13556 9880 13676 9908
rect 13282 9820 13578 9840
rect 13338 9818 13362 9820
rect 13418 9818 13442 9820
rect 13498 9818 13522 9820
rect 13360 9766 13362 9818
rect 13424 9766 13436 9818
rect 13498 9766 13500 9818
rect 13338 9764 13362 9766
rect 13418 9764 13442 9766
rect 13498 9764 13522 9766
rect 13282 9744 13578 9764
rect 13648 9704 13676 9880
rect 13556 9676 13676 9704
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 13176 9376 13228 9382
rect 13174 9344 13176 9353
rect 13228 9344 13230 9353
rect 13174 9279 13230 9288
rect 13174 9208 13230 9217
rect 13174 9143 13176 9152
rect 13228 9143 13230 9152
rect 13176 9114 13228 9120
rect 13280 9081 13308 9386
rect 13464 9178 13492 9590
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13266 9072 13322 9081
rect 13176 9036 13228 9042
rect 13556 9058 13584 9676
rect 13740 9450 13768 9930
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13556 9030 13676 9058
rect 13266 9007 13322 9016
rect 13176 8978 13228 8984
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12992 5636 13044 5642
rect 12992 5578 13044 5584
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12728 4706 12756 4966
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12636 4678 12756 4706
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12346 4040 12402 4049
rect 12346 3975 12402 3984
rect 12360 3738 12388 3975
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12452 3369 12480 3470
rect 12636 3398 12664 4678
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12624 3392 12676 3398
rect 12438 3360 12494 3369
rect 12624 3334 12676 3340
rect 12438 3295 12494 3304
rect 12346 3224 12402 3233
rect 12346 3159 12402 3168
rect 12622 3224 12678 3233
rect 12622 3159 12678 3168
rect 12360 2530 12388 3159
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 2650 12480 2790
rect 12544 2689 12572 2858
rect 12530 2680 12586 2689
rect 12440 2644 12492 2650
rect 12530 2615 12586 2624
rect 12440 2586 12492 2592
rect 12530 2544 12586 2553
rect 12360 2514 12480 2530
rect 12360 2508 12492 2514
rect 12360 2502 12440 2508
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12360 480 12388 2502
rect 12530 2479 12586 2488
rect 12440 2450 12492 2456
rect 12544 2446 12572 2479
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12636 480 12664 3159
rect 12728 2582 12756 4558
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 12820 2378 12848 4762
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 12912 3670 12940 4218
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 2428 12940 3334
rect 13004 2854 13032 5578
rect 13096 5370 13124 8298
rect 13188 8265 13216 8978
rect 13282 8732 13578 8752
rect 13338 8730 13362 8732
rect 13418 8730 13442 8732
rect 13498 8730 13522 8732
rect 13360 8678 13362 8730
rect 13424 8678 13436 8730
rect 13498 8678 13500 8730
rect 13338 8676 13362 8678
rect 13418 8676 13442 8678
rect 13498 8676 13522 8678
rect 13282 8656 13578 8676
rect 13174 8256 13230 8265
rect 13174 8191 13230 8200
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13096 5030 13124 5170
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13188 4826 13216 7890
rect 13266 7848 13322 7857
rect 13266 7783 13268 7792
rect 13320 7783 13322 7792
rect 13268 7754 13320 7760
rect 13282 7644 13578 7664
rect 13338 7642 13362 7644
rect 13418 7642 13442 7644
rect 13498 7642 13522 7644
rect 13360 7590 13362 7642
rect 13424 7590 13436 7642
rect 13498 7590 13500 7642
rect 13338 7588 13362 7590
rect 13418 7588 13442 7590
rect 13498 7588 13522 7590
rect 13282 7568 13578 7588
rect 13648 7410 13676 9030
rect 13740 8906 13768 9386
rect 13832 8922 13860 10134
rect 13924 9586 13952 13194
rect 14016 12646 14044 19520
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14292 16794 14320 17614
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14384 16454 14412 19520
rect 14556 17808 14608 17814
rect 14556 17750 14608 17756
rect 14372 16448 14424 16454
rect 14292 16408 14372 16436
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 14200 16153 14228 16186
rect 14186 16144 14242 16153
rect 14186 16079 14242 16088
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14108 14618 14136 14826
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14108 12186 14136 13670
rect 14200 13190 14228 14010
rect 14292 13258 14320 16408
rect 14372 16390 14424 16396
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14016 12158 14136 12186
rect 14016 11626 14044 12158
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14004 11620 14056 11626
rect 14004 11562 14056 11568
rect 14016 9926 14044 11562
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 13912 9580 13964 9586
rect 13964 9540 14044 9568
rect 13912 9522 13964 9528
rect 13910 9480 13966 9489
rect 13910 9415 13966 9424
rect 13924 9382 13952 9415
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13728 8900 13780 8906
rect 13832 8894 13952 8922
rect 13728 8842 13780 8848
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13636 7404 13688 7410
rect 13556 7364 13636 7392
rect 13556 6644 13584 7364
rect 13636 7346 13688 7352
rect 13740 7342 13768 8366
rect 13728 7336 13780 7342
rect 13634 7304 13690 7313
rect 13728 7278 13780 7284
rect 13634 7239 13690 7248
rect 13648 7206 13676 7239
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13728 6928 13780 6934
rect 13832 6905 13860 8774
rect 13924 8673 13952 8894
rect 13910 8664 13966 8673
rect 13910 8599 13966 8608
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13728 6870 13780 6876
rect 13818 6896 13874 6905
rect 13556 6616 13676 6644
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13452 6384 13504 6390
rect 13450 6352 13452 6361
rect 13504 6352 13506 6361
rect 13450 6287 13506 6296
rect 13648 5896 13676 6616
rect 13556 5868 13676 5896
rect 13556 5710 13584 5868
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13450 5264 13506 5273
rect 13450 5199 13506 5208
rect 13464 5098 13492 5199
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13358 4720 13414 4729
rect 13358 4655 13360 4664
rect 13412 4655 13414 4664
rect 13360 4626 13412 4632
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 13096 4146 13124 4490
rect 13282 4380 13578 4400
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 13176 4208 13228 4214
rect 13452 4208 13504 4214
rect 13176 4150 13228 4156
rect 13358 4176 13414 4185
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13096 3534 13124 4082
rect 13188 3670 13216 4150
rect 13452 4150 13504 4156
rect 13358 4111 13414 4120
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 13280 3913 13308 3946
rect 13266 3904 13322 3913
rect 13266 3839 13322 3848
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13188 3194 13216 3606
rect 13372 3466 13400 4111
rect 13464 3738 13492 4150
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 12992 2848 13044 2854
rect 13176 2848 13228 2854
rect 13044 2808 13124 2836
rect 12992 2790 13044 2796
rect 12990 2680 13046 2689
rect 12990 2615 13046 2624
rect 13004 2582 13032 2615
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 12912 2400 13032 2428
rect 12808 2372 12860 2378
rect 12808 2314 12860 2320
rect 13004 480 13032 2400
rect 13096 1562 13124 2808
rect 13176 2790 13228 2796
rect 13188 2088 13216 2790
rect 13280 2417 13308 2858
rect 13464 2666 13492 2858
rect 13648 2854 13676 5714
rect 13740 3194 13768 6870
rect 13818 6831 13874 6840
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13832 5817 13860 6666
rect 13818 5808 13874 5817
rect 13818 5743 13874 5752
rect 13924 5658 13952 8366
rect 14016 7954 14044 9540
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14004 7812 14056 7818
rect 14004 7754 14056 7760
rect 14016 6322 14044 7754
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 13832 5630 13952 5658
rect 13832 3942 13860 5630
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13924 4282 13952 5510
rect 14016 5370 14044 6054
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 14002 4584 14058 4593
rect 14002 4519 14058 4528
rect 14016 4486 14044 4519
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 14016 4026 14044 4082
rect 13924 3998 14044 4026
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13832 3074 13860 3402
rect 13740 3058 13860 3074
rect 13728 3052 13860 3058
rect 13780 3046 13860 3052
rect 13728 2994 13780 3000
rect 13636 2848 13688 2854
rect 13924 2825 13952 3998
rect 14108 3482 14136 12038
rect 14200 10130 14228 12786
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14200 8650 14228 10066
rect 14292 9042 14320 12854
rect 14384 10606 14412 14758
rect 14568 13802 14596 17750
rect 14646 17640 14702 17649
rect 14646 17575 14702 17584
rect 14556 13796 14608 13802
rect 14556 13738 14608 13744
rect 14556 12300 14608 12306
rect 14476 12260 14556 12288
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14384 9518 14412 10406
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14200 8622 14320 8650
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14200 7886 14228 8366
rect 14292 8362 14320 8622
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14200 7546 14228 7822
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14292 7018 14320 8298
rect 14200 6990 14320 7018
rect 14200 5914 14228 6990
rect 14384 6866 14412 9454
rect 14476 8566 14504 12260
rect 14556 12242 14608 12248
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14568 8430 14596 12106
rect 14660 10538 14688 17575
rect 14752 12170 14780 19520
rect 15028 16402 15056 19520
rect 15028 16374 15332 16402
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 14832 12776 14884 12782
rect 14830 12744 14832 12753
rect 14884 12744 14886 12753
rect 14830 12679 14886 12688
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14844 12306 14872 12582
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14936 11914 14964 13942
rect 15120 13274 15148 16186
rect 15028 13246 15148 13274
rect 15028 12850 15056 13246
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 14752 11886 14964 11914
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14646 10024 14702 10033
rect 14646 9959 14648 9968
rect 14700 9959 14702 9968
rect 14648 9930 14700 9936
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14568 7993 14596 8366
rect 14554 7984 14610 7993
rect 14554 7919 14610 7928
rect 14660 7834 14688 9658
rect 14568 7806 14688 7834
rect 14568 7290 14596 7806
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14660 7449 14688 7686
rect 14646 7440 14702 7449
rect 14646 7375 14702 7384
rect 14568 7262 14688 7290
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14200 5681 14228 5714
rect 14186 5672 14242 5681
rect 14186 5607 14242 5616
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14200 4622 14228 5102
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14016 3454 14136 3482
rect 13636 2790 13688 2796
rect 13910 2816 13966 2825
rect 13910 2751 13966 2760
rect 13464 2638 13768 2666
rect 13266 2408 13322 2417
rect 13266 2343 13322 2352
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 13188 2060 13400 2088
rect 13084 1556 13136 1562
rect 13084 1498 13136 1504
rect 13372 480 13400 2060
rect 13740 480 13768 2638
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 13912 2304 13964 2310
rect 13912 2246 13964 2252
rect 13832 2038 13860 2246
rect 13820 2032 13872 2038
rect 13820 1974 13872 1980
rect 13924 1834 13952 2246
rect 13912 1828 13964 1834
rect 13912 1770 13964 1776
rect 14016 480 14044 3454
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 3058 14136 3334
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14200 2650 14228 4218
rect 14292 3058 14320 6258
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14384 4282 14412 5306
rect 14476 5137 14504 5646
rect 14462 5128 14518 5137
rect 14462 5063 14518 5072
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14476 4214 14504 5063
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14384 480 14412 4082
rect 14568 4049 14596 7142
rect 14660 6866 14688 7262
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14660 5370 14688 6802
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14660 4622 14688 5170
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14648 4072 14700 4078
rect 14554 4040 14610 4049
rect 14648 4014 14700 4020
rect 14554 3975 14610 3984
rect 14462 3904 14518 3913
rect 14462 3839 14518 3848
rect 14476 3126 14504 3839
rect 14660 3641 14688 4014
rect 14646 3632 14702 3641
rect 14646 3567 14702 3576
rect 14646 3496 14702 3505
rect 14646 3431 14648 3440
rect 14700 3431 14702 3440
rect 14648 3402 14700 3408
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14476 2854 14504 3062
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14568 2446 14596 2994
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14752 480 14780 11886
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14844 2854 14872 11018
rect 14936 10033 14964 11698
rect 15028 10554 15056 12582
rect 15120 10690 15148 13126
rect 15304 11014 15332 16374
rect 15396 12918 15424 19520
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15120 10662 15240 10690
rect 15028 10526 15148 10554
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15028 10305 15056 10406
rect 15014 10296 15070 10305
rect 15014 10231 15070 10240
rect 14922 10024 14978 10033
rect 14922 9959 14978 9968
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14936 7818 14964 9862
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 15028 8945 15056 9318
rect 15014 8936 15070 8945
rect 15014 8871 15070 8880
rect 14924 7812 14976 7818
rect 14924 7754 14976 7760
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 14832 2848 14884 2854
rect 14832 2790 14884 2796
rect 14936 1766 14964 7210
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15028 6769 15056 7142
rect 15014 6760 15070 6769
rect 15014 6695 15070 6704
rect 15016 4208 15068 4214
rect 15014 4176 15016 4185
rect 15068 4176 15070 4185
rect 15014 4111 15070 4120
rect 15016 3120 15068 3126
rect 15014 3088 15016 3097
rect 15068 3088 15070 3097
rect 15014 3023 15070 3032
rect 15120 2972 15148 10526
rect 15212 9722 15240 10662
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15028 2944 15148 2972
rect 14924 1760 14976 1766
rect 14924 1702 14976 1708
rect 15028 480 15056 2944
rect 15212 2514 15240 9046
rect 15304 5234 15332 10950
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15396 480 15424 12174
rect 15488 4146 15516 14214
rect 15764 13734 15792 19520
rect 16040 17649 16068 19520
rect 16026 17640 16082 17649
rect 16026 17575 16082 17584
rect 16408 16250 16436 19520
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15580 6089 15608 8230
rect 15672 6254 15700 10134
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 15566 6080 15622 6089
rect 15566 6015 15622 6024
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15764 480 15792 12650
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16028 1964 16080 1970
rect 16028 1906 16080 1912
rect 16040 480 16068 1906
rect 16408 480 16436 11562
rect 16776 10606 16804 19520
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16762 2952 16818 2961
rect 16762 2887 16818 2896
rect 16776 480 16804 2887
rect 2870 439 2926 448
rect 3146 0 3202 480
rect 3514 0 3570 480
rect 3790 0 3846 480
rect 4158 0 4214 480
rect 4526 0 4582 480
rect 4802 0 4858 480
rect 5170 0 5226 480
rect 5538 0 5594 480
rect 5814 0 5870 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7194 0 7250 480
rect 7562 0 7618 480
rect 7930 0 7986 480
rect 8206 0 8262 480
rect 8574 0 8630 480
rect 8942 0 8998 480
rect 9218 0 9274 480
rect 9586 0 9642 480
rect 9954 0 10010 480
rect 10322 0 10378 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11610 0 11666 480
rect 11978 0 12034 480
rect 12346 0 12402 480
rect 12622 0 12678 480
rect 12990 0 13046 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14002 0 14058 480
rect 14370 0 14426 480
rect 14738 0 14794 480
rect 15014 0 15070 480
rect 15382 0 15438 480
rect 15750 0 15806 480
rect 16026 0 16082 480
rect 16394 0 16450 480
rect 16762 0 16818 480
<< via2 >>
rect 1490 19352 1546 19408
rect 1674 18400 1730 18456
rect 1214 8356 1270 8392
rect 1214 8336 1216 8356
rect 1216 8336 1268 8356
rect 1268 8336 1270 8356
rect 1674 7928 1730 7984
rect 1950 11056 2006 11112
rect 1858 10376 1914 10432
rect 1490 5344 1546 5400
rect 1858 7248 1914 7304
rect 1122 3032 1178 3088
rect 1766 3304 1822 3360
rect 1858 2916 1914 2952
rect 1858 2896 1860 2916
rect 1860 2896 1912 2916
rect 1912 2896 1914 2916
rect 2134 10648 2190 10704
rect 3421 17434 3477 17436
rect 3501 17434 3557 17436
rect 3581 17434 3637 17436
rect 3661 17434 3717 17436
rect 3421 17382 3447 17434
rect 3447 17382 3477 17434
rect 3501 17382 3511 17434
rect 3511 17382 3557 17434
rect 3581 17382 3627 17434
rect 3627 17382 3637 17434
rect 3661 17382 3691 17434
rect 3691 17382 3717 17434
rect 3421 17380 3477 17382
rect 3501 17380 3557 17382
rect 3581 17380 3637 17382
rect 3661 17380 3717 17382
rect 2962 17312 3018 17368
rect 2410 13912 2466 13968
rect 2870 16360 2926 16416
rect 2778 14456 2834 14512
rect 2870 13776 2926 13832
rect 2502 12844 2558 12880
rect 2502 12824 2504 12844
rect 2504 12824 2556 12844
rect 2556 12824 2558 12844
rect 2594 12724 2596 12744
rect 2596 12724 2648 12744
rect 2648 12724 2650 12744
rect 2594 12688 2650 12724
rect 2410 12280 2466 12336
rect 2594 10104 2650 10160
rect 2502 9560 2558 9616
rect 3330 16940 3332 16960
rect 3332 16940 3384 16960
rect 3384 16940 3386 16960
rect 3330 16904 3386 16940
rect 3421 16346 3477 16348
rect 3501 16346 3557 16348
rect 3581 16346 3637 16348
rect 3661 16346 3717 16348
rect 3421 16294 3447 16346
rect 3447 16294 3477 16346
rect 3501 16294 3511 16346
rect 3511 16294 3557 16346
rect 3581 16294 3627 16346
rect 3627 16294 3637 16346
rect 3661 16294 3691 16346
rect 3691 16294 3717 16346
rect 3421 16292 3477 16294
rect 3501 16292 3557 16294
rect 3581 16292 3637 16294
rect 3661 16292 3717 16294
rect 3606 15408 3662 15464
rect 3054 12280 3110 12336
rect 2410 8064 2466 8120
rect 2410 7928 2466 7984
rect 2134 6976 2190 7032
rect 2226 6180 2282 6216
rect 2226 6160 2228 6180
rect 2228 6160 2280 6180
rect 2280 6160 2282 6180
rect 2594 6296 2650 6352
rect 2962 8336 3018 8392
rect 3421 15258 3477 15260
rect 3501 15258 3557 15260
rect 3581 15258 3637 15260
rect 3661 15258 3717 15260
rect 3421 15206 3447 15258
rect 3447 15206 3477 15258
rect 3501 15206 3511 15258
rect 3511 15206 3557 15258
rect 3581 15206 3627 15258
rect 3627 15206 3637 15258
rect 3661 15206 3691 15258
rect 3691 15206 3717 15258
rect 3421 15204 3477 15206
rect 3501 15204 3557 15206
rect 3581 15204 3637 15206
rect 3661 15204 3717 15206
rect 3421 14170 3477 14172
rect 3501 14170 3557 14172
rect 3581 14170 3637 14172
rect 3661 14170 3717 14172
rect 3421 14118 3447 14170
rect 3447 14118 3477 14170
rect 3501 14118 3511 14170
rect 3511 14118 3557 14170
rect 3581 14118 3627 14170
rect 3627 14118 3637 14170
rect 3661 14118 3691 14170
rect 3691 14118 3717 14170
rect 3421 14116 3477 14118
rect 3501 14116 3557 14118
rect 3581 14116 3637 14118
rect 3661 14116 3717 14118
rect 3421 13082 3477 13084
rect 3501 13082 3557 13084
rect 3581 13082 3637 13084
rect 3661 13082 3717 13084
rect 3421 13030 3447 13082
rect 3447 13030 3477 13082
rect 3501 13030 3511 13082
rect 3511 13030 3557 13082
rect 3581 13030 3627 13082
rect 3627 13030 3637 13082
rect 3661 13030 3691 13082
rect 3691 13030 3717 13082
rect 3421 13028 3477 13030
rect 3501 13028 3557 13030
rect 3581 13028 3637 13030
rect 3661 13028 3717 13030
rect 3421 11994 3477 11996
rect 3501 11994 3557 11996
rect 3581 11994 3637 11996
rect 3661 11994 3717 11996
rect 3421 11942 3447 11994
rect 3447 11942 3477 11994
rect 3501 11942 3511 11994
rect 3511 11942 3557 11994
rect 3581 11942 3627 11994
rect 3627 11942 3637 11994
rect 3661 11942 3691 11994
rect 3691 11942 3717 11994
rect 3421 11940 3477 11942
rect 3501 11940 3557 11942
rect 3581 11940 3637 11942
rect 3661 11940 3717 11942
rect 3238 11328 3294 11384
rect 3054 7384 3110 7440
rect 3421 10906 3477 10908
rect 3501 10906 3557 10908
rect 3581 10906 3637 10908
rect 3661 10906 3717 10908
rect 3421 10854 3447 10906
rect 3447 10854 3477 10906
rect 3501 10854 3511 10906
rect 3511 10854 3557 10906
rect 3581 10854 3627 10906
rect 3627 10854 3637 10906
rect 3661 10854 3691 10906
rect 3691 10854 3717 10906
rect 3421 10852 3477 10854
rect 3501 10852 3557 10854
rect 3581 10852 3637 10854
rect 3661 10852 3717 10854
rect 3330 10376 3386 10432
rect 4342 15952 4398 16008
rect 4342 15000 4398 15056
rect 4986 16632 5042 16688
rect 4618 15408 4674 15464
rect 4066 14320 4122 14376
rect 4066 13504 4122 13560
rect 4894 14320 4950 14376
rect 4342 13096 4398 13152
rect 4894 12416 4950 12472
rect 3421 9818 3477 9820
rect 3501 9818 3557 9820
rect 3581 9818 3637 9820
rect 3661 9818 3717 9820
rect 3421 9766 3447 9818
rect 3447 9766 3477 9818
rect 3501 9766 3511 9818
rect 3511 9766 3557 9818
rect 3581 9766 3627 9818
rect 3627 9766 3637 9818
rect 3661 9766 3691 9818
rect 3691 9766 3717 9818
rect 3421 9764 3477 9766
rect 3501 9764 3557 9766
rect 3581 9764 3637 9766
rect 3661 9764 3717 9766
rect 3606 9288 3662 9344
rect 4066 10784 4122 10840
rect 4434 12008 4490 12064
rect 4526 11736 4582 11792
rect 4434 10376 4490 10432
rect 4434 10240 4490 10296
rect 3698 9152 3754 9208
rect 3698 9036 3754 9072
rect 3698 9016 3700 9036
rect 3700 9016 3752 9036
rect 3752 9016 3754 9036
rect 3421 8730 3477 8732
rect 3501 8730 3557 8732
rect 3581 8730 3637 8732
rect 3661 8730 3717 8732
rect 3421 8678 3447 8730
rect 3447 8678 3477 8730
rect 3501 8678 3511 8730
rect 3511 8678 3557 8730
rect 3581 8678 3627 8730
rect 3627 8678 3637 8730
rect 3661 8678 3691 8730
rect 3691 8678 3717 8730
rect 3421 8676 3477 8678
rect 3501 8676 3557 8678
rect 3581 8676 3637 8678
rect 3661 8676 3717 8678
rect 2962 6976 3018 7032
rect 2870 6432 2926 6488
rect 2134 4528 2190 4584
rect 1950 1400 2006 1456
rect 2226 3712 2282 3768
rect 2778 3984 2834 4040
rect 2962 3440 3018 3496
rect 3514 7928 3570 7984
rect 3421 7642 3477 7644
rect 3501 7642 3557 7644
rect 3581 7642 3637 7644
rect 3661 7642 3717 7644
rect 3421 7590 3447 7642
rect 3447 7590 3477 7642
rect 3501 7590 3511 7642
rect 3511 7590 3557 7642
rect 3581 7590 3627 7642
rect 3627 7590 3637 7642
rect 3661 7590 3691 7642
rect 3691 7590 3717 7642
rect 3421 7588 3477 7590
rect 3501 7588 3557 7590
rect 3581 7588 3637 7590
rect 3661 7588 3717 7590
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 3790 6160 3846 6216
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 3514 5072 3570 5128
rect 3238 4392 3294 4448
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 2870 448 2926 504
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 3974 8472 4030 8528
rect 3974 7656 4030 7712
rect 4250 9288 4306 9344
rect 4066 5652 4068 5672
rect 4068 5652 4120 5672
rect 4120 5652 4122 5672
rect 4066 5616 4122 5652
rect 4894 12008 4950 12064
rect 4710 10240 4766 10296
rect 4710 9968 4766 10024
rect 4526 9696 4582 9752
rect 4526 9288 4582 9344
rect 4434 6976 4490 7032
rect 4250 5208 4306 5264
rect 4342 4392 4398 4448
rect 4250 3304 4306 3360
rect 4342 3168 4398 3224
rect 4618 8472 4674 8528
rect 4986 9424 5042 9480
rect 5446 15544 5502 15600
rect 5886 16890 5942 16892
rect 5966 16890 6022 16892
rect 6046 16890 6102 16892
rect 6126 16890 6182 16892
rect 5886 16838 5912 16890
rect 5912 16838 5942 16890
rect 5966 16838 5976 16890
rect 5976 16838 6022 16890
rect 6046 16838 6092 16890
rect 6092 16838 6102 16890
rect 6126 16838 6156 16890
rect 6156 16838 6182 16890
rect 5886 16836 5942 16838
rect 5966 16836 6022 16838
rect 6046 16836 6102 16838
rect 6126 16836 6182 16838
rect 5814 16496 5870 16552
rect 5354 11600 5410 11656
rect 5354 10512 5410 10568
rect 5262 9716 5318 9752
rect 5262 9696 5264 9716
rect 5264 9696 5316 9716
rect 5316 9696 5318 9716
rect 4802 8900 4858 8936
rect 4802 8880 4804 8900
rect 4804 8880 4856 8900
rect 4856 8880 4858 8900
rect 4618 7928 4674 7984
rect 5170 9152 5226 9208
rect 4986 7384 5042 7440
rect 4802 7112 4858 7168
rect 4618 6452 4674 6488
rect 4618 6432 4620 6452
rect 4620 6432 4672 6452
rect 4672 6432 4674 6452
rect 4526 5752 4582 5808
rect 4066 2352 4122 2408
rect 4710 4664 4766 4720
rect 4618 3440 4674 3496
rect 5886 15802 5942 15804
rect 5966 15802 6022 15804
rect 6046 15802 6102 15804
rect 6126 15802 6182 15804
rect 5886 15750 5912 15802
rect 5912 15750 5942 15802
rect 5966 15750 5976 15802
rect 5976 15750 6022 15802
rect 6046 15750 6092 15802
rect 6092 15750 6102 15802
rect 6126 15750 6156 15802
rect 6156 15750 6182 15802
rect 5886 15748 5942 15750
rect 5966 15748 6022 15750
rect 6046 15748 6102 15750
rect 6126 15748 6182 15750
rect 6550 15544 6606 15600
rect 6550 15408 6606 15464
rect 5722 14864 5778 14920
rect 5722 13524 5778 13560
rect 5722 13504 5724 13524
rect 5724 13504 5776 13524
rect 5776 13504 5778 13524
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 6126 14714 6182 14716
rect 5886 14662 5912 14714
rect 5912 14662 5942 14714
rect 5966 14662 5976 14714
rect 5976 14662 6022 14714
rect 6046 14662 6092 14714
rect 6092 14662 6102 14714
rect 6126 14662 6156 14714
rect 6156 14662 6182 14714
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 6126 14660 6182 14662
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 6126 13626 6182 13628
rect 5886 13574 5912 13626
rect 5912 13574 5942 13626
rect 5966 13574 5976 13626
rect 5976 13574 6022 13626
rect 6046 13574 6092 13626
rect 6092 13574 6102 13626
rect 6126 13574 6156 13626
rect 6156 13574 6182 13626
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 6126 13572 6182 13574
rect 6182 12688 6238 12744
rect 6458 12552 6514 12608
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 6126 12538 6182 12540
rect 5886 12486 5912 12538
rect 5912 12486 5942 12538
rect 5966 12486 5976 12538
rect 5976 12486 6022 12538
rect 6046 12486 6092 12538
rect 6092 12486 6102 12538
rect 6126 12486 6156 12538
rect 6156 12486 6182 12538
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 6126 12484 6182 12486
rect 7286 14728 7342 14784
rect 7654 16940 7656 16960
rect 7656 16940 7708 16960
rect 7708 16940 7710 16960
rect 7654 16904 7710 16940
rect 8114 16088 8170 16144
rect 8352 17434 8408 17436
rect 8432 17434 8488 17436
rect 8512 17434 8568 17436
rect 8592 17434 8648 17436
rect 8352 17382 8378 17434
rect 8378 17382 8408 17434
rect 8432 17382 8442 17434
rect 8442 17382 8488 17434
rect 8512 17382 8558 17434
rect 8558 17382 8568 17434
rect 8592 17382 8622 17434
rect 8622 17382 8648 17434
rect 8352 17380 8408 17382
rect 8432 17380 8488 17382
rect 8512 17380 8568 17382
rect 8592 17380 8648 17382
rect 8574 16768 8630 16824
rect 8352 16346 8408 16348
rect 8432 16346 8488 16348
rect 8512 16346 8568 16348
rect 8592 16346 8648 16348
rect 8352 16294 8378 16346
rect 8378 16294 8408 16346
rect 8432 16294 8442 16346
rect 8442 16294 8488 16346
rect 8512 16294 8558 16346
rect 8558 16294 8568 16346
rect 8592 16294 8622 16346
rect 8622 16294 8648 16346
rect 8352 16292 8408 16294
rect 8432 16292 8488 16294
rect 8512 16292 8568 16294
rect 8592 16292 8648 16294
rect 8114 15408 8170 15464
rect 8352 15258 8408 15260
rect 8432 15258 8488 15260
rect 8512 15258 8568 15260
rect 8592 15258 8648 15260
rect 8352 15206 8378 15258
rect 8378 15206 8408 15258
rect 8432 15206 8442 15258
rect 8442 15206 8488 15258
rect 8512 15206 8558 15258
rect 8558 15206 8568 15258
rect 8592 15206 8622 15258
rect 8622 15206 8648 15258
rect 8352 15204 8408 15206
rect 8432 15204 8488 15206
rect 8512 15204 8568 15206
rect 8592 15204 8648 15206
rect 8942 17584 8998 17640
rect 8666 14592 8722 14648
rect 8352 14170 8408 14172
rect 8432 14170 8488 14172
rect 8512 14170 8568 14172
rect 8592 14170 8648 14172
rect 8352 14118 8378 14170
rect 8378 14118 8408 14170
rect 8432 14118 8442 14170
rect 8442 14118 8488 14170
rect 8512 14118 8558 14170
rect 8558 14118 8568 14170
rect 8592 14118 8622 14170
rect 8622 14118 8648 14170
rect 8352 14116 8408 14118
rect 8432 14116 8488 14118
rect 8512 14116 8568 14118
rect 8592 14116 8648 14118
rect 7746 13640 7802 13696
rect 7102 13504 7158 13560
rect 7010 13096 7066 13152
rect 6918 12960 6974 13016
rect 6734 12688 6790 12744
rect 5814 12144 5870 12200
rect 5630 11212 5686 11248
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 6126 11450 6182 11452
rect 5886 11398 5912 11450
rect 5912 11398 5942 11450
rect 5966 11398 5976 11450
rect 5976 11398 6022 11450
rect 6046 11398 6092 11450
rect 6092 11398 6102 11450
rect 6126 11398 6156 11450
rect 6156 11398 6182 11450
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 6126 11396 6182 11398
rect 6550 11328 6606 11384
rect 5630 11192 5632 11212
rect 5632 11192 5684 11212
rect 5684 11192 5686 11212
rect 5722 10376 5778 10432
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 6126 10362 6182 10364
rect 5886 10310 5912 10362
rect 5912 10310 5942 10362
rect 5966 10310 5976 10362
rect 5976 10310 6022 10362
rect 6046 10310 6092 10362
rect 6092 10310 6102 10362
rect 6126 10310 6156 10362
rect 6156 10310 6182 10362
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 6126 10308 6182 10310
rect 6366 9968 6422 10024
rect 5630 9832 5686 9888
rect 5446 9696 5502 9752
rect 5814 9460 5816 9480
rect 5816 9460 5868 9480
rect 5868 9460 5870 9480
rect 5814 9424 5870 9460
rect 5722 9288 5778 9344
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 6126 9274 6182 9276
rect 5886 9222 5912 9274
rect 5912 9222 5942 9274
rect 5966 9222 5976 9274
rect 5976 9222 6022 9274
rect 6046 9222 6092 9274
rect 6092 9222 6102 9274
rect 6126 9222 6156 9274
rect 6156 9222 6182 9274
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 6126 9220 6182 9222
rect 6458 8744 6514 8800
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 6126 8186 6182 8188
rect 5886 8134 5912 8186
rect 5912 8134 5942 8186
rect 5966 8134 5976 8186
rect 5976 8134 6022 8186
rect 6046 8134 6092 8186
rect 6092 8134 6102 8186
rect 6126 8134 6156 8186
rect 6156 8134 6182 8186
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 6126 8132 6182 8134
rect 6366 8064 6422 8120
rect 5722 7928 5778 7984
rect 5354 6704 5410 6760
rect 5170 6568 5226 6624
rect 5078 4120 5134 4176
rect 5078 3440 5134 3496
rect 5538 7520 5594 7576
rect 5722 7148 5724 7168
rect 5724 7148 5776 7168
rect 5776 7148 5778 7168
rect 5446 6568 5502 6624
rect 5722 7112 5778 7148
rect 6366 7112 6422 7168
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 6126 7098 6182 7100
rect 5886 7046 5912 7098
rect 5912 7046 5942 7098
rect 5966 7046 5976 7098
rect 5976 7046 6022 7098
rect 6046 7046 6092 7098
rect 6092 7046 6102 7098
rect 6126 7046 6156 7098
rect 6156 7046 6182 7098
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 6126 7044 6182 7046
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 5630 4276 5686 4312
rect 5630 4256 5632 4276
rect 5632 4256 5684 4276
rect 5684 4256 5686 4276
rect 5078 2796 5080 2816
rect 5080 2796 5132 2816
rect 5132 2796 5134 2816
rect 5078 2760 5134 2796
rect 5630 3712 5686 3768
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 7010 12416 7066 12472
rect 7102 10784 7158 10840
rect 7010 10376 7066 10432
rect 6642 10104 6698 10160
rect 7286 10668 7342 10704
rect 7286 10648 7288 10668
rect 7288 10648 7340 10668
rect 7340 10648 7342 10668
rect 6734 9968 6790 10024
rect 7194 9696 7250 9752
rect 7838 12960 7894 13016
rect 8390 13232 8446 13288
rect 8352 13082 8408 13084
rect 8432 13082 8488 13084
rect 8512 13082 8568 13084
rect 8592 13082 8648 13084
rect 8352 13030 8378 13082
rect 8378 13030 8408 13082
rect 8432 13030 8442 13082
rect 8442 13030 8488 13082
rect 8512 13030 8558 13082
rect 8558 13030 8568 13082
rect 8592 13030 8622 13082
rect 8622 13030 8648 13082
rect 8352 13028 8408 13030
rect 8432 13028 8488 13030
rect 8512 13028 8568 13030
rect 8592 13028 8648 13030
rect 8390 12164 8446 12200
rect 8390 12144 8392 12164
rect 8392 12144 8444 12164
rect 8444 12144 8446 12164
rect 8352 11994 8408 11996
rect 8432 11994 8488 11996
rect 8512 11994 8568 11996
rect 8592 11994 8648 11996
rect 8352 11942 8378 11994
rect 8378 11942 8408 11994
rect 8432 11942 8442 11994
rect 8442 11942 8488 11994
rect 8512 11942 8558 11994
rect 8558 11942 8568 11994
rect 8592 11942 8622 11994
rect 8622 11942 8648 11994
rect 8352 11940 8408 11942
rect 8432 11940 8488 11942
rect 8512 11940 8568 11942
rect 8592 11940 8648 11942
rect 8666 11464 8722 11520
rect 8352 10906 8408 10908
rect 8432 10906 8488 10908
rect 8512 10906 8568 10908
rect 8592 10906 8648 10908
rect 8352 10854 8378 10906
rect 8378 10854 8408 10906
rect 8432 10854 8442 10906
rect 8442 10854 8488 10906
rect 8512 10854 8558 10906
rect 8558 10854 8568 10906
rect 8592 10854 8622 10906
rect 8622 10854 8648 10906
rect 8352 10852 8408 10854
rect 8432 10852 8488 10854
rect 8512 10852 8568 10854
rect 8592 10852 8648 10854
rect 8022 9868 8024 9888
rect 8024 9868 8076 9888
rect 8076 9868 8078 9888
rect 8022 9832 8078 9868
rect 7654 9152 7710 9208
rect 6918 6024 6974 6080
rect 6826 3304 6882 3360
rect 7562 5616 7618 5672
rect 7470 4936 7526 4992
rect 7286 4256 7342 4312
rect 7562 3712 7618 3768
rect 8352 9818 8408 9820
rect 8432 9818 8488 9820
rect 8512 9818 8568 9820
rect 8592 9818 8648 9820
rect 8352 9766 8378 9818
rect 8378 9766 8408 9818
rect 8432 9766 8442 9818
rect 8442 9766 8488 9818
rect 8512 9766 8558 9818
rect 8558 9766 8568 9818
rect 8592 9766 8622 9818
rect 8622 9766 8648 9818
rect 8352 9764 8408 9766
rect 8432 9764 8488 9766
rect 8512 9764 8568 9766
rect 8592 9764 8648 9766
rect 8482 9424 8538 9480
rect 8758 9832 8814 9888
rect 8666 9152 8722 9208
rect 8352 8730 8408 8732
rect 8432 8730 8488 8732
rect 8512 8730 8568 8732
rect 8592 8730 8648 8732
rect 8352 8678 8378 8730
rect 8378 8678 8408 8730
rect 8432 8678 8442 8730
rect 8442 8678 8488 8730
rect 8512 8678 8558 8730
rect 8558 8678 8568 8730
rect 8592 8678 8622 8730
rect 8622 8678 8648 8730
rect 8352 8676 8408 8678
rect 8432 8676 8488 8678
rect 8512 8676 8568 8678
rect 8592 8676 8648 8678
rect 7838 6860 7894 6896
rect 7838 6840 7840 6860
rect 7840 6840 7892 6860
rect 7892 6840 7894 6860
rect 7746 5344 7802 5400
rect 7930 4120 7986 4176
rect 7654 3440 7710 3496
rect 7838 3168 7894 3224
rect 7562 2760 7618 2816
rect 7562 2488 7618 2544
rect 7838 2488 7894 2544
rect 8206 7656 8262 7712
rect 8352 7642 8408 7644
rect 8432 7642 8488 7644
rect 8512 7642 8568 7644
rect 8592 7642 8648 7644
rect 8352 7590 8378 7642
rect 8378 7590 8408 7642
rect 8432 7590 8442 7642
rect 8442 7590 8488 7642
rect 8512 7590 8558 7642
rect 8558 7590 8568 7642
rect 8592 7590 8622 7642
rect 8622 7590 8648 7642
rect 8352 7588 8408 7590
rect 8432 7588 8488 7590
rect 8512 7588 8568 7590
rect 8592 7588 8648 7590
rect 8114 7520 8170 7576
rect 8206 6604 8208 6624
rect 8208 6604 8260 6624
rect 8260 6604 8262 6624
rect 8206 6568 8262 6604
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 8114 6432 8170 6488
rect 8114 4392 8170 4448
rect 8022 3848 8078 3904
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 8666 4936 8722 4992
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 8022 2760 8078 2816
rect 8574 2760 8630 2816
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 9034 16360 9090 16416
rect 8942 15000 8998 15056
rect 9586 17448 9642 17504
rect 9126 15000 9182 15056
rect 9126 14728 9182 14784
rect 8942 12824 8998 12880
rect 8942 12552 8998 12608
rect 9218 14048 9274 14104
rect 9402 15680 9458 15736
rect 9034 10376 9090 10432
rect 9034 8608 9090 8664
rect 9034 8472 9090 8528
rect 9126 8236 9128 8256
rect 9128 8236 9180 8256
rect 9180 8236 9182 8256
rect 9126 8200 9182 8236
rect 9034 8064 9090 8120
rect 9586 16224 9642 16280
rect 9862 16360 9918 16416
rect 10138 17312 10194 17368
rect 9678 15272 9734 15328
rect 9678 15000 9734 15056
rect 9770 14728 9826 14784
rect 9770 14592 9826 14648
rect 9586 13096 9642 13152
rect 9586 12316 9588 12336
rect 9588 12316 9640 12336
rect 9640 12316 9642 12336
rect 9586 12280 9642 12316
rect 9586 11872 9642 11928
rect 9494 10240 9550 10296
rect 8942 3304 8998 3360
rect 9126 4120 9182 4176
rect 9494 9288 9550 9344
rect 10138 15000 10194 15056
rect 10138 14864 10194 14920
rect 9862 11192 9918 11248
rect 10322 15272 10378 15328
rect 10138 12180 10140 12200
rect 10140 12180 10192 12200
rect 10192 12180 10194 12200
rect 10138 12144 10194 12180
rect 10046 11464 10102 11520
rect 9954 10648 10010 10704
rect 9862 10240 9918 10296
rect 9770 9696 9826 9752
rect 9770 9288 9826 9344
rect 9586 8744 9642 8800
rect 9402 7928 9458 7984
rect 9586 7520 9642 7576
rect 9402 6432 9458 6488
rect 9402 6160 9458 6216
rect 9770 6840 9826 6896
rect 9310 5480 9366 5536
rect 9402 4936 9458 4992
rect 9402 4664 9458 4720
rect 9218 2760 9274 2816
rect 8942 2624 8998 2680
rect 10690 17312 10746 17368
rect 10598 16904 10654 16960
rect 10506 16768 10562 16824
rect 10506 16360 10562 16416
rect 10966 17176 11022 17232
rect 10817 16890 10873 16892
rect 10897 16890 10953 16892
rect 10977 16890 11033 16892
rect 11057 16890 11113 16892
rect 10817 16838 10843 16890
rect 10843 16838 10873 16890
rect 10897 16838 10907 16890
rect 10907 16838 10953 16890
rect 10977 16838 11023 16890
rect 11023 16838 11033 16890
rect 11057 16838 11087 16890
rect 11087 16838 11113 16890
rect 10817 16836 10873 16838
rect 10897 16836 10953 16838
rect 10977 16836 11033 16838
rect 11057 16836 11113 16838
rect 10817 15802 10873 15804
rect 10897 15802 10953 15804
rect 10977 15802 11033 15804
rect 11057 15802 11113 15804
rect 10817 15750 10843 15802
rect 10843 15750 10873 15802
rect 10897 15750 10907 15802
rect 10907 15750 10953 15802
rect 10977 15750 11023 15802
rect 11023 15750 11033 15802
rect 11057 15750 11087 15802
rect 11087 15750 11113 15802
rect 10817 15748 10873 15750
rect 10897 15748 10953 15750
rect 10977 15748 11033 15750
rect 11057 15748 11113 15750
rect 10506 15272 10562 15328
rect 10414 14456 10470 14512
rect 10506 14184 10562 14240
rect 10414 13640 10470 13696
rect 10414 12416 10470 12472
rect 10322 12008 10378 12064
rect 10138 9152 10194 9208
rect 10046 7384 10102 7440
rect 10046 7112 10102 7168
rect 10414 10648 10470 10704
rect 10690 15000 10746 15056
rect 10874 15000 10930 15056
rect 11150 14864 11206 14920
rect 10817 14714 10873 14716
rect 10897 14714 10953 14716
rect 10977 14714 11033 14716
rect 11057 14714 11113 14716
rect 10817 14662 10843 14714
rect 10843 14662 10873 14714
rect 10897 14662 10907 14714
rect 10907 14662 10953 14714
rect 10977 14662 11023 14714
rect 11023 14662 11033 14714
rect 11057 14662 11087 14714
rect 11087 14662 11113 14714
rect 10817 14660 10873 14662
rect 10897 14660 10953 14662
rect 10977 14660 11033 14662
rect 11057 14660 11113 14662
rect 10817 13626 10873 13628
rect 10897 13626 10953 13628
rect 10977 13626 11033 13628
rect 11057 13626 11113 13628
rect 10817 13574 10843 13626
rect 10843 13574 10873 13626
rect 10897 13574 10907 13626
rect 10907 13574 10953 13626
rect 10977 13574 11023 13626
rect 11023 13574 11033 13626
rect 11057 13574 11087 13626
rect 11087 13574 11113 13626
rect 10817 13572 10873 13574
rect 10897 13572 10953 13574
rect 10977 13572 11033 13574
rect 11057 13572 11113 13574
rect 11426 14592 11482 14648
rect 11334 14456 11390 14512
rect 11334 14340 11390 14376
rect 11334 14320 11336 14340
rect 11336 14320 11388 14340
rect 11388 14320 11390 14340
rect 11242 13232 11298 13288
rect 11150 13096 11206 13152
rect 10817 12538 10873 12540
rect 10897 12538 10953 12540
rect 10977 12538 11033 12540
rect 11057 12538 11113 12540
rect 10817 12486 10843 12538
rect 10843 12486 10873 12538
rect 10897 12486 10907 12538
rect 10907 12486 10953 12538
rect 10977 12486 11023 12538
rect 11023 12486 11033 12538
rect 11057 12486 11087 12538
rect 11087 12486 11113 12538
rect 10817 12484 10873 12486
rect 10897 12484 10953 12486
rect 10977 12484 11033 12486
rect 11057 12484 11113 12486
rect 10690 11736 10746 11792
rect 11150 11736 11206 11792
rect 10817 11450 10873 11452
rect 10897 11450 10953 11452
rect 10977 11450 11033 11452
rect 11057 11450 11113 11452
rect 10817 11398 10843 11450
rect 10843 11398 10873 11450
rect 10897 11398 10907 11450
rect 10907 11398 10953 11450
rect 10977 11398 11023 11450
rect 11023 11398 11033 11450
rect 11057 11398 11087 11450
rect 11087 11398 11113 11450
rect 10817 11396 10873 11398
rect 10897 11396 10953 11398
rect 10977 11396 11033 11398
rect 11057 11396 11113 11398
rect 11334 11736 11390 11792
rect 11150 10920 11206 10976
rect 10414 10240 10470 10296
rect 10506 9424 10562 9480
rect 10506 9324 10508 9344
rect 10508 9324 10560 9344
rect 10560 9324 10562 9344
rect 10506 9288 10562 9324
rect 10230 7656 10286 7712
rect 10414 7928 10470 7984
rect 10046 6568 10102 6624
rect 9770 6024 9826 6080
rect 10138 5752 10194 5808
rect 10322 7384 10378 7440
rect 10322 6976 10378 7032
rect 9770 5072 9826 5128
rect 9586 4392 9642 4448
rect 9954 4120 10010 4176
rect 9770 3712 9826 3768
rect 9954 2760 10010 2816
rect 9586 2624 9642 2680
rect 9862 2624 9918 2680
rect 9586 2352 9642 2408
rect 9586 2216 9642 2272
rect 10230 4800 10286 4856
rect 10322 4140 10378 4176
rect 10322 4120 10324 4140
rect 10324 4120 10376 4140
rect 10376 4120 10378 4140
rect 10414 3712 10470 3768
rect 10414 3576 10470 3632
rect 10414 3168 10470 3224
rect 11058 10512 11114 10568
rect 10817 10362 10873 10364
rect 10897 10362 10953 10364
rect 10977 10362 11033 10364
rect 11057 10362 11113 10364
rect 10817 10310 10843 10362
rect 10843 10310 10873 10362
rect 10897 10310 10907 10362
rect 10907 10310 10953 10362
rect 10977 10310 11023 10362
rect 11023 10310 11033 10362
rect 11057 10310 11087 10362
rect 11087 10310 11113 10362
rect 10817 10308 10873 10310
rect 10897 10308 10953 10310
rect 10977 10308 11033 10310
rect 11057 10308 11113 10310
rect 10782 9444 10838 9480
rect 10782 9424 10784 9444
rect 10784 9424 10836 9444
rect 10836 9424 10838 9444
rect 11242 10648 11298 10704
rect 11886 17448 11942 17504
rect 11610 13776 11666 13832
rect 11702 13096 11758 13152
rect 11610 12960 11666 13016
rect 11242 10512 11298 10568
rect 11978 12960 12034 13016
rect 11794 12824 11850 12880
rect 11702 12588 11704 12608
rect 11704 12588 11756 12608
rect 11756 12588 11758 12608
rect 11702 12552 11758 12588
rect 11702 12436 11758 12472
rect 11702 12416 11704 12436
rect 11704 12416 11756 12436
rect 11756 12416 11758 12436
rect 12162 16496 12218 16552
rect 12162 15544 12218 15600
rect 12162 15408 12218 15464
rect 12254 15156 12310 15192
rect 12254 15136 12256 15156
rect 12256 15136 12308 15156
rect 12308 15136 12310 15156
rect 11886 12416 11942 12472
rect 11334 9832 11390 9888
rect 11426 9460 11428 9480
rect 11428 9460 11480 9480
rect 11480 9460 11482 9480
rect 11426 9424 11482 9460
rect 10817 9274 10873 9276
rect 10897 9274 10953 9276
rect 10977 9274 11033 9276
rect 11057 9274 11113 9276
rect 10817 9222 10843 9274
rect 10843 9222 10873 9274
rect 10897 9222 10907 9274
rect 10907 9222 10953 9274
rect 10977 9222 11023 9274
rect 11023 9222 11033 9274
rect 11057 9222 11087 9274
rect 11087 9222 11113 9274
rect 10817 9220 10873 9222
rect 10897 9220 10953 9222
rect 10977 9220 11033 9222
rect 11057 9220 11113 9222
rect 10782 8744 10838 8800
rect 10817 8186 10873 8188
rect 10897 8186 10953 8188
rect 10977 8186 11033 8188
rect 11057 8186 11113 8188
rect 10817 8134 10843 8186
rect 10843 8134 10873 8186
rect 10897 8134 10907 8186
rect 10907 8134 10953 8186
rect 10977 8134 11023 8186
rect 11023 8134 11033 8186
rect 11057 8134 11087 8186
rect 11087 8134 11113 8186
rect 10817 8132 10873 8134
rect 10897 8132 10953 8134
rect 10977 8132 11033 8134
rect 11057 8132 11113 8134
rect 11702 9832 11758 9888
rect 11518 8064 11574 8120
rect 10874 7520 10930 7576
rect 11150 7520 11206 7576
rect 10817 7098 10873 7100
rect 10897 7098 10953 7100
rect 10977 7098 11033 7100
rect 11057 7098 11113 7100
rect 10817 7046 10843 7098
rect 10843 7046 10873 7098
rect 10897 7046 10907 7098
rect 10907 7046 10953 7098
rect 10977 7046 11023 7098
rect 11023 7046 11033 7098
rect 11057 7046 11087 7098
rect 11087 7046 11113 7098
rect 10817 7044 10873 7046
rect 10897 7044 10953 7046
rect 10977 7044 11033 7046
rect 11057 7044 11113 7046
rect 10966 6840 11022 6896
rect 11150 6840 11206 6896
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 10690 5072 10746 5128
rect 11242 5908 11298 5944
rect 11242 5888 11244 5908
rect 11244 5888 11296 5908
rect 11296 5888 11298 5908
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 11426 5344 11482 5400
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 11426 4392 11482 4448
rect 11334 4256 11390 4312
rect 11242 3848 11298 3904
rect 12070 11464 12126 11520
rect 11702 8064 11758 8120
rect 11794 7520 11850 7576
rect 12070 9832 12126 9888
rect 11978 8608 12034 8664
rect 12070 8064 12126 8120
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 11886 3984 11942 4040
rect 11518 2760 11574 2816
rect 10966 2216 11022 2272
rect 12254 12416 12310 12472
rect 12530 16496 12586 16552
rect 12622 15680 12678 15736
rect 12530 12008 12586 12064
rect 12438 11736 12494 11792
rect 12346 11600 12402 11656
rect 12438 11328 12494 11384
rect 12438 10920 12494 10976
rect 12438 10548 12440 10568
rect 12440 10548 12492 10568
rect 12492 10548 12494 10568
rect 12438 10512 12494 10548
rect 12438 9560 12494 9616
rect 12530 9424 12586 9480
rect 13282 17434 13338 17436
rect 13362 17434 13418 17436
rect 13442 17434 13498 17436
rect 13522 17434 13578 17436
rect 13282 17382 13308 17434
rect 13308 17382 13338 17434
rect 13362 17382 13372 17434
rect 13372 17382 13418 17434
rect 13442 17382 13488 17434
rect 13488 17382 13498 17434
rect 13522 17382 13552 17434
rect 13552 17382 13578 17434
rect 13282 17380 13338 17382
rect 13362 17380 13418 17382
rect 13442 17380 13498 17382
rect 13522 17380 13578 17382
rect 13358 17076 13360 17096
rect 13360 17076 13412 17096
rect 13412 17076 13414 17096
rect 13358 17040 13414 17076
rect 13174 16632 13230 16688
rect 13282 16346 13338 16348
rect 13362 16346 13418 16348
rect 13442 16346 13498 16348
rect 13522 16346 13578 16348
rect 13282 16294 13308 16346
rect 13308 16294 13338 16346
rect 13362 16294 13372 16346
rect 13372 16294 13418 16346
rect 13442 16294 13488 16346
rect 13488 16294 13498 16346
rect 13522 16294 13552 16346
rect 13552 16294 13578 16346
rect 13282 16292 13338 16294
rect 13362 16292 13418 16294
rect 13442 16292 13498 16294
rect 13522 16292 13578 16294
rect 13174 15544 13230 15600
rect 12714 11872 12770 11928
rect 13282 15258 13338 15260
rect 13362 15258 13418 15260
rect 13442 15258 13498 15260
rect 13522 15258 13578 15260
rect 13282 15206 13308 15258
rect 13308 15206 13338 15258
rect 13362 15206 13372 15258
rect 13372 15206 13418 15258
rect 13442 15206 13488 15258
rect 13488 15206 13498 15258
rect 13522 15206 13552 15258
rect 13552 15206 13578 15258
rect 13282 15204 13338 15206
rect 13362 15204 13418 15206
rect 13442 15204 13498 15206
rect 13522 15204 13578 15206
rect 13282 14170 13338 14172
rect 13362 14170 13418 14172
rect 13442 14170 13498 14172
rect 13522 14170 13578 14172
rect 13282 14118 13308 14170
rect 13308 14118 13338 14170
rect 13362 14118 13372 14170
rect 13372 14118 13418 14170
rect 13442 14118 13488 14170
rect 13488 14118 13498 14170
rect 13522 14118 13552 14170
rect 13552 14118 13578 14170
rect 13282 14116 13338 14118
rect 13362 14116 13418 14118
rect 13442 14116 13498 14118
rect 13522 14116 13578 14118
rect 12530 8744 12586 8800
rect 12530 8336 12586 8392
rect 12438 7520 12494 7576
rect 12622 8064 12678 8120
rect 12898 9152 12954 9208
rect 12806 8472 12862 8528
rect 12898 7520 12954 7576
rect 12806 7148 12808 7168
rect 12808 7148 12860 7168
rect 12860 7148 12862 7168
rect 12806 7112 12862 7148
rect 12438 6160 12494 6216
rect 12806 5616 12862 5672
rect 12714 5480 12770 5536
rect 13282 13082 13338 13084
rect 13362 13082 13418 13084
rect 13442 13082 13498 13084
rect 13522 13082 13578 13084
rect 13282 13030 13308 13082
rect 13308 13030 13338 13082
rect 13362 13030 13372 13082
rect 13372 13030 13418 13082
rect 13442 13030 13488 13082
rect 13488 13030 13498 13082
rect 13522 13030 13552 13082
rect 13552 13030 13578 13082
rect 13282 13028 13338 13030
rect 13362 13028 13418 13030
rect 13442 13028 13498 13030
rect 13522 13028 13578 13030
rect 13450 12824 13506 12880
rect 13910 15952 13966 16008
rect 13818 13912 13874 13968
rect 13726 13504 13782 13560
rect 13726 13368 13782 13424
rect 13726 13096 13782 13152
rect 13282 11994 13338 11996
rect 13362 11994 13418 11996
rect 13442 11994 13498 11996
rect 13522 11994 13578 11996
rect 13282 11942 13308 11994
rect 13308 11942 13338 11994
rect 13362 11942 13372 11994
rect 13372 11942 13418 11994
rect 13442 11942 13488 11994
rect 13488 11942 13498 11994
rect 13522 11942 13552 11994
rect 13552 11942 13578 11994
rect 13282 11940 13338 11942
rect 13362 11940 13418 11942
rect 13442 11940 13498 11942
rect 13522 11940 13578 11942
rect 13082 11056 13138 11112
rect 13282 10906 13338 10908
rect 13362 10906 13418 10908
rect 13442 10906 13498 10908
rect 13522 10906 13578 10908
rect 13282 10854 13308 10906
rect 13308 10854 13338 10906
rect 13362 10854 13372 10906
rect 13372 10854 13418 10906
rect 13442 10854 13488 10906
rect 13488 10854 13498 10906
rect 13522 10854 13552 10906
rect 13552 10854 13578 10906
rect 13282 10852 13338 10854
rect 13362 10852 13418 10854
rect 13442 10852 13498 10854
rect 13522 10852 13578 10854
rect 13450 10376 13506 10432
rect 13358 10124 13414 10160
rect 13358 10104 13360 10124
rect 13360 10104 13412 10124
rect 13412 10104 13414 10124
rect 13726 10124 13782 10160
rect 13726 10104 13728 10124
rect 13728 10104 13780 10124
rect 13780 10104 13782 10124
rect 13282 9818 13338 9820
rect 13362 9818 13418 9820
rect 13442 9818 13498 9820
rect 13522 9818 13578 9820
rect 13282 9766 13308 9818
rect 13308 9766 13338 9818
rect 13362 9766 13372 9818
rect 13372 9766 13418 9818
rect 13442 9766 13488 9818
rect 13488 9766 13498 9818
rect 13522 9766 13552 9818
rect 13552 9766 13578 9818
rect 13282 9764 13338 9766
rect 13362 9764 13418 9766
rect 13442 9764 13498 9766
rect 13522 9764 13578 9766
rect 13174 9324 13176 9344
rect 13176 9324 13228 9344
rect 13228 9324 13230 9344
rect 13174 9288 13230 9324
rect 13174 9172 13230 9208
rect 13174 9152 13176 9172
rect 13176 9152 13228 9172
rect 13228 9152 13230 9172
rect 13266 9016 13322 9072
rect 12346 3984 12402 4040
rect 12438 3304 12494 3360
rect 12346 3168 12402 3224
rect 12622 3168 12678 3224
rect 12530 2624 12586 2680
rect 12530 2488 12586 2544
rect 13282 8730 13338 8732
rect 13362 8730 13418 8732
rect 13442 8730 13498 8732
rect 13522 8730 13578 8732
rect 13282 8678 13308 8730
rect 13308 8678 13338 8730
rect 13362 8678 13372 8730
rect 13372 8678 13418 8730
rect 13442 8678 13488 8730
rect 13488 8678 13498 8730
rect 13522 8678 13552 8730
rect 13552 8678 13578 8730
rect 13282 8676 13338 8678
rect 13362 8676 13418 8678
rect 13442 8676 13498 8678
rect 13522 8676 13578 8678
rect 13174 8200 13230 8256
rect 13266 7812 13322 7848
rect 13266 7792 13268 7812
rect 13268 7792 13320 7812
rect 13320 7792 13322 7812
rect 13282 7642 13338 7644
rect 13362 7642 13418 7644
rect 13442 7642 13498 7644
rect 13522 7642 13578 7644
rect 13282 7590 13308 7642
rect 13308 7590 13338 7642
rect 13362 7590 13372 7642
rect 13372 7590 13418 7642
rect 13442 7590 13488 7642
rect 13488 7590 13498 7642
rect 13522 7590 13552 7642
rect 13552 7590 13578 7642
rect 13282 7588 13338 7590
rect 13362 7588 13418 7590
rect 13442 7588 13498 7590
rect 13522 7588 13578 7590
rect 14186 16088 14242 16144
rect 13910 9424 13966 9480
rect 13634 7248 13690 7304
rect 13910 8608 13966 8664
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 13450 6332 13452 6352
rect 13452 6332 13504 6352
rect 13504 6332 13506 6352
rect 13450 6296 13506 6332
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 13450 5208 13506 5264
rect 13358 4684 13414 4720
rect 13358 4664 13360 4684
rect 13360 4664 13412 4684
rect 13412 4664 13414 4684
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 13358 4120 13414 4176
rect 13266 3848 13322 3904
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 12990 2624 13046 2680
rect 13818 6840 13874 6896
rect 13818 5752 13874 5808
rect 14002 4528 14058 4584
rect 14646 17584 14702 17640
rect 14830 12724 14832 12744
rect 14832 12724 14884 12744
rect 14884 12724 14886 12744
rect 14830 12688 14886 12724
rect 14646 9988 14702 10024
rect 14646 9968 14648 9988
rect 14648 9968 14700 9988
rect 14700 9968 14702 9988
rect 14554 7928 14610 7984
rect 14646 7384 14702 7440
rect 14186 5616 14242 5672
rect 13910 2760 13966 2816
rect 13266 2352 13322 2408
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
rect 14462 5072 14518 5128
rect 14554 3984 14610 4040
rect 14462 3848 14518 3904
rect 14646 3576 14702 3632
rect 14646 3460 14702 3496
rect 14646 3440 14648 3460
rect 14648 3440 14700 3460
rect 14700 3440 14702 3460
rect 15014 10240 15070 10296
rect 14922 9968 14978 10024
rect 15014 8880 15070 8936
rect 15014 6704 15070 6760
rect 15014 4156 15016 4176
rect 15016 4156 15068 4176
rect 15068 4156 15070 4176
rect 15014 4120 15070 4156
rect 15014 3068 15016 3088
rect 15016 3068 15068 3088
rect 15068 3068 15070 3088
rect 15014 3032 15070 3068
rect 16026 17584 16082 17640
rect 15566 6024 15622 6080
rect 16762 2896 16818 2952
<< metal3 >>
rect 0 19410 480 19440
rect 1485 19410 1551 19413
rect 0 19408 1551 19410
rect 0 19352 1490 19408
rect 1546 19352 1551 19408
rect 0 19350 1551 19352
rect 0 19320 480 19350
rect 1485 19347 1551 19350
rect 0 18458 480 18488
rect 1669 18458 1735 18461
rect 0 18456 1735 18458
rect 0 18400 1674 18456
rect 1730 18400 1735 18456
rect 0 18398 1735 18400
rect 0 18368 480 18398
rect 1669 18395 1735 18398
rect 8937 17642 9003 17645
rect 14641 17642 14707 17645
rect 16021 17642 16087 17645
rect 8937 17640 16087 17642
rect 8937 17584 8942 17640
rect 8998 17584 14646 17640
rect 14702 17584 16026 17640
rect 16082 17584 16087 17640
rect 8937 17582 16087 17584
rect 8937 17579 9003 17582
rect 14641 17579 14707 17582
rect 16021 17579 16087 17582
rect 9581 17506 9647 17509
rect 11881 17506 11947 17509
rect 9581 17504 11947 17506
rect 9581 17448 9586 17504
rect 9642 17448 11886 17504
rect 11942 17448 11947 17504
rect 9581 17446 11947 17448
rect 9581 17443 9647 17446
rect 11881 17443 11947 17446
rect 3409 17440 3729 17441
rect 0 17370 480 17400
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 17375 3729 17376
rect 8340 17440 8660 17441
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 17375 8660 17376
rect 13270 17440 13590 17441
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 13270 17375 13590 17376
rect 2957 17370 3023 17373
rect 0 17368 3023 17370
rect 0 17312 2962 17368
rect 3018 17312 3023 17368
rect 0 17310 3023 17312
rect 0 17280 480 17310
rect 2957 17307 3023 17310
rect 10133 17370 10199 17373
rect 10685 17370 10751 17373
rect 10133 17368 10751 17370
rect 10133 17312 10138 17368
rect 10194 17312 10690 17368
rect 10746 17312 10751 17368
rect 10133 17310 10751 17312
rect 10133 17307 10199 17310
rect 10685 17307 10751 17310
rect 9622 17172 9628 17236
rect 9692 17234 9698 17236
rect 10961 17234 11027 17237
rect 9692 17232 11027 17234
rect 9692 17176 10966 17232
rect 11022 17176 11027 17232
rect 9692 17174 11027 17176
rect 9692 17172 9698 17174
rect 10961 17171 11027 17174
rect 10174 17036 10180 17100
rect 10244 17098 10250 17100
rect 13353 17098 13419 17101
rect 10244 17096 13419 17098
rect 10244 17040 13358 17096
rect 13414 17040 13419 17096
rect 10244 17038 13419 17040
rect 10244 17036 10250 17038
rect 13353 17035 13419 17038
rect 3182 16900 3188 16964
rect 3252 16962 3258 16964
rect 3325 16962 3391 16965
rect 3252 16960 3391 16962
rect 3252 16904 3330 16960
rect 3386 16904 3391 16960
rect 3252 16902 3391 16904
rect 3252 16900 3258 16902
rect 3325 16899 3391 16902
rect 7649 16962 7715 16965
rect 10593 16962 10659 16965
rect 7649 16960 10659 16962
rect 7649 16904 7654 16960
rect 7710 16904 10598 16960
rect 10654 16904 10659 16960
rect 7649 16902 10659 16904
rect 7649 16899 7715 16902
rect 10593 16899 10659 16902
rect 5874 16896 6194 16897
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6194 16896
rect 5874 16831 6194 16832
rect 10805 16896 11125 16897
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 16831 11125 16832
rect 8569 16826 8635 16829
rect 9806 16826 9812 16828
rect 8569 16824 9812 16826
rect 8569 16768 8574 16824
rect 8630 16768 9812 16824
rect 8569 16766 9812 16768
rect 8569 16763 8635 16766
rect 9806 16764 9812 16766
rect 9876 16826 9882 16828
rect 10501 16826 10567 16829
rect 9876 16824 10567 16826
rect 9876 16768 10506 16824
rect 10562 16768 10567 16824
rect 9876 16766 10567 16768
rect 9876 16764 9882 16766
rect 10501 16763 10567 16766
rect 4981 16690 5047 16693
rect 10358 16690 10364 16692
rect 4981 16688 10364 16690
rect 4981 16632 4986 16688
rect 5042 16632 10364 16688
rect 4981 16630 10364 16632
rect 4981 16627 5047 16630
rect 10358 16628 10364 16630
rect 10428 16628 10434 16692
rect 13169 16690 13235 16693
rect 13670 16690 13676 16692
rect 13169 16688 13676 16690
rect 13169 16632 13174 16688
rect 13230 16632 13676 16688
rect 13169 16630 13676 16632
rect 13169 16627 13235 16630
rect 13670 16628 13676 16630
rect 13740 16690 13746 16692
rect 16520 16690 17000 16720
rect 13740 16630 17000 16690
rect 13740 16628 13746 16630
rect 16520 16600 17000 16630
rect 5809 16554 5875 16557
rect 12157 16554 12223 16557
rect 12525 16556 12591 16557
rect 12525 16554 12572 16556
rect 5809 16552 12223 16554
rect 5809 16496 5814 16552
rect 5870 16496 12162 16552
rect 12218 16496 12223 16552
rect 5809 16494 12223 16496
rect 12480 16552 12572 16554
rect 12480 16496 12530 16552
rect 12480 16494 12572 16496
rect 5809 16491 5875 16494
rect 12157 16491 12223 16494
rect 12525 16492 12572 16494
rect 12636 16492 12642 16556
rect 12525 16491 12591 16492
rect 0 16418 480 16448
rect 2865 16418 2931 16421
rect 0 16416 2931 16418
rect 0 16360 2870 16416
rect 2926 16360 2931 16416
rect 0 16358 2931 16360
rect 0 16328 480 16358
rect 2865 16355 2931 16358
rect 9029 16418 9095 16421
rect 9857 16418 9923 16421
rect 9029 16416 9923 16418
rect 9029 16360 9034 16416
rect 9090 16360 9862 16416
rect 9918 16360 9923 16416
rect 9029 16358 9923 16360
rect 9029 16355 9095 16358
rect 9857 16355 9923 16358
rect 9990 16356 9996 16420
rect 10060 16418 10066 16420
rect 10501 16418 10567 16421
rect 10060 16416 10567 16418
rect 10060 16360 10506 16416
rect 10562 16360 10567 16416
rect 10060 16358 10567 16360
rect 10060 16356 10066 16358
rect 10501 16355 10567 16358
rect 3409 16352 3729 16353
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 16287 3729 16288
rect 8340 16352 8660 16353
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 16287 8660 16288
rect 13270 16352 13590 16353
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 16287 13590 16288
rect 9581 16282 9647 16285
rect 12566 16282 12572 16284
rect 9581 16280 12572 16282
rect 9581 16224 9586 16280
rect 9642 16224 12572 16280
rect 9581 16222 12572 16224
rect 9581 16219 9647 16222
rect 12566 16220 12572 16222
rect 12636 16220 12642 16284
rect 8109 16146 8175 16149
rect 14181 16146 14247 16149
rect 8109 16144 14247 16146
rect 8109 16088 8114 16144
rect 8170 16088 14186 16144
rect 14242 16088 14247 16144
rect 8109 16086 14247 16088
rect 8109 16083 8175 16086
rect 14181 16083 14247 16086
rect 4337 16010 4403 16013
rect 13905 16010 13971 16013
rect 4337 16008 13971 16010
rect 4337 15952 4342 16008
rect 4398 15952 13910 16008
rect 13966 15952 13971 16008
rect 4337 15950 13971 15952
rect 4337 15947 4403 15950
rect 13905 15947 13971 15950
rect 5874 15808 6194 15809
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6194 15808
rect 5874 15743 6194 15744
rect 10805 15808 11125 15809
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 15743 11125 15744
rect 9397 15740 9463 15741
rect 9397 15738 9444 15740
rect 6318 15736 9444 15738
rect 9508 15738 9514 15740
rect 6318 15680 9402 15736
rect 6318 15678 9444 15680
rect 5441 15602 5507 15605
rect 6318 15602 6378 15678
rect 9397 15676 9444 15678
rect 9508 15678 9590 15738
rect 9508 15676 9514 15678
rect 12198 15676 12204 15740
rect 12268 15738 12274 15740
rect 12617 15738 12683 15741
rect 12268 15736 12683 15738
rect 12268 15680 12622 15736
rect 12678 15680 12683 15736
rect 12268 15678 12683 15680
rect 12268 15676 12274 15678
rect 9397 15675 9463 15676
rect 12617 15675 12683 15678
rect 5441 15600 6378 15602
rect 5441 15544 5446 15600
rect 5502 15544 6378 15600
rect 5441 15542 6378 15544
rect 6545 15602 6611 15605
rect 12157 15602 12223 15605
rect 6545 15600 12223 15602
rect 6545 15544 6550 15600
rect 6606 15544 12162 15600
rect 12218 15544 12223 15600
rect 6545 15542 12223 15544
rect 5441 15539 5507 15542
rect 6545 15539 6611 15542
rect 12157 15539 12223 15542
rect 12382 15540 12388 15604
rect 12452 15602 12458 15604
rect 13169 15602 13235 15605
rect 12452 15600 13235 15602
rect 12452 15544 13174 15600
rect 13230 15544 13235 15600
rect 12452 15542 13235 15544
rect 12452 15540 12458 15542
rect 13169 15539 13235 15542
rect 0 15466 480 15496
rect 3601 15466 3667 15469
rect 0 15464 3667 15466
rect 0 15408 3606 15464
rect 3662 15408 3667 15464
rect 0 15406 3667 15408
rect 0 15376 480 15406
rect 3601 15403 3667 15406
rect 4613 15466 4679 15469
rect 6545 15466 6611 15469
rect 4613 15464 6611 15466
rect 4613 15408 4618 15464
rect 4674 15408 6550 15464
rect 6606 15408 6611 15464
rect 4613 15406 6611 15408
rect 4613 15403 4679 15406
rect 6545 15403 6611 15406
rect 8109 15466 8175 15469
rect 12157 15466 12223 15469
rect 8109 15464 12223 15466
rect 8109 15408 8114 15464
rect 8170 15408 12162 15464
rect 12218 15408 12223 15464
rect 8109 15406 12223 15408
rect 8109 15403 8175 15406
rect 12157 15403 12223 15406
rect 9673 15330 9739 15333
rect 10317 15330 10383 15333
rect 10501 15332 10567 15333
rect 10501 15330 10548 15332
rect 9673 15328 10383 15330
rect 9673 15272 9678 15328
rect 9734 15272 10322 15328
rect 10378 15272 10383 15328
rect 9673 15270 10383 15272
rect 10456 15328 10548 15330
rect 10456 15272 10506 15328
rect 10456 15270 10548 15272
rect 9673 15267 9739 15270
rect 10317 15267 10383 15270
rect 10501 15268 10548 15270
rect 10612 15268 10618 15332
rect 10501 15267 10567 15268
rect 3409 15264 3729 15265
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 15199 3729 15200
rect 8340 15264 8660 15265
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 15199 8660 15200
rect 13270 15264 13590 15265
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 15199 13590 15200
rect 9254 15132 9260 15196
rect 9324 15194 9330 15196
rect 12249 15194 12315 15197
rect 9324 15192 12315 15194
rect 9324 15136 12254 15192
rect 12310 15136 12315 15192
rect 9324 15134 12315 15136
rect 9324 15132 9330 15134
rect 12249 15131 12315 15134
rect 4337 15058 4403 15061
rect 8937 15058 9003 15061
rect 4337 15056 9003 15058
rect 4337 15000 4342 15056
rect 4398 15000 8942 15056
rect 8998 15000 9003 15056
rect 4337 14998 9003 15000
rect 4337 14995 4403 14998
rect 8937 14995 9003 14998
rect 9121 15058 9187 15061
rect 9673 15058 9739 15061
rect 9121 15056 9739 15058
rect 9121 15000 9126 15056
rect 9182 15000 9678 15056
rect 9734 15000 9739 15056
rect 9121 14998 9739 15000
rect 9121 14995 9187 14998
rect 9673 14995 9739 14998
rect 10133 15058 10199 15061
rect 10685 15058 10751 15061
rect 10133 15056 10751 15058
rect 10133 15000 10138 15056
rect 10194 15000 10690 15056
rect 10746 15000 10751 15056
rect 10133 14998 10751 15000
rect 10133 14995 10199 14998
rect 10685 14995 10751 14998
rect 10869 15058 10935 15061
rect 12750 15058 12756 15060
rect 10869 15056 12756 15058
rect 10869 15000 10874 15056
rect 10930 15000 12756 15056
rect 10869 14998 12756 15000
rect 10869 14995 10935 14998
rect 12750 14996 12756 14998
rect 12820 14996 12826 15060
rect 5717 14922 5783 14925
rect 10133 14922 10199 14925
rect 11145 14922 11211 14925
rect 5717 14920 10199 14922
rect 5717 14864 5722 14920
rect 5778 14864 10138 14920
rect 10194 14864 10199 14920
rect 5717 14862 10199 14864
rect 5717 14859 5783 14862
rect 10133 14859 10199 14862
rect 10320 14920 11211 14922
rect 10320 14864 11150 14920
rect 11206 14864 11211 14920
rect 10320 14862 11211 14864
rect 7281 14786 7347 14789
rect 9121 14786 9187 14789
rect 7281 14784 9187 14786
rect 7281 14728 7286 14784
rect 7342 14728 9126 14784
rect 9182 14728 9187 14784
rect 7281 14726 9187 14728
rect 7281 14723 7347 14726
rect 9121 14723 9187 14726
rect 9765 14786 9831 14789
rect 10320 14786 10380 14862
rect 11145 14859 11211 14862
rect 9765 14784 10380 14786
rect 9765 14728 9770 14784
rect 9826 14728 10380 14784
rect 9765 14726 10380 14728
rect 9765 14723 9831 14726
rect 5874 14720 6194 14721
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6194 14720
rect 5874 14655 6194 14656
rect 10805 14720 11125 14721
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 14655 11125 14656
rect 8661 14650 8727 14653
rect 8886 14650 8892 14652
rect 8661 14648 8892 14650
rect 8661 14592 8666 14648
rect 8722 14592 8892 14648
rect 8661 14590 8892 14592
rect 8661 14587 8727 14590
rect 8886 14588 8892 14590
rect 8956 14588 8962 14652
rect 9622 14588 9628 14652
rect 9692 14650 9698 14652
rect 9765 14650 9831 14653
rect 9692 14648 9831 14650
rect 9692 14592 9770 14648
rect 9826 14592 9831 14648
rect 9692 14590 9831 14592
rect 9692 14588 9698 14590
rect 9765 14587 9831 14590
rect 11421 14650 11487 14653
rect 12934 14650 12940 14652
rect 11421 14648 12940 14650
rect 11421 14592 11426 14648
rect 11482 14592 12940 14648
rect 11421 14590 12940 14592
rect 11421 14587 11487 14590
rect 12934 14588 12940 14590
rect 13004 14588 13010 14652
rect 2773 14514 2839 14517
rect 9070 14514 9076 14516
rect 2773 14512 9076 14514
rect 2773 14456 2778 14512
rect 2834 14456 9076 14512
rect 2773 14454 9076 14456
rect 2773 14451 2839 14454
rect 9070 14452 9076 14454
rect 9140 14452 9146 14516
rect 9622 14452 9628 14516
rect 9692 14514 9698 14516
rect 10409 14514 10475 14517
rect 11329 14516 11395 14517
rect 11278 14514 11284 14516
rect 9692 14512 10475 14514
rect 9692 14456 10414 14512
rect 10470 14456 10475 14512
rect 9692 14454 10475 14456
rect 11238 14454 11284 14514
rect 11348 14512 11395 14516
rect 11390 14456 11395 14512
rect 9692 14452 9698 14454
rect 10409 14451 10475 14454
rect 11278 14452 11284 14454
rect 11348 14452 11395 14456
rect 11329 14451 11395 14452
rect 0 14378 480 14408
rect 4061 14378 4127 14381
rect 0 14376 4127 14378
rect 0 14320 4066 14376
rect 4122 14320 4127 14376
rect 0 14318 4127 14320
rect 0 14288 480 14318
rect 4061 14315 4127 14318
rect 4889 14378 4955 14381
rect 11329 14378 11395 14381
rect 4889 14376 11395 14378
rect 4889 14320 4894 14376
rect 4950 14320 11334 14376
rect 11390 14320 11395 14376
rect 4889 14318 11395 14320
rect 4889 14315 4955 14318
rect 11329 14315 11395 14318
rect 10501 14242 10567 14245
rect 11462 14242 11468 14244
rect 10501 14240 11468 14242
rect 10501 14184 10506 14240
rect 10562 14184 11468 14240
rect 10501 14182 11468 14184
rect 10501 14179 10567 14182
rect 11462 14180 11468 14182
rect 11532 14180 11538 14244
rect 3409 14176 3729 14177
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 14111 3729 14112
rect 8340 14176 8660 14177
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 14111 8660 14112
rect 13270 14176 13590 14177
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 14111 13590 14112
rect 9070 14044 9076 14108
rect 9140 14106 9146 14108
rect 9213 14106 9279 14109
rect 12014 14106 12020 14108
rect 9140 14104 12020 14106
rect 9140 14048 9218 14104
rect 9274 14048 12020 14104
rect 9140 14046 12020 14048
rect 9140 14044 9146 14046
rect 9213 14043 9279 14046
rect 12014 14044 12020 14046
rect 12084 14044 12090 14108
rect 2405 13970 2471 13973
rect 13813 13970 13879 13973
rect 2405 13968 13879 13970
rect 2405 13912 2410 13968
rect 2466 13912 13818 13968
rect 13874 13912 13879 13968
rect 2405 13910 13879 13912
rect 2405 13907 2471 13910
rect 13813 13907 13879 13910
rect 2865 13834 2931 13837
rect 11605 13834 11671 13837
rect 2865 13832 11671 13834
rect 2865 13776 2870 13832
rect 2926 13776 11610 13832
rect 11666 13776 11671 13832
rect 2865 13774 11671 13776
rect 2865 13771 2931 13774
rect 11605 13771 11671 13774
rect 7741 13698 7807 13701
rect 9438 13698 9444 13700
rect 7741 13696 9444 13698
rect 7741 13640 7746 13696
rect 7802 13640 9444 13696
rect 7741 13638 9444 13640
rect 7741 13635 7807 13638
rect 9438 13636 9444 13638
rect 9508 13698 9514 13700
rect 10409 13698 10475 13701
rect 9508 13696 10475 13698
rect 9508 13640 10414 13696
rect 10470 13640 10475 13696
rect 9508 13638 10475 13640
rect 9508 13636 9514 13638
rect 10409 13635 10475 13638
rect 5874 13632 6194 13633
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6194 13632
rect 5874 13567 6194 13568
rect 10805 13632 11125 13633
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 13567 11125 13568
rect 4061 13562 4127 13565
rect 5717 13562 5783 13565
rect 4061 13560 5783 13562
rect 4061 13504 4066 13560
rect 4122 13504 5722 13560
rect 5778 13504 5783 13560
rect 4061 13502 5783 13504
rect 4061 13499 4127 13502
rect 5717 13499 5783 13502
rect 7097 13562 7163 13565
rect 9254 13562 9260 13564
rect 7097 13560 9260 13562
rect 7097 13504 7102 13560
rect 7158 13504 9260 13560
rect 7097 13502 9260 13504
rect 7097 13499 7163 13502
rect 9254 13500 9260 13502
rect 9324 13500 9330 13564
rect 9438 13500 9444 13564
rect 9508 13562 9514 13564
rect 9990 13562 9996 13564
rect 9508 13502 9996 13562
rect 9508 13500 9514 13502
rect 9990 13500 9996 13502
rect 10060 13500 10066 13564
rect 11646 13500 11652 13564
rect 11716 13562 11722 13564
rect 13721 13562 13787 13565
rect 11716 13560 13787 13562
rect 11716 13504 13726 13560
rect 13782 13504 13787 13560
rect 11716 13502 13787 13504
rect 11716 13500 11722 13502
rect 13721 13499 13787 13502
rect 0 13426 480 13456
rect 13721 13426 13787 13429
rect 0 13424 13787 13426
rect 0 13368 13726 13424
rect 13782 13368 13787 13424
rect 0 13366 13787 13368
rect 0 13336 480 13366
rect 13721 13363 13787 13366
rect 8385 13290 8451 13293
rect 9070 13290 9076 13292
rect 8385 13288 9076 13290
rect 8385 13232 8390 13288
rect 8446 13232 9076 13288
rect 8385 13230 9076 13232
rect 8385 13227 8451 13230
rect 9070 13228 9076 13230
rect 9140 13290 9146 13292
rect 11237 13290 11303 13293
rect 9140 13288 11303 13290
rect 9140 13232 11242 13288
rect 11298 13232 11303 13288
rect 9140 13230 11303 13232
rect 9140 13228 9146 13230
rect 11237 13227 11303 13230
rect 4337 13154 4403 13157
rect 7005 13154 7071 13157
rect 9581 13154 9647 13157
rect 11145 13154 11211 13157
rect 11697 13154 11763 13157
rect 13721 13156 13787 13157
rect 4337 13152 7071 13154
rect 4337 13096 4342 13152
rect 4398 13096 7010 13152
rect 7066 13096 7071 13152
rect 4337 13094 7071 13096
rect 4337 13091 4403 13094
rect 7005 13091 7071 13094
rect 8756 13152 11763 13154
rect 8756 13096 9586 13152
rect 9642 13096 11150 13152
rect 11206 13096 11702 13152
rect 11758 13096 11763 13152
rect 8756 13094 11763 13096
rect 3409 13088 3729 13089
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 13023 3729 13024
rect 8340 13088 8660 13089
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 13023 8660 13024
rect 6913 13018 6979 13021
rect 7833 13018 7899 13021
rect 6548 13016 7899 13018
rect 6548 12960 6918 13016
rect 6974 12960 7838 13016
rect 7894 12960 7899 13016
rect 6548 12958 7899 12960
rect 2497 12882 2563 12885
rect 6548 12882 6608 12958
rect 6913 12955 6979 12958
rect 7833 12955 7899 12958
rect 2497 12880 6608 12882
rect 2497 12824 2502 12880
rect 2558 12824 6608 12880
rect 2497 12822 6608 12824
rect 2497 12819 2563 12822
rect 6678 12820 6684 12884
rect 6748 12882 6754 12884
rect 8756 12882 8816 13094
rect 9581 13091 9647 13094
rect 11145 13091 11211 13094
rect 11697 13091 11763 13094
rect 13670 13092 13676 13156
rect 13740 13154 13787 13156
rect 13740 13152 13832 13154
rect 13782 13096 13832 13152
rect 13740 13094 13832 13096
rect 13740 13092 13787 13094
rect 13721 13091 13787 13092
rect 13270 13088 13590 13089
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 13023 13590 13024
rect 11605 13018 11671 13021
rect 11973 13018 12039 13021
rect 11605 13016 12039 13018
rect 11605 12960 11610 13016
rect 11666 12960 11978 13016
rect 12034 12960 12039 13016
rect 11605 12958 12039 12960
rect 11605 12955 11671 12958
rect 11973 12955 12039 12958
rect 6748 12822 8816 12882
rect 8937 12882 9003 12885
rect 11789 12884 11855 12885
rect 10174 12882 10180 12884
rect 8937 12880 10180 12882
rect 8937 12824 8942 12880
rect 8998 12824 10180 12880
rect 8937 12822 10180 12824
rect 6748 12820 6754 12822
rect 8937 12819 9003 12822
rect 10174 12820 10180 12822
rect 10244 12820 10250 12884
rect 11789 12882 11836 12884
rect 11744 12880 11836 12882
rect 11744 12824 11794 12880
rect 11744 12822 11836 12824
rect 11789 12820 11836 12822
rect 11900 12820 11906 12884
rect 12014 12820 12020 12884
rect 12084 12882 12090 12884
rect 13445 12882 13511 12885
rect 12084 12880 13511 12882
rect 12084 12824 13450 12880
rect 13506 12824 13511 12880
rect 12084 12822 13511 12824
rect 12084 12820 12090 12822
rect 11789 12819 11855 12820
rect 13445 12819 13511 12822
rect 2589 12746 2655 12749
rect 6177 12746 6243 12749
rect 2589 12744 6243 12746
rect 2589 12688 2594 12744
rect 2650 12688 6182 12744
rect 6238 12688 6243 12744
rect 2589 12686 6243 12688
rect 2589 12683 2655 12686
rect 6177 12683 6243 12686
rect 6729 12746 6795 12749
rect 14825 12746 14891 12749
rect 6729 12744 14891 12746
rect 6729 12688 6734 12744
rect 6790 12688 14830 12744
rect 14886 12688 14891 12744
rect 6729 12686 14891 12688
rect 6729 12683 6795 12686
rect 14825 12683 14891 12686
rect 6453 12610 6519 12613
rect 8937 12610 9003 12613
rect 6453 12608 9003 12610
rect 6453 12552 6458 12608
rect 6514 12552 8942 12608
rect 8998 12552 9003 12608
rect 6453 12550 9003 12552
rect 6453 12547 6519 12550
rect 8937 12547 9003 12550
rect 11697 12610 11763 12613
rect 12014 12610 12020 12612
rect 11697 12608 12020 12610
rect 11697 12552 11702 12608
rect 11758 12552 12020 12608
rect 11697 12550 12020 12552
rect 11697 12547 11763 12550
rect 12014 12548 12020 12550
rect 12084 12548 12090 12612
rect 5874 12544 6194 12545
rect 0 12474 480 12504
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6194 12544
rect 5874 12479 6194 12480
rect 10805 12544 11125 12545
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 12479 11125 12480
rect 4889 12474 4955 12477
rect 0 12472 4955 12474
rect 0 12416 4894 12472
rect 4950 12416 4955 12472
rect 0 12414 4955 12416
rect 0 12384 480 12414
rect 4889 12411 4955 12414
rect 7005 12474 7071 12477
rect 10409 12474 10475 12477
rect 7005 12472 10475 12474
rect 7005 12416 7010 12472
rect 7066 12416 10414 12472
rect 10470 12416 10475 12472
rect 7005 12414 10475 12416
rect 7005 12411 7071 12414
rect 10409 12411 10475 12414
rect 11462 12412 11468 12476
rect 11532 12474 11538 12476
rect 11697 12474 11763 12477
rect 11532 12472 11763 12474
rect 11532 12416 11702 12472
rect 11758 12416 11763 12472
rect 11532 12414 11763 12416
rect 11532 12412 11538 12414
rect 11697 12411 11763 12414
rect 11881 12474 11947 12477
rect 12249 12474 12315 12477
rect 11881 12472 12315 12474
rect 11881 12416 11886 12472
rect 11942 12416 12254 12472
rect 12310 12416 12315 12472
rect 11881 12414 12315 12416
rect 11881 12411 11947 12414
rect 12249 12411 12315 12414
rect 2405 12338 2471 12341
rect 3049 12338 3115 12341
rect 2405 12336 3115 12338
rect 2405 12280 2410 12336
rect 2466 12280 3054 12336
rect 3110 12280 3115 12336
rect 2405 12278 3115 12280
rect 2405 12275 2471 12278
rect 3049 12275 3115 12278
rect 9581 12338 9647 12341
rect 9806 12338 9812 12340
rect 9581 12336 9812 12338
rect 9581 12280 9586 12336
rect 9642 12280 9812 12336
rect 9581 12278 9812 12280
rect 9581 12275 9647 12278
rect 9806 12276 9812 12278
rect 9876 12338 9882 12340
rect 13670 12338 13676 12340
rect 9876 12278 13676 12338
rect 9876 12276 9882 12278
rect 13670 12276 13676 12278
rect 13740 12276 13746 12340
rect 5809 12202 5875 12205
rect 8385 12202 8451 12205
rect 5809 12200 8451 12202
rect 5809 12144 5814 12200
rect 5870 12144 8390 12200
rect 8446 12144 8451 12200
rect 5809 12142 8451 12144
rect 5809 12139 5875 12142
rect 8385 12139 8451 12142
rect 9806 12140 9812 12204
rect 9876 12202 9882 12204
rect 10133 12202 10199 12205
rect 9876 12200 10199 12202
rect 9876 12144 10138 12200
rect 10194 12144 10199 12200
rect 9876 12142 10199 12144
rect 9876 12140 9882 12142
rect 10133 12139 10199 12142
rect 4429 12066 4495 12069
rect 4889 12066 4955 12069
rect 4429 12064 4955 12066
rect 4429 12008 4434 12064
rect 4490 12008 4894 12064
rect 4950 12008 4955 12064
rect 4429 12006 4955 12008
rect 4429 12003 4495 12006
rect 4889 12003 4955 12006
rect 10174 12004 10180 12068
rect 10244 12066 10250 12068
rect 10317 12066 10383 12069
rect 12525 12066 12591 12069
rect 10244 12064 10383 12066
rect 10244 12008 10322 12064
rect 10378 12008 10383 12064
rect 10244 12006 10383 12008
rect 10244 12004 10250 12006
rect 10317 12003 10383 12006
rect 11286 12064 12591 12066
rect 11286 12008 12530 12064
rect 12586 12008 12591 12064
rect 11286 12006 12591 12008
rect 3409 12000 3729 12001
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 11935 3729 11936
rect 8340 12000 8660 12001
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 11935 8660 11936
rect 9581 11930 9647 11933
rect 11286 11932 11346 12006
rect 12525 12003 12591 12006
rect 13270 12000 13590 12001
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 11935 13590 11936
rect 11278 11930 11284 11932
rect 9581 11928 11284 11930
rect 9581 11872 9586 11928
rect 9642 11872 11284 11928
rect 9581 11870 11284 11872
rect 9581 11867 9647 11870
rect 11278 11868 11284 11870
rect 11348 11868 11354 11932
rect 12709 11930 12775 11933
rect 11608 11928 12775 11930
rect 11608 11872 12714 11928
rect 12770 11872 12775 11928
rect 11608 11870 12775 11872
rect 4521 11794 4587 11797
rect 10542 11794 10548 11796
rect 4521 11792 10548 11794
rect 4521 11736 4526 11792
rect 4582 11736 10548 11792
rect 4521 11734 10548 11736
rect 4521 11731 4587 11734
rect 10542 11732 10548 11734
rect 10612 11732 10618 11796
rect 10685 11794 10751 11797
rect 11145 11794 11211 11797
rect 11329 11794 11395 11797
rect 11608 11794 11668 11870
rect 12709 11867 12775 11870
rect 10685 11792 11395 11794
rect 10685 11736 10690 11792
rect 10746 11736 11150 11792
rect 11206 11736 11334 11792
rect 11390 11736 11395 11792
rect 10685 11734 11395 11736
rect 10685 11731 10751 11734
rect 11145 11731 11211 11734
rect 11329 11731 11395 11734
rect 11470 11734 11668 11794
rect 12433 11794 12499 11797
rect 13118 11794 13124 11796
rect 12433 11792 13124 11794
rect 12433 11736 12438 11792
rect 12494 11736 13124 11792
rect 12433 11734 13124 11736
rect 5349 11658 5415 11661
rect 11470 11658 11530 11734
rect 12433 11731 12499 11734
rect 13118 11732 13124 11734
rect 13188 11732 13194 11796
rect 5349 11656 11530 11658
rect 5349 11600 5354 11656
rect 5410 11600 11530 11656
rect 5349 11598 11530 11600
rect 12341 11658 12407 11661
rect 12341 11656 12634 11658
rect 12341 11600 12346 11656
rect 12402 11600 12634 11656
rect 12341 11598 12634 11600
rect 5349 11595 5415 11598
rect 12341 11595 12407 11598
rect 8661 11522 8727 11525
rect 8886 11522 8892 11524
rect 8661 11520 8892 11522
rect 8661 11464 8666 11520
rect 8722 11464 8892 11520
rect 8661 11462 8892 11464
rect 8661 11459 8727 11462
rect 8886 11460 8892 11462
rect 8956 11460 8962 11524
rect 9622 11460 9628 11524
rect 9692 11522 9698 11524
rect 10041 11522 10107 11525
rect 9692 11520 10107 11522
rect 9692 11464 10046 11520
rect 10102 11464 10107 11520
rect 9692 11462 10107 11464
rect 9692 11460 9698 11462
rect 10041 11459 10107 11462
rect 12065 11522 12131 11525
rect 12382 11522 12388 11524
rect 12065 11520 12388 11522
rect 12065 11464 12070 11520
rect 12126 11464 12388 11520
rect 12065 11462 12388 11464
rect 12065 11459 12131 11462
rect 12382 11460 12388 11462
rect 12452 11460 12458 11524
rect 5874 11456 6194 11457
rect 0 11386 480 11416
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6194 11456
rect 5874 11391 6194 11392
rect 10805 11456 11125 11457
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 11391 11125 11392
rect 3233 11386 3299 11389
rect 0 11384 3299 11386
rect 0 11328 3238 11384
rect 3294 11328 3299 11384
rect 0 11326 3299 11328
rect 0 11296 480 11326
rect 3233 11323 3299 11326
rect 6545 11386 6611 11389
rect 12433 11386 12499 11389
rect 6545 11384 10656 11386
rect 6545 11328 6550 11384
rect 6606 11328 10656 11384
rect 6545 11326 10656 11328
rect 6545 11323 6611 11326
rect 5625 11250 5691 11253
rect 9438 11250 9444 11252
rect 5625 11248 9444 11250
rect 5625 11192 5630 11248
rect 5686 11192 9444 11248
rect 5625 11190 9444 11192
rect 5625 11187 5691 11190
rect 9438 11188 9444 11190
rect 9508 11250 9514 11252
rect 9857 11250 9923 11253
rect 9508 11248 9923 11250
rect 9508 11192 9862 11248
rect 9918 11192 9923 11248
rect 9508 11190 9923 11192
rect 10596 11250 10656 11326
rect 11240 11384 12499 11386
rect 11240 11328 12438 11384
rect 12494 11328 12499 11384
rect 11240 11326 12499 11328
rect 11240 11250 11300 11326
rect 12433 11323 12499 11326
rect 10596 11190 11300 11250
rect 9508 11188 9514 11190
rect 9857 11187 9923 11190
rect 11462 11188 11468 11252
rect 11532 11250 11538 11252
rect 12014 11250 12020 11252
rect 11532 11190 12020 11250
rect 11532 11188 11538 11190
rect 12014 11188 12020 11190
rect 12084 11188 12090 11252
rect 12382 11188 12388 11252
rect 12452 11250 12458 11252
rect 12574 11250 12634 11598
rect 12452 11190 12634 11250
rect 12452 11188 12458 11190
rect 1945 11114 2011 11117
rect 13077 11114 13143 11117
rect 1945 11112 13143 11114
rect 1945 11056 1950 11112
rect 2006 11056 13082 11112
rect 13138 11056 13143 11112
rect 1945 11054 13143 11056
rect 1945 11051 2011 11054
rect 13077 11051 13143 11054
rect 11145 10978 11211 10981
rect 11462 10978 11468 10980
rect 11145 10976 11468 10978
rect 11145 10920 11150 10976
rect 11206 10920 11468 10976
rect 11145 10918 11468 10920
rect 11145 10915 11211 10918
rect 11462 10916 11468 10918
rect 11532 10916 11538 10980
rect 12014 10916 12020 10980
rect 12084 10978 12090 10980
rect 12433 10978 12499 10981
rect 12084 10976 12499 10978
rect 12084 10920 12438 10976
rect 12494 10920 12499 10976
rect 12084 10918 12499 10920
rect 12084 10916 12090 10918
rect 12433 10915 12499 10918
rect 3409 10912 3729 10913
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 10847 3729 10848
rect 8340 10912 8660 10913
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 10847 8660 10848
rect 13270 10912 13590 10913
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 10847 13590 10848
rect 4061 10842 4127 10845
rect 7097 10842 7163 10845
rect 4061 10840 7163 10842
rect 4061 10784 4066 10840
rect 4122 10784 7102 10840
rect 7158 10784 7163 10840
rect 4061 10782 7163 10784
rect 4061 10779 4127 10782
rect 7097 10779 7163 10782
rect 9990 10780 9996 10844
rect 10060 10842 10066 10844
rect 11462 10842 11468 10844
rect 10060 10782 11468 10842
rect 10060 10780 10066 10782
rect 11462 10780 11468 10782
rect 11532 10780 11538 10844
rect 11830 10780 11836 10844
rect 11900 10842 11906 10844
rect 11900 10782 12082 10842
rect 11900 10780 11906 10782
rect 2129 10706 2195 10709
rect 7281 10706 7347 10709
rect 9438 10706 9444 10708
rect 2129 10704 9444 10706
rect 2129 10648 2134 10704
rect 2190 10648 7286 10704
rect 7342 10648 9444 10704
rect 2129 10646 9444 10648
rect 2129 10643 2195 10646
rect 7281 10643 7347 10646
rect 9438 10644 9444 10646
rect 9508 10706 9514 10708
rect 9949 10706 10015 10709
rect 9508 10704 10015 10706
rect 9508 10648 9954 10704
rect 10010 10648 10015 10704
rect 9508 10646 10015 10648
rect 9508 10644 9514 10646
rect 9949 10643 10015 10646
rect 10409 10706 10475 10709
rect 11237 10706 11303 10709
rect 10409 10704 11303 10706
rect 10409 10648 10414 10704
rect 10470 10648 11242 10704
rect 11298 10648 11303 10704
rect 10409 10646 11303 10648
rect 10409 10643 10475 10646
rect 11237 10643 11303 10646
rect 5349 10570 5415 10573
rect 11053 10570 11119 10573
rect 5349 10568 11119 10570
rect 5349 10512 5354 10568
rect 5410 10512 11058 10568
rect 11114 10512 11119 10568
rect 5349 10510 11119 10512
rect 5349 10507 5415 10510
rect 11053 10507 11119 10510
rect 11237 10570 11303 10573
rect 12022 10570 12082 10782
rect 12433 10570 12499 10573
rect 11237 10568 12499 10570
rect 11237 10512 11242 10568
rect 11298 10512 12438 10568
rect 12494 10512 12499 10568
rect 11237 10510 12499 10512
rect 11237 10507 11303 10510
rect 12433 10507 12499 10510
rect 0 10434 480 10464
rect 1853 10434 1919 10437
rect 0 10432 1919 10434
rect 0 10376 1858 10432
rect 1914 10376 1919 10432
rect 0 10374 1919 10376
rect 0 10344 480 10374
rect 1853 10371 1919 10374
rect 3182 10372 3188 10436
rect 3252 10434 3258 10436
rect 3325 10434 3391 10437
rect 3252 10432 3391 10434
rect 3252 10376 3330 10432
rect 3386 10376 3391 10432
rect 3252 10374 3391 10376
rect 3252 10372 3258 10374
rect 3325 10371 3391 10374
rect 4429 10434 4495 10437
rect 5717 10434 5783 10437
rect 4429 10432 5783 10434
rect 4429 10376 4434 10432
rect 4490 10376 5722 10432
rect 5778 10376 5783 10432
rect 4429 10374 5783 10376
rect 4429 10371 4495 10374
rect 5717 10371 5783 10374
rect 7005 10434 7071 10437
rect 9029 10434 9095 10437
rect 7005 10432 9095 10434
rect 7005 10376 7010 10432
rect 7066 10376 9034 10432
rect 9090 10376 9095 10432
rect 7005 10374 9095 10376
rect 7005 10371 7071 10374
rect 9029 10371 9095 10374
rect 11830 10372 11836 10436
rect 11900 10434 11906 10436
rect 12382 10434 12388 10436
rect 11900 10374 12388 10434
rect 11900 10372 11906 10374
rect 12382 10372 12388 10374
rect 12452 10372 12458 10436
rect 12934 10372 12940 10436
rect 13004 10434 13010 10436
rect 13445 10434 13511 10437
rect 13004 10432 13511 10434
rect 13004 10376 13450 10432
rect 13506 10376 13511 10432
rect 13004 10374 13511 10376
rect 13004 10372 13010 10374
rect 13445 10371 13511 10374
rect 5874 10368 6194 10369
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6194 10368
rect 5874 10303 6194 10304
rect 10805 10368 11125 10369
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 10303 11125 10304
rect 4429 10298 4495 10301
rect 4705 10298 4771 10301
rect 9489 10298 9555 10301
rect 4429 10296 4771 10298
rect 4429 10240 4434 10296
rect 4490 10240 4710 10296
rect 4766 10240 4771 10296
rect 4429 10238 4771 10240
rect 4429 10235 4495 10238
rect 4705 10235 4771 10238
rect 6502 10296 9555 10298
rect 6502 10240 9494 10296
rect 9550 10240 9555 10296
rect 6502 10238 9555 10240
rect 2589 10162 2655 10165
rect 6502 10162 6562 10238
rect 9489 10235 9555 10238
rect 9857 10298 9923 10301
rect 10409 10298 10475 10301
rect 15009 10298 15075 10301
rect 9857 10296 10475 10298
rect 9857 10240 9862 10296
rect 9918 10240 10414 10296
rect 10470 10240 10475 10296
rect 9857 10238 10475 10240
rect 9857 10235 9923 10238
rect 10409 10235 10475 10238
rect 12344 10296 15075 10298
rect 12344 10240 15014 10296
rect 15070 10240 15075 10296
rect 12344 10238 15075 10240
rect 2589 10160 6562 10162
rect 2589 10104 2594 10160
rect 2650 10104 6562 10160
rect 2589 10102 6562 10104
rect 6637 10162 6703 10165
rect 12344 10162 12404 10238
rect 15009 10235 15075 10238
rect 6637 10160 12404 10162
rect 6637 10104 6642 10160
rect 6698 10104 12404 10160
rect 6637 10102 12404 10104
rect 2589 10099 2655 10102
rect 6637 10099 6703 10102
rect 12750 10100 12756 10164
rect 12820 10162 12826 10164
rect 13353 10162 13419 10165
rect 13721 10164 13787 10165
rect 13670 10162 13676 10164
rect 12820 10160 13419 10162
rect 12820 10104 13358 10160
rect 13414 10104 13419 10160
rect 12820 10102 13419 10104
rect 13630 10102 13676 10162
rect 13740 10160 13787 10164
rect 13782 10104 13787 10160
rect 12820 10100 12826 10102
rect 13353 10099 13419 10102
rect 13670 10100 13676 10102
rect 13740 10100 13787 10104
rect 13721 10099 13787 10100
rect 4705 10026 4771 10029
rect 6361 10026 6427 10029
rect 4705 10024 6427 10026
rect 4705 9968 4710 10024
rect 4766 9968 6366 10024
rect 6422 9968 6427 10024
rect 4705 9966 6427 9968
rect 4705 9963 4771 9966
rect 6361 9963 6427 9966
rect 6729 10026 6795 10029
rect 14641 10026 14707 10029
rect 6729 10024 14707 10026
rect 6729 9968 6734 10024
rect 6790 9968 14646 10024
rect 14702 9968 14707 10024
rect 6729 9966 14707 9968
rect 6729 9963 6795 9966
rect 14641 9963 14707 9966
rect 14917 10026 14983 10029
rect 16520 10026 17000 10056
rect 14917 10024 17000 10026
rect 14917 9968 14922 10024
rect 14978 9968 17000 10024
rect 14917 9966 17000 9968
rect 14917 9963 14983 9966
rect 16520 9936 17000 9966
rect 5625 9890 5691 9893
rect 8017 9890 8083 9893
rect 5625 9888 8083 9890
rect 5625 9832 5630 9888
rect 5686 9832 8022 9888
rect 8078 9832 8083 9888
rect 5625 9830 8083 9832
rect 5625 9827 5691 9830
rect 8017 9827 8083 9830
rect 8753 9890 8819 9893
rect 11329 9890 11395 9893
rect 11697 9892 11763 9893
rect 8753 9888 11395 9890
rect 8753 9832 8758 9888
rect 8814 9832 11334 9888
rect 11390 9832 11395 9888
rect 8753 9830 11395 9832
rect 8753 9827 8819 9830
rect 11329 9827 11395 9830
rect 11646 9828 11652 9892
rect 11716 9890 11763 9892
rect 12065 9890 12131 9893
rect 12198 9890 12204 9892
rect 11716 9888 11808 9890
rect 11758 9832 11808 9888
rect 11716 9830 11808 9832
rect 12065 9888 12204 9890
rect 12065 9832 12070 9888
rect 12126 9832 12204 9888
rect 12065 9830 12204 9832
rect 11716 9828 11763 9830
rect 11697 9827 11763 9828
rect 12065 9827 12131 9830
rect 12198 9828 12204 9830
rect 12268 9828 12274 9892
rect 3409 9824 3729 9825
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 9759 3729 9760
rect 8340 9824 8660 9825
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 9759 8660 9760
rect 13270 9824 13590 9825
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 9759 13590 9760
rect 4521 9754 4587 9757
rect 5257 9754 5323 9757
rect 4521 9752 5323 9754
rect 4521 9696 4526 9752
rect 4582 9696 5262 9752
rect 5318 9696 5323 9752
rect 4521 9694 5323 9696
rect 4521 9691 4587 9694
rect 5257 9691 5323 9694
rect 5441 9754 5507 9757
rect 7189 9754 7255 9757
rect 5441 9752 7255 9754
rect 5441 9696 5446 9752
rect 5502 9696 7194 9752
rect 7250 9696 7255 9752
rect 5441 9694 7255 9696
rect 5441 9691 5507 9694
rect 7189 9691 7255 9694
rect 9070 9692 9076 9756
rect 9140 9754 9146 9756
rect 9765 9754 9831 9757
rect 9140 9752 9831 9754
rect 9140 9696 9770 9752
rect 9826 9696 9831 9752
rect 9140 9694 9831 9696
rect 9140 9692 9146 9694
rect 9765 9691 9831 9694
rect 9990 9692 9996 9756
rect 10060 9754 10066 9756
rect 10060 9694 12772 9754
rect 10060 9692 10066 9694
rect 2497 9618 2563 9621
rect 12433 9618 12499 9621
rect 2497 9616 12499 9618
rect 2497 9560 2502 9616
rect 2558 9560 12438 9616
rect 12494 9560 12499 9616
rect 2497 9558 12499 9560
rect 2497 9555 2563 9558
rect 12433 9555 12499 9558
rect 0 9482 480 9512
rect 4981 9482 5047 9485
rect 5809 9482 5875 9485
rect 0 9422 2330 9482
rect 0 9392 480 9422
rect 2270 8938 2330 9422
rect 4981 9480 5875 9482
rect 4981 9424 4986 9480
rect 5042 9424 5814 9480
rect 5870 9424 5875 9480
rect 4981 9422 5875 9424
rect 4981 9419 5047 9422
rect 5809 9419 5875 9422
rect 8477 9482 8543 9485
rect 10501 9482 10567 9485
rect 8477 9480 10567 9482
rect 8477 9424 8482 9480
rect 8538 9424 10506 9480
rect 10562 9424 10567 9480
rect 8477 9422 10567 9424
rect 8477 9419 8543 9422
rect 10501 9419 10567 9422
rect 10777 9482 10843 9485
rect 11421 9482 11487 9485
rect 10777 9480 11487 9482
rect 10777 9424 10782 9480
rect 10838 9424 11426 9480
rect 11482 9424 11487 9480
rect 10777 9422 11487 9424
rect 10777 9419 10843 9422
rect 11421 9419 11487 9422
rect 12198 9420 12204 9484
rect 12268 9482 12274 9484
rect 12525 9482 12591 9485
rect 12268 9480 12591 9482
rect 12268 9424 12530 9480
rect 12586 9424 12591 9480
rect 12268 9422 12591 9424
rect 12712 9482 12772 9694
rect 13905 9482 13971 9485
rect 12712 9480 13971 9482
rect 12712 9424 13910 9480
rect 13966 9424 13971 9480
rect 12712 9422 13971 9424
rect 12268 9420 12274 9422
rect 12525 9419 12591 9422
rect 13905 9419 13971 9422
rect 3601 9346 3667 9349
rect 4245 9346 4311 9349
rect 3601 9344 4311 9346
rect 3601 9288 3606 9344
rect 3662 9288 4250 9344
rect 4306 9288 4311 9344
rect 3601 9286 4311 9288
rect 3601 9283 3667 9286
rect 4245 9283 4311 9286
rect 4521 9346 4587 9349
rect 5717 9346 5783 9349
rect 9489 9348 9555 9349
rect 4521 9344 5783 9346
rect 4521 9288 4526 9344
rect 4582 9288 5722 9344
rect 5778 9288 5783 9344
rect 4521 9286 5783 9288
rect 4521 9283 4587 9286
rect 5717 9283 5783 9286
rect 9438 9284 9444 9348
rect 9508 9346 9555 9348
rect 9765 9346 9831 9349
rect 10501 9346 10567 9349
rect 9508 9344 9600 9346
rect 9550 9288 9600 9344
rect 9508 9286 9600 9288
rect 9765 9344 10567 9346
rect 9765 9288 9770 9344
rect 9826 9288 10506 9344
rect 10562 9288 10567 9344
rect 9765 9286 10567 9288
rect 9508 9284 9555 9286
rect 9489 9283 9555 9284
rect 9765 9283 9831 9286
rect 10501 9283 10567 9286
rect 5874 9280 6194 9281
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6194 9280
rect 5874 9215 6194 9216
rect 10805 9280 11125 9281
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 9215 11125 9216
rect 3693 9210 3759 9213
rect 5165 9210 5231 9213
rect 3693 9208 5231 9210
rect 3693 9152 3698 9208
rect 3754 9152 5170 9208
rect 5226 9152 5231 9208
rect 3693 9150 5231 9152
rect 3693 9147 3759 9150
rect 5165 9147 5231 9150
rect 7649 9210 7715 9213
rect 8661 9210 8727 9213
rect 7649 9208 8727 9210
rect 7649 9152 7654 9208
rect 7710 9152 8666 9208
rect 8722 9152 8727 9208
rect 7649 9150 8727 9152
rect 7649 9147 7715 9150
rect 8661 9147 8727 9150
rect 10133 9212 10199 9213
rect 10133 9208 10180 9212
rect 10244 9210 10250 9212
rect 11424 9210 11484 9419
rect 11830 9284 11836 9348
rect 11900 9346 11906 9348
rect 13169 9346 13235 9349
rect 11900 9344 13235 9346
rect 11900 9288 13174 9344
rect 13230 9288 13235 9344
rect 11900 9286 13235 9288
rect 11900 9284 11906 9286
rect 13169 9283 13235 9286
rect 12382 9210 12388 9212
rect 10133 9152 10138 9208
rect 10133 9148 10180 9152
rect 10244 9150 10290 9210
rect 11424 9150 12388 9210
rect 10244 9148 10250 9150
rect 12382 9148 12388 9150
rect 12452 9148 12458 9212
rect 12893 9210 12959 9213
rect 13169 9210 13235 9213
rect 12893 9208 13235 9210
rect 12893 9152 12898 9208
rect 12954 9152 13174 9208
rect 13230 9152 13235 9208
rect 12893 9150 13235 9152
rect 10133 9147 10199 9148
rect 12893 9147 12959 9150
rect 13169 9147 13235 9150
rect 2446 9012 2452 9076
rect 2516 9074 2522 9076
rect 3693 9074 3759 9077
rect 9622 9074 9628 9076
rect 2516 9072 9628 9074
rect 2516 9016 3698 9072
rect 3754 9016 9628 9072
rect 2516 9014 9628 9016
rect 2516 9012 2522 9014
rect 3693 9011 3759 9014
rect 9622 9012 9628 9014
rect 9692 9074 9698 9076
rect 11278 9074 11284 9076
rect 9692 9014 11284 9074
rect 9692 9012 9698 9014
rect 11278 9012 11284 9014
rect 11348 9074 11354 9076
rect 13261 9074 13327 9077
rect 11348 9072 13327 9074
rect 11348 9016 13266 9072
rect 13322 9016 13327 9072
rect 11348 9014 13327 9016
rect 11348 9012 11354 9014
rect 13261 9011 13327 9014
rect 4797 8938 4863 8941
rect 15009 8938 15075 8941
rect 2270 8936 4863 8938
rect 2270 8880 4802 8936
rect 4858 8880 4863 8936
rect 2270 8878 4863 8880
rect 4797 8875 4863 8878
rect 7238 8936 15075 8938
rect 7238 8880 15014 8936
rect 15070 8880 15075 8936
rect 7238 8878 15075 8880
rect 6453 8802 6519 8805
rect 7238 8802 7298 8878
rect 15009 8875 15075 8878
rect 6453 8800 7298 8802
rect 6453 8744 6458 8800
rect 6514 8744 7298 8800
rect 6453 8742 7298 8744
rect 9581 8802 9647 8805
rect 10777 8802 10843 8805
rect 9581 8800 10843 8802
rect 9581 8744 9586 8800
rect 9642 8744 10782 8800
rect 10838 8744 10843 8800
rect 9581 8742 10843 8744
rect 6453 8739 6519 8742
rect 9581 8739 9647 8742
rect 10777 8739 10843 8742
rect 11646 8740 11652 8804
rect 11716 8802 11722 8804
rect 12525 8802 12591 8805
rect 13118 8802 13124 8804
rect 11716 8742 12450 8802
rect 11716 8740 11722 8742
rect 3409 8736 3729 8737
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 8671 3729 8672
rect 8340 8736 8660 8737
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 8671 8660 8672
rect 9029 8666 9095 8669
rect 11973 8666 12039 8669
rect 9029 8664 12039 8666
rect 9029 8608 9034 8664
rect 9090 8608 11978 8664
rect 12034 8608 12039 8664
rect 9029 8606 12039 8608
rect 12390 8666 12450 8742
rect 12525 8800 13124 8802
rect 12525 8744 12530 8800
rect 12586 8744 13124 8800
rect 12525 8742 13124 8744
rect 12525 8739 12591 8742
rect 13118 8740 13124 8742
rect 13188 8740 13194 8804
rect 13270 8736 13590 8737
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 8671 13590 8672
rect 12566 8666 12572 8668
rect 12390 8606 12572 8666
rect 9029 8603 9095 8606
rect 11973 8603 12039 8606
rect 12566 8604 12572 8606
rect 12636 8604 12642 8668
rect 13905 8666 13971 8669
rect 14406 8666 14412 8668
rect 13905 8664 14412 8666
rect 13905 8608 13910 8664
rect 13966 8608 14412 8664
rect 13905 8606 14412 8608
rect 13905 8603 13971 8606
rect 14406 8604 14412 8606
rect 14476 8604 14482 8668
rect 3969 8530 4035 8533
rect 4613 8530 4679 8533
rect 6678 8530 6684 8532
rect 3969 8528 6684 8530
rect 3969 8472 3974 8528
rect 4030 8472 4618 8528
rect 4674 8472 6684 8528
rect 3969 8470 6684 8472
rect 3969 8467 4035 8470
rect 4613 8467 4679 8470
rect 6678 8468 6684 8470
rect 6748 8530 6754 8532
rect 8886 8530 8892 8532
rect 6748 8470 8892 8530
rect 6748 8468 6754 8470
rect 8886 8468 8892 8470
rect 8956 8468 8962 8532
rect 9029 8530 9095 8533
rect 9806 8530 9812 8532
rect 9029 8528 9812 8530
rect 9029 8472 9034 8528
rect 9090 8472 9812 8528
rect 9029 8470 9812 8472
rect 9029 8467 9095 8470
rect 9806 8468 9812 8470
rect 9876 8530 9882 8532
rect 12014 8530 12020 8532
rect 9876 8470 12020 8530
rect 9876 8468 9882 8470
rect 12014 8468 12020 8470
rect 12084 8468 12090 8532
rect 12566 8468 12572 8532
rect 12636 8530 12642 8532
rect 12801 8530 12867 8533
rect 12636 8528 12867 8530
rect 12636 8472 12806 8528
rect 12862 8472 12867 8528
rect 12636 8470 12867 8472
rect 12636 8468 12642 8470
rect 12801 8467 12867 8470
rect 0 8394 480 8424
rect 1209 8394 1275 8397
rect 0 8392 1275 8394
rect 0 8336 1214 8392
rect 1270 8336 1275 8392
rect 0 8334 1275 8336
rect 0 8304 480 8334
rect 1209 8331 1275 8334
rect 2957 8394 3023 8397
rect 12525 8394 12591 8397
rect 2957 8392 12591 8394
rect 2957 8336 2962 8392
rect 3018 8336 12530 8392
rect 12586 8336 12591 8392
rect 2957 8334 12591 8336
rect 2957 8331 3023 8334
rect 12525 8331 12591 8334
rect 9121 8260 9187 8261
rect 9070 8196 9076 8260
rect 9140 8258 9187 8260
rect 9140 8256 9232 8258
rect 9182 8200 9232 8256
rect 9140 8198 9232 8200
rect 9140 8196 9187 8198
rect 11278 8196 11284 8260
rect 11348 8258 11354 8260
rect 13169 8258 13235 8261
rect 11348 8256 13235 8258
rect 11348 8200 13174 8256
rect 13230 8200 13235 8256
rect 11348 8198 13235 8200
rect 11348 8196 11354 8198
rect 9121 8195 9187 8196
rect 13169 8195 13235 8198
rect 5874 8192 6194 8193
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6194 8192
rect 5874 8127 6194 8128
rect 10805 8192 11125 8193
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 8127 11125 8128
rect 2405 8122 2471 8125
rect 6361 8122 6427 8125
rect 9029 8122 9095 8125
rect 11513 8124 11579 8125
rect 2405 8120 2744 8122
rect 2405 8064 2410 8120
rect 2466 8064 2744 8120
rect 2405 8062 2744 8064
rect 2405 8059 2471 8062
rect 1669 7986 1735 7989
rect 2405 7986 2471 7989
rect 1669 7984 2471 7986
rect 1669 7928 1674 7984
rect 1730 7928 2410 7984
rect 2466 7928 2471 7984
rect 1669 7926 2471 7928
rect 1669 7923 1735 7926
rect 2405 7923 2471 7926
rect 2684 7850 2744 8062
rect 6361 8120 9095 8122
rect 6361 8064 6366 8120
rect 6422 8064 9034 8120
rect 9090 8064 9095 8120
rect 6361 8062 9095 8064
rect 6361 8059 6427 8062
rect 9029 8059 9095 8062
rect 11462 8060 11468 8124
rect 11532 8122 11579 8124
rect 11697 8122 11763 8125
rect 12065 8122 12131 8125
rect 11532 8120 11624 8122
rect 11574 8064 11624 8120
rect 11532 8062 11624 8064
rect 11697 8120 12131 8122
rect 11697 8064 11702 8120
rect 11758 8064 12070 8120
rect 12126 8064 12131 8120
rect 11697 8062 12131 8064
rect 11532 8060 11579 8062
rect 11513 8059 11579 8060
rect 11697 8059 11763 8062
rect 12065 8059 12131 8062
rect 12617 8122 12683 8125
rect 13670 8122 13676 8124
rect 12617 8120 13676 8122
rect 12617 8064 12622 8120
rect 12678 8064 13676 8120
rect 12617 8062 13676 8064
rect 12617 8059 12683 8062
rect 13670 8060 13676 8062
rect 13740 8060 13746 8124
rect 3509 7986 3575 7989
rect 4613 7986 4679 7989
rect 3509 7984 4679 7986
rect 3509 7928 3514 7984
rect 3570 7928 4618 7984
rect 4674 7928 4679 7984
rect 3509 7926 4679 7928
rect 3509 7923 3575 7926
rect 4613 7923 4679 7926
rect 5717 7986 5783 7989
rect 9397 7986 9463 7989
rect 5717 7984 9463 7986
rect 5717 7928 5722 7984
rect 5778 7928 9402 7984
rect 9458 7928 9463 7984
rect 5717 7926 9463 7928
rect 5717 7923 5783 7926
rect 9397 7923 9463 7926
rect 10409 7986 10475 7989
rect 14549 7986 14615 7989
rect 10409 7984 14615 7986
rect 10409 7928 10414 7984
rect 10470 7928 14554 7984
rect 14610 7928 14615 7984
rect 10409 7926 14615 7928
rect 10409 7923 10475 7926
rect 14549 7923 14615 7926
rect 13261 7850 13327 7853
rect 2684 7848 13327 7850
rect 2684 7792 13266 7848
rect 13322 7792 13327 7848
rect 2684 7790 13327 7792
rect 13261 7787 13327 7790
rect 3969 7714 4035 7717
rect 8201 7714 8267 7717
rect 3969 7712 8267 7714
rect 3969 7656 3974 7712
rect 4030 7656 8206 7712
rect 8262 7656 8267 7712
rect 3969 7654 8267 7656
rect 3969 7651 4035 7654
rect 8201 7651 8267 7654
rect 10225 7714 10291 7717
rect 12750 7714 12756 7716
rect 10225 7712 12756 7714
rect 10225 7656 10230 7712
rect 10286 7656 12756 7712
rect 10225 7654 12756 7656
rect 10225 7651 10291 7654
rect 12750 7652 12756 7654
rect 12820 7652 12826 7716
rect 3409 7648 3729 7649
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 7583 3729 7584
rect 8340 7648 8660 7649
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 7583 8660 7584
rect 13270 7648 13590 7649
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 7583 13590 7584
rect 5533 7578 5599 7581
rect 8109 7578 8175 7581
rect 5533 7576 8175 7578
rect 5533 7520 5538 7576
rect 5594 7520 8114 7576
rect 8170 7520 8175 7576
rect 5533 7518 8175 7520
rect 5533 7515 5599 7518
rect 8109 7515 8175 7518
rect 9581 7578 9647 7581
rect 10869 7578 10935 7581
rect 9581 7576 10935 7578
rect 9581 7520 9586 7576
rect 9642 7520 10874 7576
rect 10930 7520 10935 7576
rect 9581 7518 10935 7520
rect 9581 7515 9647 7518
rect 10869 7515 10935 7518
rect 11145 7578 11211 7581
rect 11278 7578 11284 7580
rect 11145 7576 11284 7578
rect 11145 7520 11150 7576
rect 11206 7520 11284 7576
rect 11145 7518 11284 7520
rect 11145 7515 11211 7518
rect 11278 7516 11284 7518
rect 11348 7516 11354 7580
rect 11789 7578 11855 7581
rect 12014 7578 12020 7580
rect 11789 7576 12020 7578
rect 11789 7520 11794 7576
rect 11850 7520 12020 7576
rect 11789 7518 12020 7520
rect 11789 7515 11855 7518
rect 12014 7516 12020 7518
rect 12084 7516 12090 7580
rect 12198 7516 12204 7580
rect 12268 7578 12274 7580
rect 12433 7578 12499 7581
rect 12268 7576 12499 7578
rect 12268 7520 12438 7576
rect 12494 7520 12499 7576
rect 12268 7518 12499 7520
rect 12268 7516 12274 7518
rect 12433 7515 12499 7518
rect 12566 7516 12572 7580
rect 12636 7578 12642 7580
rect 12893 7578 12959 7581
rect 12636 7576 12959 7578
rect 12636 7520 12898 7576
rect 12954 7520 12959 7576
rect 12636 7518 12959 7520
rect 12636 7516 12642 7518
rect 12893 7515 12959 7518
rect 0 7442 480 7472
rect 3049 7442 3115 7445
rect 0 7440 3115 7442
rect 0 7384 3054 7440
rect 3110 7384 3115 7440
rect 0 7382 3115 7384
rect 0 7352 480 7382
rect 3049 7379 3115 7382
rect 4981 7442 5047 7445
rect 10041 7442 10107 7445
rect 4981 7440 10107 7442
rect 4981 7384 4986 7440
rect 5042 7384 10046 7440
rect 10102 7384 10107 7440
rect 4981 7382 10107 7384
rect 4981 7379 5047 7382
rect 10041 7379 10107 7382
rect 10317 7442 10383 7445
rect 14641 7442 14707 7445
rect 10317 7440 14707 7442
rect 10317 7384 10322 7440
rect 10378 7384 14646 7440
rect 14702 7384 14707 7440
rect 10317 7382 14707 7384
rect 10317 7379 10383 7382
rect 14641 7379 14707 7382
rect 1853 7306 1919 7309
rect 13629 7306 13695 7309
rect 1853 7304 13695 7306
rect 1853 7248 1858 7304
rect 1914 7248 13634 7304
rect 13690 7248 13695 7304
rect 1853 7246 13695 7248
rect 1853 7243 1919 7246
rect 13629 7243 13695 7246
rect 4797 7170 4863 7173
rect 5717 7170 5783 7173
rect 4797 7168 5783 7170
rect 4797 7112 4802 7168
rect 4858 7112 5722 7168
rect 5778 7112 5783 7168
rect 4797 7110 5783 7112
rect 4797 7107 4863 7110
rect 5717 7107 5783 7110
rect 6361 7170 6427 7173
rect 10041 7170 10107 7173
rect 6361 7168 10107 7170
rect 6361 7112 6366 7168
rect 6422 7112 10046 7168
rect 10102 7112 10107 7168
rect 6361 7110 10107 7112
rect 6361 7107 6427 7110
rect 10041 7107 10107 7110
rect 12801 7170 12867 7173
rect 13118 7170 13124 7172
rect 12801 7168 13124 7170
rect 12801 7112 12806 7168
rect 12862 7112 13124 7168
rect 12801 7110 13124 7112
rect 12801 7107 12867 7110
rect 13118 7108 13124 7110
rect 13188 7108 13194 7172
rect 5874 7104 6194 7105
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6194 7104
rect 5874 7039 6194 7040
rect 10805 7104 11125 7105
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 7039 11125 7040
rect 2129 7034 2195 7037
rect 2957 7034 3023 7037
rect 2129 7032 3023 7034
rect 2129 6976 2134 7032
rect 2190 6976 2962 7032
rect 3018 6976 3023 7032
rect 2129 6974 3023 6976
rect 2129 6971 2195 6974
rect 2957 6971 3023 6974
rect 4429 7034 4495 7037
rect 10317 7034 10383 7037
rect 4429 7032 5642 7034
rect 4429 6976 4434 7032
rect 4490 6976 5642 7032
rect 4429 6974 5642 6976
rect 4429 6971 4495 6974
rect 5582 6898 5642 6974
rect 6318 7032 10383 7034
rect 6318 6976 10322 7032
rect 10378 6976 10383 7032
rect 6318 6974 10383 6976
rect 6318 6898 6378 6974
rect 10317 6971 10383 6974
rect 5582 6838 6378 6898
rect 7833 6898 7899 6901
rect 9765 6898 9831 6901
rect 10961 6898 11027 6901
rect 7833 6896 11027 6898
rect 7833 6840 7838 6896
rect 7894 6840 9770 6896
rect 9826 6840 10966 6896
rect 11022 6840 11027 6896
rect 7833 6838 11027 6840
rect 7833 6835 7899 6838
rect 9765 6835 9831 6838
rect 10961 6835 11027 6838
rect 11145 6898 11211 6901
rect 11462 6898 11468 6900
rect 11145 6896 11468 6898
rect 11145 6840 11150 6896
rect 11206 6840 11468 6896
rect 11145 6838 11468 6840
rect 11145 6835 11211 6838
rect 11462 6836 11468 6838
rect 11532 6836 11538 6900
rect 13813 6898 13879 6901
rect 12942 6896 13879 6898
rect 12942 6840 13818 6896
rect 13874 6840 13879 6896
rect 12942 6838 13879 6840
rect 5349 6762 5415 6765
rect 12942 6762 13002 6838
rect 13813 6835 13879 6838
rect 15009 6762 15075 6765
rect 5349 6760 13002 6762
rect 5349 6704 5354 6760
rect 5410 6704 13002 6760
rect 5349 6702 13002 6704
rect 13126 6760 15075 6762
rect 13126 6704 15014 6760
rect 15070 6704 15075 6760
rect 13126 6702 15075 6704
rect 5349 6699 5415 6702
rect 5165 6626 5231 6629
rect 5441 6626 5507 6629
rect 8201 6626 8267 6629
rect 5165 6624 8267 6626
rect 5165 6568 5170 6624
rect 5226 6568 5446 6624
rect 5502 6568 8206 6624
rect 8262 6568 8267 6624
rect 5165 6566 8267 6568
rect 5165 6563 5231 6566
rect 5441 6563 5507 6566
rect 8201 6563 8267 6566
rect 9254 6564 9260 6628
rect 9324 6626 9330 6628
rect 10041 6626 10107 6629
rect 9324 6624 10107 6626
rect 9324 6568 10046 6624
rect 10102 6568 10107 6624
rect 9324 6566 10107 6568
rect 9324 6564 9330 6566
rect 10041 6563 10107 6566
rect 3409 6560 3729 6561
rect 0 6490 480 6520
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 2865 6490 2931 6493
rect 0 6488 2931 6490
rect 0 6432 2870 6488
rect 2926 6432 2931 6488
rect 0 6430 2931 6432
rect 0 6400 480 6430
rect 2865 6427 2931 6430
rect 4613 6490 4679 6493
rect 8109 6490 8175 6493
rect 4613 6488 8175 6490
rect 4613 6432 4618 6488
rect 4674 6432 8114 6488
rect 8170 6432 8175 6488
rect 4613 6430 8175 6432
rect 4613 6427 4679 6430
rect 8109 6427 8175 6430
rect 9397 6490 9463 6493
rect 13126 6490 13186 6702
rect 15009 6699 15075 6702
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 9397 6488 13186 6490
rect 9397 6432 9402 6488
rect 9458 6432 13186 6488
rect 9397 6430 13186 6432
rect 9397 6427 9463 6430
rect 2589 6354 2655 6357
rect 13445 6354 13511 6357
rect 2589 6352 13511 6354
rect 2589 6296 2594 6352
rect 2650 6296 13450 6352
rect 13506 6296 13511 6352
rect 2589 6294 13511 6296
rect 2589 6291 2655 6294
rect 13445 6291 13511 6294
rect 2221 6218 2287 6221
rect 2446 6218 2452 6220
rect 2221 6216 2452 6218
rect 2221 6160 2226 6216
rect 2282 6160 2452 6216
rect 2221 6158 2452 6160
rect 2221 6155 2287 6158
rect 2446 6156 2452 6158
rect 2516 6156 2522 6220
rect 3785 6218 3851 6221
rect 9397 6218 9463 6221
rect 12433 6220 12499 6221
rect 3785 6216 9463 6218
rect 3785 6160 3790 6216
rect 3846 6160 9402 6216
rect 9458 6160 9463 6216
rect 3785 6158 9463 6160
rect 3785 6155 3851 6158
rect 9397 6155 9463 6158
rect 9998 6158 11300 6218
rect 6913 6082 6979 6085
rect 9765 6082 9831 6085
rect 6913 6080 9831 6082
rect 6913 6024 6918 6080
rect 6974 6024 9770 6080
rect 9826 6024 9831 6080
rect 6913 6022 9831 6024
rect 6913 6019 6979 6022
rect 9765 6019 9831 6022
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 4521 5810 4587 5813
rect 9998 5810 10058 6158
rect 11240 6082 11300 6158
rect 12382 6156 12388 6220
rect 12452 6218 12499 6220
rect 12452 6216 12544 6218
rect 12494 6160 12544 6216
rect 12452 6158 12544 6160
rect 12452 6156 12499 6158
rect 12433 6155 12499 6156
rect 15561 6082 15627 6085
rect 11240 6080 15627 6082
rect 11240 6024 15566 6080
rect 15622 6024 15627 6080
rect 11240 6022 15627 6024
rect 15561 6019 15627 6022
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 11237 5946 11303 5949
rect 13670 5946 13676 5948
rect 11237 5944 13676 5946
rect 11237 5888 11242 5944
rect 11298 5888 13676 5944
rect 11237 5886 13676 5888
rect 11237 5883 11303 5886
rect 13670 5884 13676 5886
rect 13740 5884 13746 5948
rect 4521 5808 10058 5810
rect 4521 5752 4526 5808
rect 4582 5752 10058 5808
rect 4521 5750 10058 5752
rect 10133 5810 10199 5813
rect 13813 5810 13879 5813
rect 10133 5808 13879 5810
rect 10133 5752 10138 5808
rect 10194 5752 13818 5808
rect 13874 5752 13879 5808
rect 10133 5750 13879 5752
rect 4521 5747 4587 5750
rect 10133 5747 10199 5750
rect 13813 5747 13879 5750
rect 4061 5672 4127 5677
rect 4061 5616 4066 5672
rect 4122 5616 4127 5672
rect 4061 5611 4127 5616
rect 7557 5674 7623 5677
rect 12801 5674 12867 5677
rect 7557 5672 12867 5674
rect 7557 5616 7562 5672
rect 7618 5616 12806 5672
rect 12862 5616 12867 5672
rect 7557 5614 12867 5616
rect 7557 5611 7623 5614
rect 12801 5611 12867 5614
rect 14038 5612 14044 5676
rect 14108 5674 14114 5676
rect 14181 5674 14247 5677
rect 14108 5672 14247 5674
rect 14108 5616 14186 5672
rect 14242 5616 14247 5672
rect 14108 5614 14247 5616
rect 14108 5612 14114 5614
rect 14181 5611 14247 5614
rect 3409 5472 3729 5473
rect 0 5402 480 5432
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 1485 5402 1551 5405
rect 0 5400 1551 5402
rect 0 5344 1490 5400
rect 1546 5344 1551 5400
rect 0 5342 1551 5344
rect 4064 5402 4124 5611
rect 9305 5538 9371 5541
rect 9622 5538 9628 5540
rect 9305 5536 9628 5538
rect 9305 5480 9310 5536
rect 9366 5480 9628 5536
rect 9305 5478 9628 5480
rect 9305 5475 9371 5478
rect 9622 5476 9628 5478
rect 9692 5476 9698 5540
rect 12566 5476 12572 5540
rect 12636 5538 12642 5540
rect 12709 5538 12775 5541
rect 12636 5536 12775 5538
rect 12636 5480 12714 5536
rect 12770 5480 12775 5536
rect 12636 5478 12775 5480
rect 12636 5476 12642 5478
rect 12709 5475 12775 5478
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 7741 5402 7807 5405
rect 4064 5400 7807 5402
rect 4064 5344 7746 5400
rect 7802 5344 7807 5400
rect 4064 5342 7807 5344
rect 0 5312 480 5342
rect 1485 5339 1551 5342
rect 7741 5339 7807 5342
rect 8886 5340 8892 5404
rect 8956 5402 8962 5404
rect 11421 5402 11487 5405
rect 8956 5400 11487 5402
rect 8956 5344 11426 5400
rect 11482 5344 11487 5400
rect 8956 5342 11487 5344
rect 8956 5340 8962 5342
rect 11421 5339 11487 5342
rect 4245 5266 4311 5269
rect 13445 5266 13511 5269
rect 4245 5264 13511 5266
rect 4245 5208 4250 5264
rect 4306 5208 13450 5264
rect 13506 5208 13511 5264
rect 4245 5206 13511 5208
rect 4245 5203 4311 5206
rect 13445 5203 13511 5206
rect 3509 5130 3575 5133
rect 9765 5130 9831 5133
rect 3509 5128 9831 5130
rect 3509 5072 3514 5128
rect 3570 5072 9770 5128
rect 9826 5072 9831 5128
rect 3509 5070 9831 5072
rect 3509 5067 3575 5070
rect 9765 5067 9831 5070
rect 10685 5130 10751 5133
rect 14457 5130 14523 5133
rect 10685 5128 14523 5130
rect 10685 5072 10690 5128
rect 10746 5072 14462 5128
rect 14518 5072 14523 5128
rect 10685 5070 14523 5072
rect 10685 5067 10751 5070
rect 14457 5067 14523 5070
rect 7465 4994 7531 4997
rect 8661 4994 8727 4997
rect 9397 4996 9463 4997
rect 9397 4994 9444 4996
rect 7465 4992 8727 4994
rect 7465 4936 7470 4992
rect 7526 4936 8666 4992
rect 8722 4936 8727 4992
rect 7465 4934 8727 4936
rect 9352 4992 9444 4994
rect 9352 4936 9402 4992
rect 9352 4934 9444 4936
rect 7465 4931 7531 4934
rect 8661 4931 8727 4934
rect 9397 4932 9444 4934
rect 9508 4932 9514 4996
rect 9397 4931 9463 4932
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 10225 4858 10291 4861
rect 6318 4856 10291 4858
rect 6318 4800 10230 4856
rect 10286 4800 10291 4856
rect 6318 4798 10291 4800
rect 4705 4722 4771 4725
rect 6318 4722 6378 4798
rect 10225 4795 10291 4798
rect 4705 4720 6378 4722
rect 4705 4664 4710 4720
rect 4766 4664 6378 4720
rect 4705 4662 6378 4664
rect 9397 4722 9463 4725
rect 12934 4722 12940 4724
rect 9397 4720 12940 4722
rect 9397 4664 9402 4720
rect 9458 4664 12940 4720
rect 9397 4662 12940 4664
rect 4705 4659 4771 4662
rect 9397 4659 9463 4662
rect 12934 4660 12940 4662
rect 13004 4722 13010 4724
rect 13353 4722 13419 4725
rect 13004 4720 13419 4722
rect 13004 4664 13358 4720
rect 13414 4664 13419 4720
rect 13004 4662 13419 4664
rect 13004 4660 13010 4662
rect 13353 4659 13419 4662
rect 2129 4586 2195 4589
rect 13997 4586 14063 4589
rect 2129 4584 14063 4586
rect 2129 4528 2134 4584
rect 2190 4528 14002 4584
rect 14058 4528 14063 4584
rect 2129 4526 14063 4528
rect 2129 4523 2195 4526
rect 13997 4523 14063 4526
rect 0 4450 480 4480
rect 3233 4450 3299 4453
rect 0 4448 3299 4450
rect 0 4392 3238 4448
rect 3294 4392 3299 4448
rect 0 4390 3299 4392
rect 0 4360 480 4390
rect 3233 4387 3299 4390
rect 4337 4450 4403 4453
rect 8109 4450 8175 4453
rect 4337 4448 8175 4450
rect 4337 4392 4342 4448
rect 4398 4392 8114 4448
rect 8170 4392 8175 4448
rect 4337 4390 8175 4392
rect 4337 4387 4403 4390
rect 8109 4387 8175 4390
rect 9581 4450 9647 4453
rect 10542 4450 10548 4452
rect 9581 4448 10548 4450
rect 9581 4392 9586 4448
rect 9642 4392 10548 4448
rect 9581 4390 10548 4392
rect 9581 4387 9647 4390
rect 10542 4388 10548 4390
rect 10612 4450 10618 4452
rect 11421 4450 11487 4453
rect 10612 4448 11487 4450
rect 10612 4392 11426 4448
rect 11482 4392 11487 4448
rect 10612 4390 11487 4392
rect 10612 4388 10618 4390
rect 11421 4387 11487 4390
rect 3409 4384 3729 4385
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 4319 13590 4320
rect 5625 4314 5691 4317
rect 7281 4314 7347 4317
rect 11329 4316 11395 4317
rect 11278 4314 11284 4316
rect 5625 4312 7347 4314
rect 5625 4256 5630 4312
rect 5686 4256 7286 4312
rect 7342 4256 7347 4312
rect 5625 4254 7347 4256
rect 5625 4251 5691 4254
rect 7281 4251 7347 4254
rect 8940 4254 11284 4314
rect 11348 4312 11395 4316
rect 11390 4256 11395 4312
rect 5073 4178 5139 4181
rect 7925 4178 7991 4181
rect 8940 4178 9000 4254
rect 11278 4252 11284 4254
rect 11348 4252 11395 4256
rect 11329 4251 11395 4252
rect 5073 4176 9000 4178
rect 5073 4120 5078 4176
rect 5134 4120 7930 4176
rect 7986 4120 9000 4176
rect 5073 4118 9000 4120
rect 9121 4178 9187 4181
rect 9949 4178 10015 4181
rect 9121 4176 10015 4178
rect 9121 4120 9126 4176
rect 9182 4120 9954 4176
rect 10010 4120 10015 4176
rect 9121 4118 10015 4120
rect 5073 4115 5139 4118
rect 7925 4115 7991 4118
rect 9121 4115 9187 4118
rect 9949 4115 10015 4118
rect 10317 4178 10383 4181
rect 11830 4178 11836 4180
rect 10317 4176 11836 4178
rect 10317 4120 10322 4176
rect 10378 4120 11836 4176
rect 10317 4118 11836 4120
rect 10317 4115 10383 4118
rect 11830 4116 11836 4118
rect 11900 4116 11906 4180
rect 13353 4178 13419 4181
rect 15009 4178 15075 4181
rect 13353 4176 15075 4178
rect 13353 4120 13358 4176
rect 13414 4120 15014 4176
rect 15070 4120 15075 4176
rect 13353 4118 15075 4120
rect 13353 4115 13419 4118
rect 15009 4115 15075 4118
rect 2773 4042 2839 4045
rect 11881 4042 11947 4045
rect 2773 4040 11947 4042
rect 2773 3984 2778 4040
rect 2834 3984 11886 4040
rect 11942 3984 11947 4040
rect 2773 3982 11947 3984
rect 2773 3979 2839 3982
rect 11881 3979 11947 3982
rect 12341 4042 12407 4045
rect 14549 4042 14615 4045
rect 12341 4040 14615 4042
rect 12341 3984 12346 4040
rect 12402 3984 14554 4040
rect 14610 3984 14615 4040
rect 12341 3982 14615 3984
rect 12341 3979 12407 3982
rect 14549 3979 14615 3982
rect 8017 3906 8083 3909
rect 11237 3906 11303 3909
rect 13261 3906 13327 3909
rect 14457 3908 14523 3909
rect 8017 3904 10610 3906
rect 8017 3848 8022 3904
rect 8078 3848 10610 3904
rect 8017 3846 10610 3848
rect 8017 3843 8083 3846
rect 5874 3840 6194 3841
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 2221 3770 2287 3773
rect 5625 3770 5691 3773
rect 2221 3768 5691 3770
rect 2221 3712 2226 3768
rect 2282 3712 5630 3768
rect 5686 3712 5691 3768
rect 2221 3710 5691 3712
rect 2221 3707 2287 3710
rect 5625 3707 5691 3710
rect 7557 3770 7623 3773
rect 9438 3770 9444 3772
rect 7557 3768 9444 3770
rect 7557 3712 7562 3768
rect 7618 3712 9444 3768
rect 7557 3710 9444 3712
rect 7557 3707 7623 3710
rect 9438 3708 9444 3710
rect 9508 3708 9514 3772
rect 9765 3770 9831 3773
rect 10409 3770 10475 3773
rect 9765 3768 10475 3770
rect 9765 3712 9770 3768
rect 9826 3712 10414 3768
rect 10470 3712 10475 3768
rect 9765 3710 10475 3712
rect 9765 3707 9831 3710
rect 10409 3707 10475 3710
rect 10409 3634 10475 3637
rect 3144 3632 10475 3634
rect 3144 3576 10414 3632
rect 10470 3576 10475 3632
rect 3144 3574 10475 3576
rect 10550 3634 10610 3846
rect 11237 3904 13327 3906
rect 11237 3848 11242 3904
rect 11298 3848 13266 3904
rect 13322 3848 13327 3904
rect 11237 3846 13327 3848
rect 11237 3843 11303 3846
rect 13261 3843 13327 3846
rect 14406 3844 14412 3908
rect 14476 3906 14523 3908
rect 14476 3904 14568 3906
rect 14518 3848 14568 3904
rect 14476 3846 14568 3848
rect 14476 3844 14523 3846
rect 14457 3843 14523 3844
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 12382 3708 12388 3772
rect 12452 3770 12458 3772
rect 12452 3710 14842 3770
rect 12452 3708 12458 3710
rect 14641 3634 14707 3637
rect 10550 3632 14707 3634
rect 10550 3576 14646 3632
rect 14702 3576 14707 3632
rect 10550 3574 14707 3576
rect 0 3498 480 3528
rect 2957 3498 3023 3501
rect 0 3496 3023 3498
rect 0 3440 2962 3496
rect 3018 3440 3023 3496
rect 0 3438 3023 3440
rect 0 3408 480 3438
rect 2957 3435 3023 3438
rect 1761 3362 1827 3365
rect 3144 3362 3204 3574
rect 10409 3571 10475 3574
rect 14641 3571 14707 3574
rect 4613 3498 4679 3501
rect 5073 3498 5139 3501
rect 7649 3498 7715 3501
rect 14641 3498 14707 3501
rect 4613 3496 5139 3498
rect 4613 3440 4618 3496
rect 4674 3440 5078 3496
rect 5134 3440 5139 3496
rect 4613 3438 5139 3440
rect 4613 3435 4679 3438
rect 5073 3435 5139 3438
rect 5214 3496 7715 3498
rect 5214 3440 7654 3496
rect 7710 3440 7715 3496
rect 5214 3438 7715 3440
rect 1761 3360 3204 3362
rect 1761 3304 1766 3360
rect 1822 3304 3204 3360
rect 1761 3302 3204 3304
rect 4245 3362 4311 3365
rect 5214 3362 5274 3438
rect 7649 3435 7715 3438
rect 7974 3496 14707 3498
rect 7974 3440 14646 3496
rect 14702 3440 14707 3496
rect 7974 3438 14707 3440
rect 4245 3360 5274 3362
rect 4245 3304 4250 3360
rect 4306 3304 5274 3360
rect 4245 3302 5274 3304
rect 6821 3362 6887 3365
rect 7974 3362 8034 3438
rect 14641 3435 14707 3438
rect 6821 3360 8034 3362
rect 6821 3304 6826 3360
rect 6882 3304 8034 3360
rect 6821 3302 8034 3304
rect 8937 3362 9003 3365
rect 12433 3362 12499 3365
rect 8937 3360 12499 3362
rect 8937 3304 8942 3360
rect 8998 3304 12438 3360
rect 12494 3304 12499 3360
rect 8937 3302 12499 3304
rect 14782 3362 14842 3710
rect 16520 3362 17000 3392
rect 14782 3302 17000 3362
rect 1761 3299 1827 3302
rect 4245 3299 4311 3302
rect 6821 3299 6887 3302
rect 8937 3299 9003 3302
rect 12433 3299 12499 3302
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 16520 3272 17000 3302
rect 13270 3231 13590 3232
rect 4337 3226 4403 3229
rect 7833 3226 7899 3229
rect 10409 3228 10475 3229
rect 4337 3224 7899 3226
rect 4337 3168 4342 3224
rect 4398 3168 7838 3224
rect 7894 3168 7899 3224
rect 4337 3166 7899 3168
rect 4337 3163 4403 3166
rect 7833 3163 7899 3166
rect 10358 3164 10364 3228
rect 10428 3226 10475 3228
rect 10428 3224 10520 3226
rect 10470 3168 10520 3224
rect 10428 3166 10520 3168
rect 10428 3164 10475 3166
rect 11646 3164 11652 3228
rect 11716 3226 11722 3228
rect 12341 3226 12407 3229
rect 11716 3224 12407 3226
rect 11716 3168 12346 3224
rect 12402 3168 12407 3224
rect 11716 3166 12407 3168
rect 11716 3164 11722 3166
rect 10409 3163 10475 3164
rect 12341 3163 12407 3166
rect 12617 3226 12683 3229
rect 12750 3226 12756 3228
rect 12617 3224 12756 3226
rect 12617 3168 12622 3224
rect 12678 3168 12756 3224
rect 12617 3166 12756 3168
rect 12617 3163 12683 3166
rect 12750 3164 12756 3166
rect 12820 3164 12826 3228
rect 1117 3090 1183 3093
rect 15009 3090 15075 3093
rect 1117 3088 15075 3090
rect 1117 3032 1122 3088
rect 1178 3032 15014 3088
rect 15070 3032 15075 3088
rect 1117 3030 15075 3032
rect 1117 3027 1183 3030
rect 15009 3027 15075 3030
rect 1853 2954 1919 2957
rect 16757 2954 16823 2957
rect 1853 2952 16823 2954
rect 1853 2896 1858 2952
rect 1914 2896 16762 2952
rect 16818 2896 16823 2952
rect 1853 2894 16823 2896
rect 1853 2891 1919 2894
rect 16757 2891 16823 2894
rect 5073 2818 5139 2821
rect 5030 2816 5139 2818
rect 5030 2760 5078 2816
rect 5134 2760 5139 2816
rect 5030 2755 5139 2760
rect 7557 2818 7623 2821
rect 8017 2818 8083 2821
rect 7557 2816 8083 2818
rect 7557 2760 7562 2816
rect 7618 2760 8022 2816
rect 8078 2760 8083 2816
rect 7557 2758 8083 2760
rect 7557 2755 7623 2758
rect 8017 2755 8083 2758
rect 8569 2818 8635 2821
rect 9213 2820 9279 2821
rect 9949 2820 10015 2821
rect 9070 2818 9076 2820
rect 8569 2816 9076 2818
rect 8569 2760 8574 2816
rect 8630 2760 9076 2816
rect 8569 2758 9076 2760
rect 8569 2755 8635 2758
rect 9070 2756 9076 2758
rect 9140 2756 9146 2820
rect 9213 2816 9260 2820
rect 9324 2818 9330 2820
rect 9213 2760 9218 2816
rect 9213 2756 9260 2760
rect 9324 2758 9370 2818
rect 9949 2816 9996 2820
rect 10060 2818 10066 2820
rect 11513 2818 11579 2821
rect 13118 2818 13124 2820
rect 9949 2760 9954 2816
rect 9324 2756 9330 2758
rect 9949 2756 9996 2760
rect 10060 2758 10106 2818
rect 11513 2816 13124 2818
rect 11513 2760 11518 2816
rect 11574 2760 13124 2816
rect 11513 2758 13124 2760
rect 10060 2756 10066 2758
rect 9213 2755 9279 2756
rect 9949 2755 10015 2756
rect 11513 2755 11579 2758
rect 13118 2756 13124 2758
rect 13188 2818 13194 2820
rect 13905 2818 13971 2821
rect 13188 2816 13971 2818
rect 13188 2760 13910 2816
rect 13966 2760 13971 2816
rect 13188 2758 13971 2760
rect 13188 2756 13194 2758
rect 13905 2755 13971 2758
rect 5030 2546 5090 2755
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 8937 2682 9003 2685
rect 9581 2682 9647 2685
rect 8937 2680 9647 2682
rect 8937 2624 8942 2680
rect 8998 2624 9586 2680
rect 9642 2624 9647 2680
rect 8937 2622 9647 2624
rect 8937 2619 9003 2622
rect 9581 2619 9647 2622
rect 9857 2682 9923 2685
rect 10174 2682 10180 2684
rect 9857 2680 10180 2682
rect 9857 2624 9862 2680
rect 9918 2624 10180 2680
rect 9857 2622 10180 2624
rect 9857 2619 9923 2622
rect 10174 2620 10180 2622
rect 10244 2620 10250 2684
rect 12525 2682 12591 2685
rect 12985 2682 13051 2685
rect 12525 2680 13051 2682
rect 12525 2624 12530 2680
rect 12586 2624 12990 2680
rect 13046 2624 13051 2680
rect 12525 2622 13051 2624
rect 12525 2619 12591 2622
rect 12985 2619 13051 2622
rect 7557 2546 7623 2549
rect 5030 2544 7623 2546
rect 5030 2488 7562 2544
rect 7618 2488 7623 2544
rect 5030 2486 7623 2488
rect 7557 2483 7623 2486
rect 7833 2546 7899 2549
rect 12525 2546 12591 2549
rect 7833 2544 12591 2546
rect 7833 2488 7838 2544
rect 7894 2488 12530 2544
rect 12586 2488 12591 2544
rect 7833 2486 12591 2488
rect 7833 2483 7899 2486
rect 12525 2483 12591 2486
rect 0 2410 480 2440
rect 4061 2410 4127 2413
rect 0 2408 4127 2410
rect 0 2352 4066 2408
rect 4122 2352 4127 2408
rect 0 2350 4127 2352
rect 0 2320 480 2350
rect 4061 2347 4127 2350
rect 9581 2410 9647 2413
rect 9806 2410 9812 2412
rect 9581 2408 9812 2410
rect 9581 2352 9586 2408
rect 9642 2352 9812 2408
rect 9581 2350 9812 2352
rect 9581 2347 9647 2350
rect 9806 2348 9812 2350
rect 9876 2410 9882 2412
rect 13261 2410 13327 2413
rect 14038 2410 14044 2412
rect 9876 2408 14044 2410
rect 9876 2352 13266 2408
rect 13322 2352 14044 2408
rect 9876 2350 14044 2352
rect 9876 2348 9882 2350
rect 13261 2347 13327 2350
rect 14038 2348 14044 2350
rect 14108 2348 14114 2412
rect 9438 2212 9444 2276
rect 9508 2274 9514 2276
rect 9581 2274 9647 2277
rect 9508 2272 9647 2274
rect 9508 2216 9586 2272
rect 9642 2216 9647 2272
rect 9508 2214 9647 2216
rect 9508 2212 9514 2214
rect 9581 2211 9647 2214
rect 10961 2274 11027 2277
rect 12198 2274 12204 2276
rect 10961 2272 12204 2274
rect 10961 2216 10966 2272
rect 11022 2216 12204 2272
rect 10961 2214 12204 2216
rect 10961 2211 11027 2214
rect 12198 2212 12204 2214
rect 12268 2212 12274 2276
rect 3409 2208 3729 2209
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
rect 0 1458 480 1488
rect 1945 1458 2011 1461
rect 0 1456 2011 1458
rect 0 1400 1950 1456
rect 2006 1400 2011 1456
rect 0 1398 2011 1400
rect 0 1368 480 1398
rect 1945 1395 2011 1398
rect 0 506 480 536
rect 2865 506 2931 509
rect 0 504 2931 506
rect 0 448 2870 504
rect 2926 448 2931 504
rect 0 446 2931 448
rect 0 416 480 446
rect 2865 443 2931 446
<< via3 >>
rect 3417 17436 3481 17440
rect 3417 17380 3421 17436
rect 3421 17380 3477 17436
rect 3477 17380 3481 17436
rect 3417 17376 3481 17380
rect 3497 17436 3561 17440
rect 3497 17380 3501 17436
rect 3501 17380 3557 17436
rect 3557 17380 3561 17436
rect 3497 17376 3561 17380
rect 3577 17436 3641 17440
rect 3577 17380 3581 17436
rect 3581 17380 3637 17436
rect 3637 17380 3641 17436
rect 3577 17376 3641 17380
rect 3657 17436 3721 17440
rect 3657 17380 3661 17436
rect 3661 17380 3717 17436
rect 3717 17380 3721 17436
rect 3657 17376 3721 17380
rect 8348 17436 8412 17440
rect 8348 17380 8352 17436
rect 8352 17380 8408 17436
rect 8408 17380 8412 17436
rect 8348 17376 8412 17380
rect 8428 17436 8492 17440
rect 8428 17380 8432 17436
rect 8432 17380 8488 17436
rect 8488 17380 8492 17436
rect 8428 17376 8492 17380
rect 8508 17436 8572 17440
rect 8508 17380 8512 17436
rect 8512 17380 8568 17436
rect 8568 17380 8572 17436
rect 8508 17376 8572 17380
rect 8588 17436 8652 17440
rect 8588 17380 8592 17436
rect 8592 17380 8648 17436
rect 8648 17380 8652 17436
rect 8588 17376 8652 17380
rect 13278 17436 13342 17440
rect 13278 17380 13282 17436
rect 13282 17380 13338 17436
rect 13338 17380 13342 17436
rect 13278 17376 13342 17380
rect 13358 17436 13422 17440
rect 13358 17380 13362 17436
rect 13362 17380 13418 17436
rect 13418 17380 13422 17436
rect 13358 17376 13422 17380
rect 13438 17436 13502 17440
rect 13438 17380 13442 17436
rect 13442 17380 13498 17436
rect 13498 17380 13502 17436
rect 13438 17376 13502 17380
rect 13518 17436 13582 17440
rect 13518 17380 13522 17436
rect 13522 17380 13578 17436
rect 13578 17380 13582 17436
rect 13518 17376 13582 17380
rect 9628 17172 9692 17236
rect 10180 17036 10244 17100
rect 3188 16900 3252 16964
rect 5882 16892 5946 16896
rect 5882 16836 5886 16892
rect 5886 16836 5942 16892
rect 5942 16836 5946 16892
rect 5882 16832 5946 16836
rect 5962 16892 6026 16896
rect 5962 16836 5966 16892
rect 5966 16836 6022 16892
rect 6022 16836 6026 16892
rect 5962 16832 6026 16836
rect 6042 16892 6106 16896
rect 6042 16836 6046 16892
rect 6046 16836 6102 16892
rect 6102 16836 6106 16892
rect 6042 16832 6106 16836
rect 6122 16892 6186 16896
rect 6122 16836 6126 16892
rect 6126 16836 6182 16892
rect 6182 16836 6186 16892
rect 6122 16832 6186 16836
rect 10813 16892 10877 16896
rect 10813 16836 10817 16892
rect 10817 16836 10873 16892
rect 10873 16836 10877 16892
rect 10813 16832 10877 16836
rect 10893 16892 10957 16896
rect 10893 16836 10897 16892
rect 10897 16836 10953 16892
rect 10953 16836 10957 16892
rect 10893 16832 10957 16836
rect 10973 16892 11037 16896
rect 10973 16836 10977 16892
rect 10977 16836 11033 16892
rect 11033 16836 11037 16892
rect 10973 16832 11037 16836
rect 11053 16892 11117 16896
rect 11053 16836 11057 16892
rect 11057 16836 11113 16892
rect 11113 16836 11117 16892
rect 11053 16832 11117 16836
rect 9812 16764 9876 16828
rect 10364 16628 10428 16692
rect 13676 16628 13740 16692
rect 12572 16552 12636 16556
rect 12572 16496 12586 16552
rect 12586 16496 12636 16552
rect 12572 16492 12636 16496
rect 9996 16356 10060 16420
rect 3417 16348 3481 16352
rect 3417 16292 3421 16348
rect 3421 16292 3477 16348
rect 3477 16292 3481 16348
rect 3417 16288 3481 16292
rect 3497 16348 3561 16352
rect 3497 16292 3501 16348
rect 3501 16292 3557 16348
rect 3557 16292 3561 16348
rect 3497 16288 3561 16292
rect 3577 16348 3641 16352
rect 3577 16292 3581 16348
rect 3581 16292 3637 16348
rect 3637 16292 3641 16348
rect 3577 16288 3641 16292
rect 3657 16348 3721 16352
rect 3657 16292 3661 16348
rect 3661 16292 3717 16348
rect 3717 16292 3721 16348
rect 3657 16288 3721 16292
rect 8348 16348 8412 16352
rect 8348 16292 8352 16348
rect 8352 16292 8408 16348
rect 8408 16292 8412 16348
rect 8348 16288 8412 16292
rect 8428 16348 8492 16352
rect 8428 16292 8432 16348
rect 8432 16292 8488 16348
rect 8488 16292 8492 16348
rect 8428 16288 8492 16292
rect 8508 16348 8572 16352
rect 8508 16292 8512 16348
rect 8512 16292 8568 16348
rect 8568 16292 8572 16348
rect 8508 16288 8572 16292
rect 8588 16348 8652 16352
rect 8588 16292 8592 16348
rect 8592 16292 8648 16348
rect 8648 16292 8652 16348
rect 8588 16288 8652 16292
rect 13278 16348 13342 16352
rect 13278 16292 13282 16348
rect 13282 16292 13338 16348
rect 13338 16292 13342 16348
rect 13278 16288 13342 16292
rect 13358 16348 13422 16352
rect 13358 16292 13362 16348
rect 13362 16292 13418 16348
rect 13418 16292 13422 16348
rect 13358 16288 13422 16292
rect 13438 16348 13502 16352
rect 13438 16292 13442 16348
rect 13442 16292 13498 16348
rect 13498 16292 13502 16348
rect 13438 16288 13502 16292
rect 13518 16348 13582 16352
rect 13518 16292 13522 16348
rect 13522 16292 13578 16348
rect 13578 16292 13582 16348
rect 13518 16288 13582 16292
rect 12572 16220 12636 16284
rect 5882 15804 5946 15808
rect 5882 15748 5886 15804
rect 5886 15748 5942 15804
rect 5942 15748 5946 15804
rect 5882 15744 5946 15748
rect 5962 15804 6026 15808
rect 5962 15748 5966 15804
rect 5966 15748 6022 15804
rect 6022 15748 6026 15804
rect 5962 15744 6026 15748
rect 6042 15804 6106 15808
rect 6042 15748 6046 15804
rect 6046 15748 6102 15804
rect 6102 15748 6106 15804
rect 6042 15744 6106 15748
rect 6122 15804 6186 15808
rect 6122 15748 6126 15804
rect 6126 15748 6182 15804
rect 6182 15748 6186 15804
rect 6122 15744 6186 15748
rect 10813 15804 10877 15808
rect 10813 15748 10817 15804
rect 10817 15748 10873 15804
rect 10873 15748 10877 15804
rect 10813 15744 10877 15748
rect 10893 15804 10957 15808
rect 10893 15748 10897 15804
rect 10897 15748 10953 15804
rect 10953 15748 10957 15804
rect 10893 15744 10957 15748
rect 10973 15804 11037 15808
rect 10973 15748 10977 15804
rect 10977 15748 11033 15804
rect 11033 15748 11037 15804
rect 10973 15744 11037 15748
rect 11053 15804 11117 15808
rect 11053 15748 11057 15804
rect 11057 15748 11113 15804
rect 11113 15748 11117 15804
rect 11053 15744 11117 15748
rect 9444 15736 9508 15740
rect 9444 15680 9458 15736
rect 9458 15680 9508 15736
rect 9444 15676 9508 15680
rect 12204 15676 12268 15740
rect 12388 15540 12452 15604
rect 10548 15328 10612 15332
rect 10548 15272 10562 15328
rect 10562 15272 10612 15328
rect 10548 15268 10612 15272
rect 3417 15260 3481 15264
rect 3417 15204 3421 15260
rect 3421 15204 3477 15260
rect 3477 15204 3481 15260
rect 3417 15200 3481 15204
rect 3497 15260 3561 15264
rect 3497 15204 3501 15260
rect 3501 15204 3557 15260
rect 3557 15204 3561 15260
rect 3497 15200 3561 15204
rect 3577 15260 3641 15264
rect 3577 15204 3581 15260
rect 3581 15204 3637 15260
rect 3637 15204 3641 15260
rect 3577 15200 3641 15204
rect 3657 15260 3721 15264
rect 3657 15204 3661 15260
rect 3661 15204 3717 15260
rect 3717 15204 3721 15260
rect 3657 15200 3721 15204
rect 8348 15260 8412 15264
rect 8348 15204 8352 15260
rect 8352 15204 8408 15260
rect 8408 15204 8412 15260
rect 8348 15200 8412 15204
rect 8428 15260 8492 15264
rect 8428 15204 8432 15260
rect 8432 15204 8488 15260
rect 8488 15204 8492 15260
rect 8428 15200 8492 15204
rect 8508 15260 8572 15264
rect 8508 15204 8512 15260
rect 8512 15204 8568 15260
rect 8568 15204 8572 15260
rect 8508 15200 8572 15204
rect 8588 15260 8652 15264
rect 8588 15204 8592 15260
rect 8592 15204 8648 15260
rect 8648 15204 8652 15260
rect 8588 15200 8652 15204
rect 13278 15260 13342 15264
rect 13278 15204 13282 15260
rect 13282 15204 13338 15260
rect 13338 15204 13342 15260
rect 13278 15200 13342 15204
rect 13358 15260 13422 15264
rect 13358 15204 13362 15260
rect 13362 15204 13418 15260
rect 13418 15204 13422 15260
rect 13358 15200 13422 15204
rect 13438 15260 13502 15264
rect 13438 15204 13442 15260
rect 13442 15204 13498 15260
rect 13498 15204 13502 15260
rect 13438 15200 13502 15204
rect 13518 15260 13582 15264
rect 13518 15204 13522 15260
rect 13522 15204 13578 15260
rect 13578 15204 13582 15260
rect 13518 15200 13582 15204
rect 9260 15132 9324 15196
rect 12756 14996 12820 15060
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 6122 14716 6186 14720
rect 6122 14660 6126 14716
rect 6126 14660 6182 14716
rect 6182 14660 6186 14716
rect 6122 14656 6186 14660
rect 10813 14716 10877 14720
rect 10813 14660 10817 14716
rect 10817 14660 10873 14716
rect 10873 14660 10877 14716
rect 10813 14656 10877 14660
rect 10893 14716 10957 14720
rect 10893 14660 10897 14716
rect 10897 14660 10953 14716
rect 10953 14660 10957 14716
rect 10893 14656 10957 14660
rect 10973 14716 11037 14720
rect 10973 14660 10977 14716
rect 10977 14660 11033 14716
rect 11033 14660 11037 14716
rect 10973 14656 11037 14660
rect 11053 14716 11117 14720
rect 11053 14660 11057 14716
rect 11057 14660 11113 14716
rect 11113 14660 11117 14716
rect 11053 14656 11117 14660
rect 8892 14588 8956 14652
rect 9628 14588 9692 14652
rect 12940 14588 13004 14652
rect 9076 14452 9140 14516
rect 9628 14452 9692 14516
rect 11284 14512 11348 14516
rect 11284 14456 11334 14512
rect 11334 14456 11348 14512
rect 11284 14452 11348 14456
rect 11468 14180 11532 14244
rect 3417 14172 3481 14176
rect 3417 14116 3421 14172
rect 3421 14116 3477 14172
rect 3477 14116 3481 14172
rect 3417 14112 3481 14116
rect 3497 14172 3561 14176
rect 3497 14116 3501 14172
rect 3501 14116 3557 14172
rect 3557 14116 3561 14172
rect 3497 14112 3561 14116
rect 3577 14172 3641 14176
rect 3577 14116 3581 14172
rect 3581 14116 3637 14172
rect 3637 14116 3641 14172
rect 3577 14112 3641 14116
rect 3657 14172 3721 14176
rect 3657 14116 3661 14172
rect 3661 14116 3717 14172
rect 3717 14116 3721 14172
rect 3657 14112 3721 14116
rect 8348 14172 8412 14176
rect 8348 14116 8352 14172
rect 8352 14116 8408 14172
rect 8408 14116 8412 14172
rect 8348 14112 8412 14116
rect 8428 14172 8492 14176
rect 8428 14116 8432 14172
rect 8432 14116 8488 14172
rect 8488 14116 8492 14172
rect 8428 14112 8492 14116
rect 8508 14172 8572 14176
rect 8508 14116 8512 14172
rect 8512 14116 8568 14172
rect 8568 14116 8572 14172
rect 8508 14112 8572 14116
rect 8588 14172 8652 14176
rect 8588 14116 8592 14172
rect 8592 14116 8648 14172
rect 8648 14116 8652 14172
rect 8588 14112 8652 14116
rect 13278 14172 13342 14176
rect 13278 14116 13282 14172
rect 13282 14116 13338 14172
rect 13338 14116 13342 14172
rect 13278 14112 13342 14116
rect 13358 14172 13422 14176
rect 13358 14116 13362 14172
rect 13362 14116 13418 14172
rect 13418 14116 13422 14172
rect 13358 14112 13422 14116
rect 13438 14172 13502 14176
rect 13438 14116 13442 14172
rect 13442 14116 13498 14172
rect 13498 14116 13502 14172
rect 13438 14112 13502 14116
rect 13518 14172 13582 14176
rect 13518 14116 13522 14172
rect 13522 14116 13578 14172
rect 13578 14116 13582 14172
rect 13518 14112 13582 14116
rect 9076 14044 9140 14108
rect 12020 14044 12084 14108
rect 9444 13636 9508 13700
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 6122 13628 6186 13632
rect 6122 13572 6126 13628
rect 6126 13572 6182 13628
rect 6182 13572 6186 13628
rect 6122 13568 6186 13572
rect 10813 13628 10877 13632
rect 10813 13572 10817 13628
rect 10817 13572 10873 13628
rect 10873 13572 10877 13628
rect 10813 13568 10877 13572
rect 10893 13628 10957 13632
rect 10893 13572 10897 13628
rect 10897 13572 10953 13628
rect 10953 13572 10957 13628
rect 10893 13568 10957 13572
rect 10973 13628 11037 13632
rect 10973 13572 10977 13628
rect 10977 13572 11033 13628
rect 11033 13572 11037 13628
rect 10973 13568 11037 13572
rect 11053 13628 11117 13632
rect 11053 13572 11057 13628
rect 11057 13572 11113 13628
rect 11113 13572 11117 13628
rect 11053 13568 11117 13572
rect 9260 13500 9324 13564
rect 9444 13500 9508 13564
rect 9996 13500 10060 13564
rect 11652 13500 11716 13564
rect 9076 13228 9140 13292
rect 3417 13084 3481 13088
rect 3417 13028 3421 13084
rect 3421 13028 3477 13084
rect 3477 13028 3481 13084
rect 3417 13024 3481 13028
rect 3497 13084 3561 13088
rect 3497 13028 3501 13084
rect 3501 13028 3557 13084
rect 3557 13028 3561 13084
rect 3497 13024 3561 13028
rect 3577 13084 3641 13088
rect 3577 13028 3581 13084
rect 3581 13028 3637 13084
rect 3637 13028 3641 13084
rect 3577 13024 3641 13028
rect 3657 13084 3721 13088
rect 3657 13028 3661 13084
rect 3661 13028 3717 13084
rect 3717 13028 3721 13084
rect 3657 13024 3721 13028
rect 8348 13084 8412 13088
rect 8348 13028 8352 13084
rect 8352 13028 8408 13084
rect 8408 13028 8412 13084
rect 8348 13024 8412 13028
rect 8428 13084 8492 13088
rect 8428 13028 8432 13084
rect 8432 13028 8488 13084
rect 8488 13028 8492 13084
rect 8428 13024 8492 13028
rect 8508 13084 8572 13088
rect 8508 13028 8512 13084
rect 8512 13028 8568 13084
rect 8568 13028 8572 13084
rect 8508 13024 8572 13028
rect 8588 13084 8652 13088
rect 8588 13028 8592 13084
rect 8592 13028 8648 13084
rect 8648 13028 8652 13084
rect 8588 13024 8652 13028
rect 6684 12820 6748 12884
rect 13676 13152 13740 13156
rect 13676 13096 13726 13152
rect 13726 13096 13740 13152
rect 13676 13092 13740 13096
rect 13278 13084 13342 13088
rect 13278 13028 13282 13084
rect 13282 13028 13338 13084
rect 13338 13028 13342 13084
rect 13278 13024 13342 13028
rect 13358 13084 13422 13088
rect 13358 13028 13362 13084
rect 13362 13028 13418 13084
rect 13418 13028 13422 13084
rect 13358 13024 13422 13028
rect 13438 13084 13502 13088
rect 13438 13028 13442 13084
rect 13442 13028 13498 13084
rect 13498 13028 13502 13084
rect 13438 13024 13502 13028
rect 13518 13084 13582 13088
rect 13518 13028 13522 13084
rect 13522 13028 13578 13084
rect 13578 13028 13582 13084
rect 13518 13024 13582 13028
rect 10180 12820 10244 12884
rect 11836 12880 11900 12884
rect 11836 12824 11850 12880
rect 11850 12824 11900 12880
rect 11836 12820 11900 12824
rect 12020 12820 12084 12884
rect 12020 12548 12084 12612
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 6122 12540 6186 12544
rect 6122 12484 6126 12540
rect 6126 12484 6182 12540
rect 6182 12484 6186 12540
rect 6122 12480 6186 12484
rect 10813 12540 10877 12544
rect 10813 12484 10817 12540
rect 10817 12484 10873 12540
rect 10873 12484 10877 12540
rect 10813 12480 10877 12484
rect 10893 12540 10957 12544
rect 10893 12484 10897 12540
rect 10897 12484 10953 12540
rect 10953 12484 10957 12540
rect 10893 12480 10957 12484
rect 10973 12540 11037 12544
rect 10973 12484 10977 12540
rect 10977 12484 11033 12540
rect 11033 12484 11037 12540
rect 10973 12480 11037 12484
rect 11053 12540 11117 12544
rect 11053 12484 11057 12540
rect 11057 12484 11113 12540
rect 11113 12484 11117 12540
rect 11053 12480 11117 12484
rect 11468 12412 11532 12476
rect 9812 12276 9876 12340
rect 13676 12276 13740 12340
rect 9812 12140 9876 12204
rect 10180 12004 10244 12068
rect 3417 11996 3481 12000
rect 3417 11940 3421 11996
rect 3421 11940 3477 11996
rect 3477 11940 3481 11996
rect 3417 11936 3481 11940
rect 3497 11996 3561 12000
rect 3497 11940 3501 11996
rect 3501 11940 3557 11996
rect 3557 11940 3561 11996
rect 3497 11936 3561 11940
rect 3577 11996 3641 12000
rect 3577 11940 3581 11996
rect 3581 11940 3637 11996
rect 3637 11940 3641 11996
rect 3577 11936 3641 11940
rect 3657 11996 3721 12000
rect 3657 11940 3661 11996
rect 3661 11940 3717 11996
rect 3717 11940 3721 11996
rect 3657 11936 3721 11940
rect 8348 11996 8412 12000
rect 8348 11940 8352 11996
rect 8352 11940 8408 11996
rect 8408 11940 8412 11996
rect 8348 11936 8412 11940
rect 8428 11996 8492 12000
rect 8428 11940 8432 11996
rect 8432 11940 8488 11996
rect 8488 11940 8492 11996
rect 8428 11936 8492 11940
rect 8508 11996 8572 12000
rect 8508 11940 8512 11996
rect 8512 11940 8568 11996
rect 8568 11940 8572 11996
rect 8508 11936 8572 11940
rect 8588 11996 8652 12000
rect 8588 11940 8592 11996
rect 8592 11940 8648 11996
rect 8648 11940 8652 11996
rect 8588 11936 8652 11940
rect 13278 11996 13342 12000
rect 13278 11940 13282 11996
rect 13282 11940 13338 11996
rect 13338 11940 13342 11996
rect 13278 11936 13342 11940
rect 13358 11996 13422 12000
rect 13358 11940 13362 11996
rect 13362 11940 13418 11996
rect 13418 11940 13422 11996
rect 13358 11936 13422 11940
rect 13438 11996 13502 12000
rect 13438 11940 13442 11996
rect 13442 11940 13498 11996
rect 13498 11940 13502 11996
rect 13438 11936 13502 11940
rect 13518 11996 13582 12000
rect 13518 11940 13522 11996
rect 13522 11940 13578 11996
rect 13578 11940 13582 11996
rect 13518 11936 13582 11940
rect 11284 11868 11348 11932
rect 10548 11732 10612 11796
rect 13124 11732 13188 11796
rect 8892 11460 8956 11524
rect 9628 11460 9692 11524
rect 12388 11460 12452 11524
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 6122 11452 6186 11456
rect 6122 11396 6126 11452
rect 6126 11396 6182 11452
rect 6182 11396 6186 11452
rect 6122 11392 6186 11396
rect 10813 11452 10877 11456
rect 10813 11396 10817 11452
rect 10817 11396 10873 11452
rect 10873 11396 10877 11452
rect 10813 11392 10877 11396
rect 10893 11452 10957 11456
rect 10893 11396 10897 11452
rect 10897 11396 10953 11452
rect 10953 11396 10957 11452
rect 10893 11392 10957 11396
rect 10973 11452 11037 11456
rect 10973 11396 10977 11452
rect 10977 11396 11033 11452
rect 11033 11396 11037 11452
rect 10973 11392 11037 11396
rect 11053 11452 11117 11456
rect 11053 11396 11057 11452
rect 11057 11396 11113 11452
rect 11113 11396 11117 11452
rect 11053 11392 11117 11396
rect 9444 11188 9508 11252
rect 11468 11188 11532 11252
rect 12020 11188 12084 11252
rect 12388 11188 12452 11252
rect 11468 10916 11532 10980
rect 12020 10916 12084 10980
rect 3417 10908 3481 10912
rect 3417 10852 3421 10908
rect 3421 10852 3477 10908
rect 3477 10852 3481 10908
rect 3417 10848 3481 10852
rect 3497 10908 3561 10912
rect 3497 10852 3501 10908
rect 3501 10852 3557 10908
rect 3557 10852 3561 10908
rect 3497 10848 3561 10852
rect 3577 10908 3641 10912
rect 3577 10852 3581 10908
rect 3581 10852 3637 10908
rect 3637 10852 3641 10908
rect 3577 10848 3641 10852
rect 3657 10908 3721 10912
rect 3657 10852 3661 10908
rect 3661 10852 3717 10908
rect 3717 10852 3721 10908
rect 3657 10848 3721 10852
rect 8348 10908 8412 10912
rect 8348 10852 8352 10908
rect 8352 10852 8408 10908
rect 8408 10852 8412 10908
rect 8348 10848 8412 10852
rect 8428 10908 8492 10912
rect 8428 10852 8432 10908
rect 8432 10852 8488 10908
rect 8488 10852 8492 10908
rect 8428 10848 8492 10852
rect 8508 10908 8572 10912
rect 8508 10852 8512 10908
rect 8512 10852 8568 10908
rect 8568 10852 8572 10908
rect 8508 10848 8572 10852
rect 8588 10908 8652 10912
rect 8588 10852 8592 10908
rect 8592 10852 8648 10908
rect 8648 10852 8652 10908
rect 8588 10848 8652 10852
rect 13278 10908 13342 10912
rect 13278 10852 13282 10908
rect 13282 10852 13338 10908
rect 13338 10852 13342 10908
rect 13278 10848 13342 10852
rect 13358 10908 13422 10912
rect 13358 10852 13362 10908
rect 13362 10852 13418 10908
rect 13418 10852 13422 10908
rect 13358 10848 13422 10852
rect 13438 10908 13502 10912
rect 13438 10852 13442 10908
rect 13442 10852 13498 10908
rect 13498 10852 13502 10908
rect 13438 10848 13502 10852
rect 13518 10908 13582 10912
rect 13518 10852 13522 10908
rect 13522 10852 13578 10908
rect 13578 10852 13582 10908
rect 13518 10848 13582 10852
rect 9996 10780 10060 10844
rect 11468 10780 11532 10844
rect 11836 10780 11900 10844
rect 9444 10644 9508 10708
rect 3188 10372 3252 10436
rect 11836 10372 11900 10436
rect 12388 10372 12452 10436
rect 12940 10372 13004 10436
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 6122 10364 6186 10368
rect 6122 10308 6126 10364
rect 6126 10308 6182 10364
rect 6182 10308 6186 10364
rect 6122 10304 6186 10308
rect 10813 10364 10877 10368
rect 10813 10308 10817 10364
rect 10817 10308 10873 10364
rect 10873 10308 10877 10364
rect 10813 10304 10877 10308
rect 10893 10364 10957 10368
rect 10893 10308 10897 10364
rect 10897 10308 10953 10364
rect 10953 10308 10957 10364
rect 10893 10304 10957 10308
rect 10973 10364 11037 10368
rect 10973 10308 10977 10364
rect 10977 10308 11033 10364
rect 11033 10308 11037 10364
rect 10973 10304 11037 10308
rect 11053 10364 11117 10368
rect 11053 10308 11057 10364
rect 11057 10308 11113 10364
rect 11113 10308 11117 10364
rect 11053 10304 11117 10308
rect 12756 10100 12820 10164
rect 13676 10160 13740 10164
rect 13676 10104 13726 10160
rect 13726 10104 13740 10160
rect 13676 10100 13740 10104
rect 11652 9888 11716 9892
rect 11652 9832 11702 9888
rect 11702 9832 11716 9888
rect 11652 9828 11716 9832
rect 12204 9828 12268 9892
rect 3417 9820 3481 9824
rect 3417 9764 3421 9820
rect 3421 9764 3477 9820
rect 3477 9764 3481 9820
rect 3417 9760 3481 9764
rect 3497 9820 3561 9824
rect 3497 9764 3501 9820
rect 3501 9764 3557 9820
rect 3557 9764 3561 9820
rect 3497 9760 3561 9764
rect 3577 9820 3641 9824
rect 3577 9764 3581 9820
rect 3581 9764 3637 9820
rect 3637 9764 3641 9820
rect 3577 9760 3641 9764
rect 3657 9820 3721 9824
rect 3657 9764 3661 9820
rect 3661 9764 3717 9820
rect 3717 9764 3721 9820
rect 3657 9760 3721 9764
rect 8348 9820 8412 9824
rect 8348 9764 8352 9820
rect 8352 9764 8408 9820
rect 8408 9764 8412 9820
rect 8348 9760 8412 9764
rect 8428 9820 8492 9824
rect 8428 9764 8432 9820
rect 8432 9764 8488 9820
rect 8488 9764 8492 9820
rect 8428 9760 8492 9764
rect 8508 9820 8572 9824
rect 8508 9764 8512 9820
rect 8512 9764 8568 9820
rect 8568 9764 8572 9820
rect 8508 9760 8572 9764
rect 8588 9820 8652 9824
rect 8588 9764 8592 9820
rect 8592 9764 8648 9820
rect 8648 9764 8652 9820
rect 8588 9760 8652 9764
rect 13278 9820 13342 9824
rect 13278 9764 13282 9820
rect 13282 9764 13338 9820
rect 13338 9764 13342 9820
rect 13278 9760 13342 9764
rect 13358 9820 13422 9824
rect 13358 9764 13362 9820
rect 13362 9764 13418 9820
rect 13418 9764 13422 9820
rect 13358 9760 13422 9764
rect 13438 9820 13502 9824
rect 13438 9764 13442 9820
rect 13442 9764 13498 9820
rect 13498 9764 13502 9820
rect 13438 9760 13502 9764
rect 13518 9820 13582 9824
rect 13518 9764 13522 9820
rect 13522 9764 13578 9820
rect 13578 9764 13582 9820
rect 13518 9760 13582 9764
rect 9076 9692 9140 9756
rect 9996 9692 10060 9756
rect 12204 9420 12268 9484
rect 9444 9344 9508 9348
rect 9444 9288 9494 9344
rect 9494 9288 9508 9344
rect 9444 9284 9508 9288
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 6122 9276 6186 9280
rect 6122 9220 6126 9276
rect 6126 9220 6182 9276
rect 6182 9220 6186 9276
rect 6122 9216 6186 9220
rect 10813 9276 10877 9280
rect 10813 9220 10817 9276
rect 10817 9220 10873 9276
rect 10873 9220 10877 9276
rect 10813 9216 10877 9220
rect 10893 9276 10957 9280
rect 10893 9220 10897 9276
rect 10897 9220 10953 9276
rect 10953 9220 10957 9276
rect 10893 9216 10957 9220
rect 10973 9276 11037 9280
rect 10973 9220 10977 9276
rect 10977 9220 11033 9276
rect 11033 9220 11037 9276
rect 10973 9216 11037 9220
rect 11053 9276 11117 9280
rect 11053 9220 11057 9276
rect 11057 9220 11113 9276
rect 11113 9220 11117 9276
rect 11053 9216 11117 9220
rect 10180 9208 10244 9212
rect 11836 9284 11900 9348
rect 10180 9152 10194 9208
rect 10194 9152 10244 9208
rect 10180 9148 10244 9152
rect 12388 9148 12452 9212
rect 2452 9012 2516 9076
rect 9628 9012 9692 9076
rect 11284 9012 11348 9076
rect 11652 8740 11716 8804
rect 3417 8732 3481 8736
rect 3417 8676 3421 8732
rect 3421 8676 3477 8732
rect 3477 8676 3481 8732
rect 3417 8672 3481 8676
rect 3497 8732 3561 8736
rect 3497 8676 3501 8732
rect 3501 8676 3557 8732
rect 3557 8676 3561 8732
rect 3497 8672 3561 8676
rect 3577 8732 3641 8736
rect 3577 8676 3581 8732
rect 3581 8676 3637 8732
rect 3637 8676 3641 8732
rect 3577 8672 3641 8676
rect 3657 8732 3721 8736
rect 3657 8676 3661 8732
rect 3661 8676 3717 8732
rect 3717 8676 3721 8732
rect 3657 8672 3721 8676
rect 8348 8732 8412 8736
rect 8348 8676 8352 8732
rect 8352 8676 8408 8732
rect 8408 8676 8412 8732
rect 8348 8672 8412 8676
rect 8428 8732 8492 8736
rect 8428 8676 8432 8732
rect 8432 8676 8488 8732
rect 8488 8676 8492 8732
rect 8428 8672 8492 8676
rect 8508 8732 8572 8736
rect 8508 8676 8512 8732
rect 8512 8676 8568 8732
rect 8568 8676 8572 8732
rect 8508 8672 8572 8676
rect 8588 8732 8652 8736
rect 8588 8676 8592 8732
rect 8592 8676 8648 8732
rect 8648 8676 8652 8732
rect 8588 8672 8652 8676
rect 13124 8740 13188 8804
rect 13278 8732 13342 8736
rect 13278 8676 13282 8732
rect 13282 8676 13338 8732
rect 13338 8676 13342 8732
rect 13278 8672 13342 8676
rect 13358 8732 13422 8736
rect 13358 8676 13362 8732
rect 13362 8676 13418 8732
rect 13418 8676 13422 8732
rect 13358 8672 13422 8676
rect 13438 8732 13502 8736
rect 13438 8676 13442 8732
rect 13442 8676 13498 8732
rect 13498 8676 13502 8732
rect 13438 8672 13502 8676
rect 13518 8732 13582 8736
rect 13518 8676 13522 8732
rect 13522 8676 13578 8732
rect 13578 8676 13582 8732
rect 13518 8672 13582 8676
rect 12572 8604 12636 8668
rect 14412 8604 14476 8668
rect 6684 8468 6748 8532
rect 8892 8468 8956 8532
rect 9812 8468 9876 8532
rect 12020 8468 12084 8532
rect 12572 8468 12636 8532
rect 9076 8256 9140 8260
rect 9076 8200 9126 8256
rect 9126 8200 9140 8256
rect 9076 8196 9140 8200
rect 11284 8196 11348 8260
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 6122 8188 6186 8192
rect 6122 8132 6126 8188
rect 6126 8132 6182 8188
rect 6182 8132 6186 8188
rect 6122 8128 6186 8132
rect 10813 8188 10877 8192
rect 10813 8132 10817 8188
rect 10817 8132 10873 8188
rect 10873 8132 10877 8188
rect 10813 8128 10877 8132
rect 10893 8188 10957 8192
rect 10893 8132 10897 8188
rect 10897 8132 10953 8188
rect 10953 8132 10957 8188
rect 10893 8128 10957 8132
rect 10973 8188 11037 8192
rect 10973 8132 10977 8188
rect 10977 8132 11033 8188
rect 11033 8132 11037 8188
rect 10973 8128 11037 8132
rect 11053 8188 11117 8192
rect 11053 8132 11057 8188
rect 11057 8132 11113 8188
rect 11113 8132 11117 8188
rect 11053 8128 11117 8132
rect 11468 8120 11532 8124
rect 11468 8064 11518 8120
rect 11518 8064 11532 8120
rect 11468 8060 11532 8064
rect 13676 8060 13740 8124
rect 12756 7652 12820 7716
rect 3417 7644 3481 7648
rect 3417 7588 3421 7644
rect 3421 7588 3477 7644
rect 3477 7588 3481 7644
rect 3417 7584 3481 7588
rect 3497 7644 3561 7648
rect 3497 7588 3501 7644
rect 3501 7588 3557 7644
rect 3557 7588 3561 7644
rect 3497 7584 3561 7588
rect 3577 7644 3641 7648
rect 3577 7588 3581 7644
rect 3581 7588 3637 7644
rect 3637 7588 3641 7644
rect 3577 7584 3641 7588
rect 3657 7644 3721 7648
rect 3657 7588 3661 7644
rect 3661 7588 3717 7644
rect 3717 7588 3721 7644
rect 3657 7584 3721 7588
rect 8348 7644 8412 7648
rect 8348 7588 8352 7644
rect 8352 7588 8408 7644
rect 8408 7588 8412 7644
rect 8348 7584 8412 7588
rect 8428 7644 8492 7648
rect 8428 7588 8432 7644
rect 8432 7588 8488 7644
rect 8488 7588 8492 7644
rect 8428 7584 8492 7588
rect 8508 7644 8572 7648
rect 8508 7588 8512 7644
rect 8512 7588 8568 7644
rect 8568 7588 8572 7644
rect 8508 7584 8572 7588
rect 8588 7644 8652 7648
rect 8588 7588 8592 7644
rect 8592 7588 8648 7644
rect 8648 7588 8652 7644
rect 8588 7584 8652 7588
rect 13278 7644 13342 7648
rect 13278 7588 13282 7644
rect 13282 7588 13338 7644
rect 13338 7588 13342 7644
rect 13278 7584 13342 7588
rect 13358 7644 13422 7648
rect 13358 7588 13362 7644
rect 13362 7588 13418 7644
rect 13418 7588 13422 7644
rect 13358 7584 13422 7588
rect 13438 7644 13502 7648
rect 13438 7588 13442 7644
rect 13442 7588 13498 7644
rect 13498 7588 13502 7644
rect 13438 7584 13502 7588
rect 13518 7644 13582 7648
rect 13518 7588 13522 7644
rect 13522 7588 13578 7644
rect 13578 7588 13582 7644
rect 13518 7584 13582 7588
rect 11284 7516 11348 7580
rect 12020 7516 12084 7580
rect 12204 7516 12268 7580
rect 12572 7516 12636 7580
rect 13124 7108 13188 7172
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 6122 7100 6186 7104
rect 6122 7044 6126 7100
rect 6126 7044 6182 7100
rect 6182 7044 6186 7100
rect 6122 7040 6186 7044
rect 10813 7100 10877 7104
rect 10813 7044 10817 7100
rect 10817 7044 10873 7100
rect 10873 7044 10877 7100
rect 10813 7040 10877 7044
rect 10893 7100 10957 7104
rect 10893 7044 10897 7100
rect 10897 7044 10953 7100
rect 10953 7044 10957 7100
rect 10893 7040 10957 7044
rect 10973 7100 11037 7104
rect 10973 7044 10977 7100
rect 10977 7044 11033 7100
rect 11033 7044 11037 7100
rect 10973 7040 11037 7044
rect 11053 7100 11117 7104
rect 11053 7044 11057 7100
rect 11057 7044 11113 7100
rect 11113 7044 11117 7100
rect 11053 7040 11117 7044
rect 11468 6836 11532 6900
rect 9260 6564 9324 6628
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 2452 6156 2516 6220
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 12388 6216 12452 6220
rect 12388 6160 12438 6216
rect 12438 6160 12452 6216
rect 12388 6156 12452 6160
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 13676 5884 13740 5948
rect 14044 5612 14108 5676
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 9628 5476 9692 5540
rect 12572 5476 12636 5540
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 8892 5340 8956 5404
rect 9444 4992 9508 4996
rect 9444 4936 9458 4992
rect 9458 4936 9508 4992
rect 9444 4932 9508 4936
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 12940 4660 13004 4724
rect 10548 4388 10612 4452
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 11284 4312 11348 4316
rect 11284 4256 11334 4312
rect 11334 4256 11348 4312
rect 11284 4252 11348 4256
rect 11836 4116 11900 4180
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 9444 3708 9508 3772
rect 14412 3904 14476 3908
rect 14412 3848 14462 3904
rect 14462 3848 14476 3904
rect 14412 3844 14476 3848
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 12388 3708 12452 3772
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 10364 3224 10428 3228
rect 10364 3168 10414 3224
rect 10414 3168 10428 3224
rect 10364 3164 10428 3168
rect 11652 3164 11716 3228
rect 12756 3164 12820 3228
rect 9076 2756 9140 2820
rect 9260 2816 9324 2820
rect 9260 2760 9274 2816
rect 9274 2760 9324 2816
rect 9260 2756 9324 2760
rect 9996 2816 10060 2820
rect 9996 2760 10010 2816
rect 10010 2760 10060 2816
rect 9996 2756 10060 2760
rect 13124 2756 13188 2820
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 10180 2620 10244 2684
rect 9812 2348 9876 2412
rect 14044 2348 14108 2412
rect 9444 2212 9508 2276
rect 12204 2212 12268 2276
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
<< metal4 >>
rect 3409 17440 3729 17456
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3187 16964 3253 16965
rect 3187 16900 3188 16964
rect 3252 16900 3253 16964
rect 3187 16899 3253 16900
rect 3190 10437 3250 16899
rect 3409 16352 3729 17376
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 15264 3729 16288
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 14176 3729 15200
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 13088 3729 14112
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 12000 3729 13024
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 10912 3729 11936
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3187 10436 3253 10437
rect 3187 10372 3188 10436
rect 3252 10372 3253 10436
rect 3187 10371 3253 10372
rect 3409 9824 3729 10848
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 2451 9076 2517 9077
rect 2451 9012 2452 9076
rect 2516 9012 2517 9076
rect 2451 9011 2517 9012
rect 2454 6221 2514 9011
rect 3409 8736 3729 9760
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 7648 3729 8672
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 6560 3729 7584
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 2451 6220 2517 6221
rect 2451 6156 2452 6220
rect 2516 6156 2517 6220
rect 2451 6155 2517 6156
rect 3409 5472 3729 6496
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 3296 3729 4320
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 2208 3729 3232
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 5874 16896 6195 17456
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6195 16896
rect 5874 15808 6195 16832
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6195 15808
rect 5874 14720 6195 15744
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6195 14720
rect 5874 13632 6195 14656
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6195 13632
rect 5874 12544 6195 13568
rect 8340 17440 8660 17456
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 16352 8660 17376
rect 9627 17236 9693 17237
rect 9627 17172 9628 17236
rect 9692 17172 9693 17236
rect 9627 17171 9693 17172
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 15264 8660 16288
rect 9443 15740 9509 15741
rect 9443 15676 9444 15740
rect 9508 15676 9509 15740
rect 9443 15675 9509 15676
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 14176 8660 15200
rect 9259 15196 9325 15197
rect 9259 15132 9260 15196
rect 9324 15132 9325 15196
rect 9259 15131 9325 15132
rect 8891 14652 8957 14653
rect 8891 14588 8892 14652
rect 8956 14588 8957 14652
rect 8891 14587 8957 14588
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 13088 8660 14112
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 6683 12884 6749 12885
rect 6683 12820 6684 12884
rect 6748 12820 6749 12884
rect 6683 12819 6749 12820
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6195 12544
rect 5874 11456 6195 12480
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6195 11456
rect 5874 10368 6195 11392
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6195 10368
rect 5874 9280 6195 10304
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6195 9280
rect 5874 8192 6195 9216
rect 6686 8533 6746 12819
rect 8340 12000 8660 13024
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 10912 8660 11936
rect 8894 11525 8954 14587
rect 9075 14516 9141 14517
rect 9075 14452 9076 14516
rect 9140 14452 9141 14516
rect 9075 14451 9141 14452
rect 9078 14109 9138 14451
rect 9075 14108 9141 14109
rect 9075 14044 9076 14108
rect 9140 14044 9141 14108
rect 9075 14043 9141 14044
rect 9262 13565 9322 15131
rect 9446 13701 9506 15675
rect 9630 14653 9690 17171
rect 10179 17100 10245 17101
rect 10179 17036 10180 17100
rect 10244 17036 10245 17100
rect 10179 17035 10245 17036
rect 9811 16828 9877 16829
rect 9811 16764 9812 16828
rect 9876 16764 9877 16828
rect 9811 16763 9877 16764
rect 9627 14652 9693 14653
rect 9627 14588 9628 14652
rect 9692 14588 9693 14652
rect 9627 14587 9693 14588
rect 9627 14516 9693 14517
rect 9627 14452 9628 14516
rect 9692 14452 9693 14516
rect 9627 14451 9693 14452
rect 9443 13700 9509 13701
rect 9443 13636 9444 13700
rect 9508 13636 9509 13700
rect 9443 13635 9509 13636
rect 9259 13564 9325 13565
rect 9259 13500 9260 13564
rect 9324 13500 9325 13564
rect 9259 13499 9325 13500
rect 9443 13564 9509 13565
rect 9443 13500 9444 13564
rect 9508 13500 9509 13564
rect 9443 13499 9509 13500
rect 9075 13292 9141 13293
rect 9075 13228 9076 13292
rect 9140 13228 9141 13292
rect 9075 13227 9141 13228
rect 8891 11524 8957 11525
rect 8891 11460 8892 11524
rect 8956 11460 8957 11524
rect 8891 11459 8957 11460
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 9824 8660 10848
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 8736 8660 9760
rect 9078 9757 9138 13227
rect 9446 11253 9506 13499
rect 9630 11525 9690 14451
rect 9814 12341 9874 16763
rect 9995 16420 10061 16421
rect 9995 16356 9996 16420
rect 10060 16356 10061 16420
rect 9995 16355 10061 16356
rect 9998 13565 10058 16355
rect 9995 13564 10061 13565
rect 9995 13500 9996 13564
rect 10060 13500 10061 13564
rect 9995 13499 10061 13500
rect 9811 12340 9877 12341
rect 9811 12276 9812 12340
rect 9876 12276 9877 12340
rect 9811 12275 9877 12276
rect 9811 12204 9877 12205
rect 9811 12140 9812 12204
rect 9876 12140 9877 12204
rect 9811 12139 9877 12140
rect 9627 11524 9693 11525
rect 9627 11460 9628 11524
rect 9692 11460 9693 11524
rect 9627 11459 9693 11460
rect 9443 11252 9509 11253
rect 9443 11188 9444 11252
rect 9508 11188 9509 11252
rect 9443 11187 9509 11188
rect 9443 10708 9509 10709
rect 9443 10644 9444 10708
rect 9508 10644 9509 10708
rect 9814 10706 9874 12139
rect 9998 10845 10058 13499
rect 10182 12885 10242 17035
rect 10805 16896 11125 17456
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10363 16692 10429 16693
rect 10363 16628 10364 16692
rect 10428 16628 10429 16692
rect 10363 16627 10429 16628
rect 10179 12884 10245 12885
rect 10179 12820 10180 12884
rect 10244 12820 10245 12884
rect 10179 12819 10245 12820
rect 10182 12069 10242 12819
rect 10179 12068 10245 12069
rect 10179 12004 10180 12068
rect 10244 12004 10245 12068
rect 10179 12003 10245 12004
rect 9995 10844 10061 10845
rect 9995 10780 9996 10844
rect 10060 10780 10061 10844
rect 9995 10779 10061 10780
rect 9814 10646 10058 10706
rect 9443 10643 9509 10644
rect 9075 9756 9141 9757
rect 9075 9692 9076 9756
rect 9140 9692 9141 9756
rect 9075 9691 9141 9692
rect 9446 9349 9506 10643
rect 9998 9757 10058 10646
rect 9995 9756 10061 9757
rect 9995 9692 9996 9756
rect 10060 9692 10061 9756
rect 9995 9691 10061 9692
rect 9443 9348 9509 9349
rect 9443 9284 9444 9348
rect 9508 9284 9509 9348
rect 9443 9283 9509 9284
rect 9627 9076 9693 9077
rect 9627 9012 9628 9076
rect 9692 9012 9693 9076
rect 9627 9011 9693 9012
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 6683 8532 6749 8533
rect 6683 8468 6684 8532
rect 6748 8468 6749 8532
rect 6683 8467 6749 8468
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6195 8192
rect 5874 7104 6195 8128
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6195 7104
rect 5874 6016 6195 7040
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5874 3840 6195 4864
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5874 2752 6195 3776
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 5874 2128 6195 2688
rect 8340 7648 8660 8672
rect 8891 8532 8957 8533
rect 8891 8468 8892 8532
rect 8956 8468 8957 8532
rect 8891 8467 8957 8468
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 6560 8660 7584
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 5472 8660 6496
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8894 5405 8954 8467
rect 9075 8260 9141 8261
rect 9075 8196 9076 8260
rect 9140 8196 9141 8260
rect 9075 8195 9141 8196
rect 8891 5404 8957 5405
rect 8891 5340 8892 5404
rect 8956 5340 8957 5404
rect 8891 5339 8957 5340
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 3296 8660 4320
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 2208 8660 3232
rect 9078 2821 9138 8195
rect 9259 6628 9325 6629
rect 9259 6564 9260 6628
rect 9324 6564 9325 6628
rect 9259 6563 9325 6564
rect 9262 2821 9322 6563
rect 9630 5541 9690 9011
rect 9811 8532 9877 8533
rect 9811 8468 9812 8532
rect 9876 8468 9877 8532
rect 9811 8467 9877 8468
rect 9627 5540 9693 5541
rect 9627 5476 9628 5540
rect 9692 5476 9693 5540
rect 9627 5475 9693 5476
rect 9443 4996 9509 4997
rect 9443 4932 9444 4996
rect 9508 4932 9509 4996
rect 9443 4931 9509 4932
rect 9446 3773 9506 4931
rect 9443 3772 9509 3773
rect 9443 3708 9444 3772
rect 9508 3708 9509 3772
rect 9443 3707 9509 3708
rect 9075 2820 9141 2821
rect 9075 2756 9076 2820
rect 9140 2756 9141 2820
rect 9075 2755 9141 2756
rect 9259 2820 9325 2821
rect 9259 2756 9260 2820
rect 9324 2756 9325 2820
rect 9259 2755 9325 2756
rect 9446 2277 9506 3707
rect 9814 2413 9874 8467
rect 9998 2821 10058 9691
rect 10179 9212 10245 9213
rect 10179 9148 10180 9212
rect 10244 9148 10245 9212
rect 10179 9147 10245 9148
rect 9995 2820 10061 2821
rect 9995 2756 9996 2820
rect 10060 2756 10061 2820
rect 9995 2755 10061 2756
rect 10182 2685 10242 9147
rect 10366 3229 10426 16627
rect 10805 15808 11125 16832
rect 13270 17440 13590 17456
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 12571 16556 12637 16557
rect 12571 16492 12572 16556
rect 12636 16492 12637 16556
rect 12571 16491 12637 16492
rect 12574 16285 12634 16491
rect 13270 16352 13590 17376
rect 13675 16692 13741 16693
rect 13675 16628 13676 16692
rect 13740 16628 13741 16692
rect 13675 16627 13741 16628
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 12571 16284 12637 16285
rect 12571 16220 12572 16284
rect 12636 16220 12637 16284
rect 12571 16219 12637 16220
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10547 15332 10613 15333
rect 10547 15268 10548 15332
rect 10612 15268 10613 15332
rect 10547 15267 10613 15268
rect 10550 11797 10610 15267
rect 10805 14720 11125 15744
rect 12203 15740 12269 15741
rect 12203 15676 12204 15740
rect 12268 15676 12269 15740
rect 12203 15675 12269 15676
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 13632 11125 14656
rect 11283 14516 11349 14517
rect 11283 14452 11284 14516
rect 11348 14452 11349 14516
rect 11283 14451 11349 14452
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 12544 11125 13568
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10547 11796 10613 11797
rect 10547 11732 10548 11796
rect 10612 11732 10613 11796
rect 10547 11731 10613 11732
rect 10550 4453 10610 11731
rect 10805 11456 11125 12480
rect 11286 11933 11346 14451
rect 11467 14244 11533 14245
rect 11467 14180 11468 14244
rect 11532 14180 11533 14244
rect 11467 14179 11533 14180
rect 11470 12477 11530 14179
rect 12019 14108 12085 14109
rect 12019 14044 12020 14108
rect 12084 14044 12085 14108
rect 12019 14043 12085 14044
rect 11651 13564 11717 13565
rect 11651 13500 11652 13564
rect 11716 13500 11717 13564
rect 11651 13499 11717 13500
rect 11467 12476 11533 12477
rect 11467 12412 11468 12476
rect 11532 12412 11533 12476
rect 11467 12411 11533 12412
rect 11283 11932 11349 11933
rect 11283 11868 11284 11932
rect 11348 11868 11349 11932
rect 11283 11867 11349 11868
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 10368 11125 11392
rect 11470 11386 11530 12411
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 9280 11125 10304
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 8192 11125 9216
rect 11286 11326 11530 11386
rect 11286 9077 11346 11326
rect 11467 11252 11533 11253
rect 11467 11188 11468 11252
rect 11532 11188 11533 11252
rect 11467 11187 11533 11188
rect 11470 10981 11530 11187
rect 11467 10980 11533 10981
rect 11467 10916 11468 10980
rect 11532 10916 11533 10980
rect 11467 10915 11533 10916
rect 11467 10844 11533 10845
rect 11467 10780 11468 10844
rect 11532 10780 11533 10844
rect 11467 10779 11533 10780
rect 11283 9076 11349 9077
rect 11283 9012 11284 9076
rect 11348 9012 11349 9076
rect 11283 9011 11349 9012
rect 11470 8530 11530 10779
rect 11654 9893 11714 13499
rect 12022 12885 12082 14043
rect 11835 12884 11901 12885
rect 11835 12820 11836 12884
rect 11900 12820 11901 12884
rect 11835 12819 11901 12820
rect 12019 12884 12085 12885
rect 12019 12820 12020 12884
rect 12084 12820 12085 12884
rect 12019 12819 12085 12820
rect 11838 10845 11898 12819
rect 12019 12612 12085 12613
rect 12019 12548 12020 12612
rect 12084 12548 12085 12612
rect 12019 12547 12085 12548
rect 12022 11253 12082 12547
rect 12019 11252 12085 11253
rect 12019 11188 12020 11252
rect 12084 11188 12085 11252
rect 12019 11187 12085 11188
rect 12019 10980 12085 10981
rect 12019 10916 12020 10980
rect 12084 10916 12085 10980
rect 12019 10915 12085 10916
rect 11835 10844 11901 10845
rect 11835 10780 11836 10844
rect 11900 10780 11901 10844
rect 11835 10779 11901 10780
rect 11835 10436 11901 10437
rect 11835 10372 11836 10436
rect 11900 10372 11901 10436
rect 11835 10371 11901 10372
rect 11651 9892 11717 9893
rect 11651 9828 11652 9892
rect 11716 9828 11717 9892
rect 11651 9827 11717 9828
rect 11838 9349 11898 10371
rect 11835 9348 11901 9349
rect 11835 9284 11836 9348
rect 11900 9284 11901 9348
rect 11835 9283 11901 9284
rect 11651 8804 11717 8805
rect 11651 8740 11652 8804
rect 11716 8740 11717 8804
rect 11651 8739 11717 8740
rect 11286 8470 11530 8530
rect 11286 8261 11346 8470
rect 11283 8260 11349 8261
rect 11283 8196 11284 8260
rect 11348 8196 11349 8260
rect 11283 8195 11349 8196
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 7104 11125 8128
rect 11286 7581 11346 8195
rect 11467 8124 11533 8125
rect 11467 8060 11468 8124
rect 11532 8060 11533 8124
rect 11467 8059 11533 8060
rect 11283 7580 11349 7581
rect 11283 7516 11284 7580
rect 11348 7516 11349 7580
rect 11283 7515 11349 7516
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 6016 11125 7040
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10547 4452 10613 4453
rect 10547 4388 10548 4452
rect 10612 4388 10613 4452
rect 10547 4387 10613 4388
rect 10805 3840 11125 4864
rect 11286 4317 11346 7515
rect 11470 6901 11530 8059
rect 11467 6900 11533 6901
rect 11467 6836 11468 6900
rect 11532 6836 11533 6900
rect 11467 6835 11533 6836
rect 11283 4316 11349 4317
rect 11283 4252 11284 4316
rect 11348 4252 11349 4316
rect 11283 4251 11349 4252
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10363 3228 10429 3229
rect 10363 3164 10364 3228
rect 10428 3164 10429 3228
rect 10363 3163 10429 3164
rect 10805 2752 11125 3776
rect 11654 3229 11714 8739
rect 11838 4181 11898 9283
rect 12022 8533 12082 10915
rect 12206 9893 12266 15675
rect 12387 15604 12453 15605
rect 12387 15540 12388 15604
rect 12452 15540 12453 15604
rect 12387 15539 12453 15540
rect 12390 11525 12450 15539
rect 12387 11524 12453 11525
rect 12387 11460 12388 11524
rect 12452 11460 12453 11524
rect 12387 11459 12453 11460
rect 12387 11252 12453 11253
rect 12387 11188 12388 11252
rect 12452 11188 12453 11252
rect 12387 11187 12453 11188
rect 12390 10437 12450 11187
rect 12387 10436 12453 10437
rect 12387 10372 12388 10436
rect 12452 10372 12453 10436
rect 12387 10371 12453 10372
rect 12203 9892 12269 9893
rect 12203 9828 12204 9892
rect 12268 9828 12269 9892
rect 12203 9827 12269 9828
rect 12203 9484 12269 9485
rect 12203 9420 12204 9484
rect 12268 9420 12269 9484
rect 12203 9419 12269 9420
rect 12019 8532 12085 8533
rect 12019 8468 12020 8532
rect 12084 8468 12085 8532
rect 12019 8467 12085 8468
rect 12206 7850 12266 9419
rect 12387 9212 12453 9213
rect 12387 9148 12388 9212
rect 12452 9148 12453 9212
rect 12387 9147 12453 9148
rect 12022 7790 12266 7850
rect 12022 7581 12082 7790
rect 12019 7580 12085 7581
rect 12019 7516 12020 7580
rect 12084 7516 12085 7580
rect 12019 7515 12085 7516
rect 12203 7580 12269 7581
rect 12203 7516 12204 7580
rect 12268 7516 12269 7580
rect 12203 7515 12269 7516
rect 11835 4180 11901 4181
rect 11835 4116 11836 4180
rect 11900 4116 11901 4180
rect 11835 4115 11901 4116
rect 11651 3228 11717 3229
rect 11651 3164 11652 3228
rect 11716 3164 11717 3228
rect 11651 3163 11717 3164
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10179 2684 10245 2685
rect 10179 2620 10180 2684
rect 10244 2620 10245 2684
rect 10179 2619 10245 2620
rect 9811 2412 9877 2413
rect 9811 2348 9812 2412
rect 9876 2348 9877 2412
rect 9811 2347 9877 2348
rect 9443 2276 9509 2277
rect 9443 2212 9444 2276
rect 9508 2212 9509 2276
rect 9443 2211 9509 2212
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 10805 2128 11125 2688
rect 12206 2277 12266 7515
rect 12390 7170 12450 9147
rect 12574 8669 12634 16219
rect 13270 15264 13590 16288
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 12755 15060 12821 15061
rect 12755 14996 12756 15060
rect 12820 14996 12821 15060
rect 12755 14995 12821 14996
rect 12758 10165 12818 14995
rect 12939 14652 13005 14653
rect 12939 14588 12940 14652
rect 13004 14588 13005 14652
rect 12939 14587 13005 14588
rect 12942 10437 13002 14587
rect 13270 14176 13590 15200
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 13088 13590 14112
rect 13678 13157 13738 16627
rect 13675 13156 13741 13157
rect 13675 13092 13676 13156
rect 13740 13092 13741 13156
rect 13675 13091 13741 13092
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 12000 13590 13024
rect 13675 12340 13741 12341
rect 13675 12276 13676 12340
rect 13740 12276 13741 12340
rect 13675 12275 13741 12276
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13123 11796 13189 11797
rect 13123 11732 13124 11796
rect 13188 11732 13189 11796
rect 13123 11731 13189 11732
rect 12939 10436 13005 10437
rect 12939 10372 12940 10436
rect 13004 10372 13005 10436
rect 12939 10371 13005 10372
rect 12755 10164 12821 10165
rect 12755 10100 12756 10164
rect 12820 10100 12821 10164
rect 12755 10099 12821 10100
rect 12571 8668 12637 8669
rect 12571 8604 12572 8668
rect 12636 8604 12637 8668
rect 12571 8603 12637 8604
rect 12571 8532 12637 8533
rect 12571 8468 12572 8532
rect 12636 8468 12637 8532
rect 12571 8467 12637 8468
rect 12574 7581 12634 8467
rect 12758 7717 12818 10099
rect 13126 8805 13186 11731
rect 13270 10912 13590 11936
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 9824 13590 10848
rect 13678 10165 13738 12275
rect 13675 10164 13741 10165
rect 13675 10100 13676 10164
rect 13740 10100 13741 10164
rect 13675 10099 13741 10100
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13123 8804 13189 8805
rect 13123 8802 13124 8804
rect 12942 8742 13124 8802
rect 12755 7716 12821 7717
rect 12755 7652 12756 7716
rect 12820 7652 12821 7716
rect 12755 7651 12821 7652
rect 12571 7580 12637 7581
rect 12571 7516 12572 7580
rect 12636 7516 12637 7580
rect 12571 7515 12637 7516
rect 12390 7110 12634 7170
rect 12387 6220 12453 6221
rect 12387 6156 12388 6220
rect 12452 6156 12453 6220
rect 12387 6155 12453 6156
rect 12390 3773 12450 6155
rect 12574 5541 12634 7110
rect 12571 5540 12637 5541
rect 12571 5476 12572 5540
rect 12636 5476 12637 5540
rect 12571 5475 12637 5476
rect 12387 3772 12453 3773
rect 12387 3708 12388 3772
rect 12452 3708 12453 3772
rect 12387 3707 12453 3708
rect 12758 3229 12818 7651
rect 12942 4725 13002 8742
rect 13123 8740 13124 8742
rect 13188 8740 13189 8804
rect 13123 8739 13189 8740
rect 13270 8736 13590 9760
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 7648 13590 8672
rect 14411 8668 14477 8669
rect 14411 8604 14412 8668
rect 14476 8604 14477 8668
rect 14411 8603 14477 8604
rect 13675 8124 13741 8125
rect 13675 8060 13676 8124
rect 13740 8060 13741 8124
rect 13675 8059 13741 8060
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13123 7172 13189 7173
rect 13123 7108 13124 7172
rect 13188 7108 13189 7172
rect 13123 7107 13189 7108
rect 12939 4724 13005 4725
rect 12939 4660 12940 4724
rect 13004 4660 13005 4724
rect 12939 4659 13005 4660
rect 12755 3228 12821 3229
rect 12755 3164 12756 3228
rect 12820 3164 12821 3228
rect 12755 3163 12821 3164
rect 13126 2821 13186 7107
rect 13270 6560 13590 7584
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 5472 13590 6496
rect 13678 5949 13738 8059
rect 13675 5948 13741 5949
rect 13675 5884 13676 5948
rect 13740 5884 13741 5948
rect 13675 5883 13741 5884
rect 14043 5676 14109 5677
rect 14043 5612 14044 5676
rect 14108 5612 14109 5676
rect 14043 5611 14109 5612
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 3296 13590 4320
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13123 2820 13189 2821
rect 13123 2756 13124 2820
rect 13188 2756 13189 2820
rect 13123 2755 13189 2756
rect 12203 2276 12269 2277
rect 12203 2212 12204 2276
rect 12268 2212 12269 2276
rect 12203 2211 12269 2212
rect 13270 2208 13590 3232
rect 14046 2413 14106 5611
rect 14414 3909 14474 8603
rect 14411 3908 14477 3909
rect 14411 3844 14412 3908
rect 14476 3844 14477 3908
rect 14411 3843 14477 3844
rect 14043 2412 14109 2413
rect 14043 2348 14044 2412
rect 14108 2348 14109 2412
rect 14043 2347 14109 2348
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2128 13590 2144
use sky130_fd_sc_hd__buf_2  _53_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2116 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2484 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_S_FTB01 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1564 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1606256979
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4876 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1606256979
transform 1 0 3680 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1606256979
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1606256979
transform 1 0 4600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 1606256979
transform 1 0 3312 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1606256979
transform 1 0 4508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4968 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58
timestamp 1606256979
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1606256979
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1606256979
transform 1 0 8648 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1606256979
transform 1 0 7728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1606256979
transform 1 0 8280 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1606256979
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1606256979
transform 1 0 8924 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_right_ipin_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9292 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1606256979
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1606256979
transform 1 0 9844 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_104
timestamp 1606256979
transform 1 0 10672 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11040 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1606256979
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1606256979
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1606256979
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116
timestamp 1606256979
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 12144 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13616 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_134
timestamp 1606256979
transform 1 0 13432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1606256979
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1606256979
transform 1 0 14444 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606256979
transform 1 0 14812 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 14996 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_147
timestamp 1606256979
transform 1 0 14628 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1606256979
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_153
timestamp 1606256979
transform 1 0 15180 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1564 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2760 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1606256979
transform 1 0 2392 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4508 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606256979
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_36
timestamp 1606256979
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5704 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_46
timestamp 1606256979
transform 1 0 5336 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7544 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1606256979
transform 1 0 7176 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9016 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1606256979
transform 1 0 10488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10856 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12052 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1606256979
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1606256979
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 13248 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1606256979
transform 1 0 12880 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1606256979
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1606256979
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1606256979
transform 1 0 1840 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1606256979
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_17
timestamp 1606256979
transform 1 0 2668 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 3036 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4876 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1606256979
transform 1 0 4508 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1606256979
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8648 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1606256979
transform 1 0 8280 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1606256979
transform 1 0 9844 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_91
timestamp 1606256979
transform 1 0 9476 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_104
timestamp 1606256979
transform 1 0 10672 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11040 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1606256979
transform 1 0 11868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1606256979
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13616 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1606256979
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1606256979
transform 1 0 14444 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606256979
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_153
timestamp 1606256979
transform 1 0 15180 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2116 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1606256979
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606256979
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1606256979
transform 1 0 4876 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5244 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_61
timestamp 1606256979
transform 1 0 6716 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7084 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_81
timestamp 1606256979
transform 1 0 8556 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _16_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 8924 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1606256979
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1606256979
transform 1 0 10488 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10856 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_115
timestamp 1606256979
transform 1 0 11684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1606256979
transform 1 0 14444 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13248 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp 1606256979
transform 1 0 12880 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1606256979
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1606256979
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1840 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1606256979
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_17
timestamp 1606256979
transform 1 0 2668 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4876 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 3036 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1606256979
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1606256979
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8648 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1606256979
transform 1 0 8280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10488 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_98
timestamp 1606256979
transform 1 0 10120 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1606256979
transform 1 0 11684 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_111
timestamp 1606256979
transform 1 0 11316 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1606256979
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13616 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1606256979
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_132
timestamp 1606256979
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1606256979
transform 1 0 14444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1606256979
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_153
timestamp 1606256979
transform 1 0 15180 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2116 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1606256979
transform 1 0 1840 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1606256979
transform 1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1606256979
transform 1 0 1748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1606256979
transform 1 0 2668 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 3036 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4876 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1606256979
transform 1 0 4232 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606256979
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1606256979
transform 1 0 4508 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5428 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_43
timestamp 1606256979
transform 1 0 5060 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1606256979
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7268 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 8648 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_63
timestamp 1606256979
transform 1 0 6900 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_83
timestamp 1606256979
transform 1 0 8740 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1606256979
transform 1 0 8280 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1606256979
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1606256979
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1606256979
transform 1 0 10120 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1606256979
transform 1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1606256979
transform 1 0 11500 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1606256979
transform 1 0 11132 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_122
timestamp 1606256979
transform 1 0 12328 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_111
timestamp 1606256979
transform 1 0 11316 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1606256979
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13616 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13892 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1606256979
transform 1 0 12696 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1606256979
transform 1 0 13524 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1606256979
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1606256979
transform 1 0 14444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1606256979
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_148
timestamp 1606256979
transform 1 0 14720 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1606256979
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1606256979
transform 1 0 15180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2116 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1606256979
transform 1 0 1748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4232 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606256979
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 5704 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_46
timestamp 1606256979
transform 1 0 5336 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7544 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_66
timestamp 1606256979
transform 1 0 7176 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_86
timestamp 1606256979
transform 1 0 9016 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_102
timestamp 1606256979
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1606256979
transform 1 0 10856 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1606256979
transform 1 0 12052 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_115
timestamp 1606256979
transform 1 0 11684 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1606256979
transform 1 0 14444 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13248 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1606256979
transform 1 0 12880 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1606256979
transform 1 0 14076 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1606256979
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1840 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1606256979
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_17
timestamp 1606256979
transform 1 0 2668 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 3036 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4876 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_37
timestamp 1606256979
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1606256979
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8648 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_78
timestamp 1606256979
transform 1 0 8280 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1606256979
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1606256979
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1606256979
transform 1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_111
timestamp 1606256979
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1606256979
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1606256979
transform 1 0 13616 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1606256979
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_145
timestamp 1606256979
transform 1 0 14444 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1606256979
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1606256979
transform 1 0 15180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2760 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 1564 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1606256979
transform 1 0 2392 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606256979
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5888 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1606256979
transform 1 0 5520 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7728 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 1606256979
transform 1 0 7360 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1606256979
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_102
timestamp 1606256979
transform 1 0 10488 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1606256979
transform 1 0 10856 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12052 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_115
timestamp 1606256979
transform 1 0 11684 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1606256979
transform 1 0 14444 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13248 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_128
timestamp 1606256979
transform 1 0 12880 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1606256979
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1606256979
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2484 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1606256979
transform 1 0 2116 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4876 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1606256979
transform 1 0 3680 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1606256979
transform 1 0 3312 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_37
timestamp 1606256979
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1606256979
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8648 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_78
timestamp 1606256979
transform 1 0 8280 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1606256979
transform 1 0 9844 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1606256979
transform 1 0 9476 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_104
timestamp 1606256979
transform 1 0 10672 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11040 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1606256979
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1606256979
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1606256979
transform 1 0 13616 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp 1606256979
transform 1 0 13248 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_145
timestamp 1606256979
transform 1 0 14444 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1606256979
transform 1 0 14812 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1606256979
transform 1 0 15180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 1564 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 2760 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_14
timestamp 1606256979
transform 1 0 2392 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4232 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1606256979
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_right_ipin_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5888 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_12_43 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5060 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_51
timestamp 1606256979
transform 1 0 5796 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1606256979
transform 1 0 7728 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8556 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1606256979
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1606256979
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1606256979
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1606256979
transform 1 0 12052 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1606256979
transform 1 0 10856 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_115
timestamp 1606256979
transform 1 0 11684 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1606256979
transform 1 0 14444 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13248 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_128
timestamp 1606256979
transform 1 0 12880 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1606256979
transform 1 0 14076 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1606256979
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1606256979
transform 1 0 2392 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2760 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2116 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2944 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 3772 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4232 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606256979
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5428 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5244 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_43
timestamp 1606256979
transform 1 0 5060 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7268 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8648 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1606256979
transform 1 0 8280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_63
timestamp 1606256979
transform 1 0 6900 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_83
timestamp 1606256979
transform 1 0 8740 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1606256979
transform 1 0 9844 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 1606256979
transform 1 0 9476 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_104
timestamp 1606256979
transform 1 0 10672 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606256979
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1606256979
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12052 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1606256979
transform 1 0 11040 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1606256979
transform 1 0 10856 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_117
timestamp 1606256979
transform 1 0 11868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1606256979
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_115
timestamp 1606256979
transform 1 0 11684 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1606256979
transform 1 0 14444 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13616 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1606256979
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1606256979
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1606256979
transform 1 0 14444 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_128
timestamp 1606256979
transform 1 0 12880 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1606256979
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1606256979
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1606256979
transform 1 0 15180 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1606256979
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2484 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_11
timestamp 1606256979
transform 1 0 2116 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4876 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1606256979
transform 1 0 3680 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1606256979
transform 1 0 3312 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_37
timestamp 1606256979
transform 1 0 4508 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1606256979
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 8464 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 8004 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_71
timestamp 1606256979
transform 1 0 7636 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1606256979
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1606256979
transform 1 0 10304 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1606256979
transform 1 0 9936 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1606256979
transform 1 0 11500 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_109
timestamp 1606256979
transform 1 0 11132 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_117
timestamp 1606256979
transform 1 0 11868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1606256979
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13616 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1606256979
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_145
timestamp 1606256979
transform 1 0 14444 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1606256979
transform 1 0 14812 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1606256979
transform 1 0 15180 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1606256979
transform 1 0 2760 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1564 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_14
timestamp 1606256979
transform 1 0 2392 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4600 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606256979
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_32
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5796 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_47
timestamp 1606256979
transform 1 0 5428 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7636 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1606256979
transform 1 0 7268 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1606256979
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1606256979
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_102
timestamp 1606256979
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1606256979
transform 1 0 10856 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12052 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_115
timestamp 1606256979
transform 1 0 11684 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1606256979
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1606256979
transform 1 0 13248 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_128
timestamp 1606256979
transform 1 0 12880 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1606256979
transform 1 0 14076 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1606256979
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2484 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_11
timestamp 1606256979
transform 1 0 2116 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4876 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1606256979
transform 1 0 3680 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_24
timestamp 1606256979
transform 1 0 3312 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_37
timestamp 1606256979
transform 1 0 4508 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1606256979
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_62
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7360 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9200 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1606256979
transform 1 0 10396 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_84
timestamp 1606256979
transform 1 0 8832 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_97
timestamp 1606256979
transform 1 0 10028 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1606256979
transform 1 0 11592 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_110
timestamp 1606256979
transform 1 0 11224 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1606256979
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  Test_en_E_FTB01
timestamp 1606256979
transform 1 0 13616 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1606256979
transform 1 0 13248 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp 1606256979
transform 1 0 14168 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1606256979
transform 1 0 14536 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_152
timestamp 1606256979
transform 1 0 15088 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_156
timestamp 1606256979
transform 1 0 15456 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1606256979
transform 1 0 1564 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2760 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1606256979
transform 1 0 2392 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4324 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606256979
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_32
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5520 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_44
timestamp 1606256979
transform 1 0 5152 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7360 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_64
timestamp 1606256979
transform 1 0 6992 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 9200 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_84
timestamp 1606256979
transform 1 0 8832 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1606256979
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 1606256979
transform 1 0 10488 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10856 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12052 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_115
timestamp 1606256979
transform 1 0 11684 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606256979
transform 1 0 14444 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_2_S_FTB01
timestamp 1606256979
transform 1 0 13524 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 13248 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_128
timestamp 1606256979
transform 1 0 12880 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1606256979
transform 1 0 14076 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1606256979
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1606256979
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1606256979
transform 1 0 1564 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1606256979
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_14
timestamp 1606256979
transform 1 0 2392 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_17
timestamp 1606256979
transform 1 0 2668 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2760 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3036 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4324 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4876 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_37
timestamp 1606256979
transform 1 0 4508 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1606256979
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6164 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1606256979
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_51
timestamp 1606256979
transform 1 0 5796 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8648 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1606256979
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_78
timestamp 1606256979
transform 1 0 8280 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_71
timestamp 1606256979
transform 1 0 7636 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1606256979
transform 1 0 10488 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 9200 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1606256979
transform 1 0 10120 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_84
timestamp 1606256979
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606256979
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1606256979
transform 1 0 11684 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1606256979
transform 1 0 11500 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_111
timestamp 1606256979
transform 1 0 11316 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1606256979
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_109
timestamp 1606256979
transform 1 0 11132 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_122
timestamp 1606256979
transform 1 0 12328 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_3_S_FTB01
timestamp 1606256979
transform 1 0 13892 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12696 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13892 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 13616 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1606256979
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1606256979
transform 1 0 14444 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1606256979
transform 1 0 13524 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1606256979
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1606256979
transform 1 0 14812 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1606256979
transform 1 0 15180 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2484 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_11
timestamp 1606256979
transform 1 0 2116 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4876 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1606256979
transform 1 0 3680 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_24
timestamp 1606256979
transform 1 0 3312 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_37
timestamp 1606256979
transform 1 0 4508 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1606256979
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8648 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_78
timestamp 1606256979
transform 1 0 8280 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10488 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1606256979
transform 1 0 10120 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1606256979
transform 1 0 11684 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_111
timestamp 1606256979
transform 1 0 11316 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1606256979
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606256979
transform 1 0 13800 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_132
timestamp 1606256979
transform 1 0 13248 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_142
timestamp 1606256979
transform 1 0 14168 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1606256979
transform 1 0 14536 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1606256979
transform 1 0 14812 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2760 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1840 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1606256979
transform 1 0 1748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_14
timestamp 1606256979
transform 1 0 2392 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4416 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606256979
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5612 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_45
timestamp 1606256979
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7452 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_65
timestamp 1606256979
transform 1 0 7084 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1606256979
transform 1 0 8924 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1606256979
transform 1 0 10488 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12052 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1606256979
transform 1 0 10856 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_115
timestamp 1606256979
transform 1 0 11684 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_125
timestamp 1606256979
transform 1 0 12604 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1606256979
transform 1 0 14076 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606256979
transform 1 0 13340 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_137
timestamp 1606256979
transform 1 0 13708 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_144
timestamp 1606256979
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1606256979
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1606256979
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1748 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2668 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1606256979
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_13
timestamp 1606256979
transform 1 0 2300 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4876 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1606256979
transform 1 0 3680 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_23
timestamp 1606256979
transform 1 0 3220 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_27
timestamp 1606256979
transform 1 0 3588 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_37
timestamp 1606256979
transform 1 0 4508 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1606256979
transform 1 0 6348 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8648 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_78
timestamp 1606256979
transform 1 0 8280 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9844 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1606256979
transform 1 0 9476 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_104
timestamp 1606256979
transform 1 0 10672 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1606256979
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1606256979
transform 1 0 11040 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1606256979
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1606256979
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1606256979
transform 1 0 13064 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1606256979
transform 1 0 13708 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1606256979
transform 1 0 14352 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_126
timestamp 1606256979
transform 1 0 12696 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_133
timestamp 1606256979
transform 1 0 13340 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 1606256979
transform 1 0 13984 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp 1606256979
transform 1 0 14628 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1606256979
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2300 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1380 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_9
timestamp 1606256979
transform 1 0 1932 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_19
timestamp 1606256979
transform 1 0 2852 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1606256979
transform 1 0 3220 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4600 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1606256979
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_32
timestamp 1606256979
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5796 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_47
timestamp 1606256979
transform 1 0 5428 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1606256979
transform 1 0 7636 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_67
timestamp 1606256979
transform 1 0 7268 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1606256979
transform 1 0 8464 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606256979
transform 1 0 8832 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1606256979
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1606256979
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1606256979
transform 1 0 10488 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606256979
transform 1 0 10856 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606256979
transform 1 0 11592 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606256979
transform 1 0 12328 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1606256979
transform 1 0 11224 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_118
timestamp 1606256979
transform 1 0 11960 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1606256979
transform 1 0 13064 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1606256979
transform 1 0 13708 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_126
timestamp 1606256979
transform 1 0 12696 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_133
timestamp 1606256979
transform 1 0 13340 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_140 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 13984 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1606256979
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1606256979
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  clk_2_N_FTB01
timestamp 1606256979
transform 1 0 1472 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1606256979
transform 1 0 2392 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1606256979
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_10
timestamp 1606256979
transform 1 0 2024 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_20
timestamp 1606256979
transform 1 0 2944 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4324 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 3312 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 1606256979
transform 1 0 3864 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_34
timestamp 1606256979
transform 1 0 4232 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1606256979
transform 1 0 5520 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_44
timestamp 1606256979
transform 1 0 5152 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1606256979
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8004 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_71
timestamp 1606256979
transform 1 0 7636 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606256979
transform 1 0 10396 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1606256979
transform 1 0 9200 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_84
timestamp 1606256979
transform 1 0 8832 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1606256979
transform 1 0 10028 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606256979
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1606256979
transform 1 0 11132 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_105
timestamp 1606256979
transform 1 0 10764 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1606256979
transform 1 0 11500 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1606256979
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606256979
transform 1 0 13156 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_127
timestamp 1606256979
transform 1 0 12788 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1606256979
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_147
timestamp 1606256979
transform 1 0 14628 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1606256979
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1606256979
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1606256979
transform 1 0 1472 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  Test_en_W_FTB01
timestamp 1606256979
transform 1 0 1380 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_10
timestamp 1606256979
transform 1 0 2024 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_9
timestamp 1606256979
transform 1 0 1932 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_20
timestamp 1606256979
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 2484 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1606256979
transform 1 0 2760 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1606256979
transform 1 0 2392 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1606256979
transform 1 0 3588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1606256979
transform 1 0 3312 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606256979
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1606256979
transform 1 0 3312 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 4048 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01
timestamp 1606256979
transform 1 0 4048 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1606256979
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_38
timestamp 1606256979
transform 1 0 4600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606256979
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1606256979
transform 1 0 4968 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5612 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1606256979
transform 1 0 6256 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4968 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_51
timestamp 1606256979
transform 1 0 5796 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_55
timestamp 1606256979
transform 1 0 6164 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1606256979
transform 1 0 5244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_58
timestamp 1606256979
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8648 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6900 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1606256979
transform 1 0 8096 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1606256979
transform 1 0 7452 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_65
timestamp 1606256979
transform 1 0 7084 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_78
timestamp 1606256979
transform 1 0 8280 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_72
timestamp 1606256979
transform 1 0 7728 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1606256979
transform 1 0 8924 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1606256979
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_92
timestamp 1606256979
transform 1 0 9568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_right_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 9292 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606256979
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp 1606256979
transform 1 0 10028 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606256979
transform 1 0 9752 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_98
timestamp 1606256979
transform 1 0 10120 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606256979
transform 1 0 10396 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606256979
transform 1 0 10488 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_106
timestamp 1606256979
transform 1 0 10856 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_113
timestamp 1606256979
transform 1 0 11500 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_105
timestamp 1606256979
transform 1 0 10764 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606256979
transform 1 0 11132 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606256979
transform 1 0 11224 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_114
timestamp 1606256979
transform 1 0 11592 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_121
timestamp 1606256979
transform 1 0 12236 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606256979
transform 1 0 11868 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_122
timestamp 1606256979
transform 1 0 12328 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606256979
transform 1 0 12604 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606256979
transform 1 0 12604 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606256979
transform 1 0 13340 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606256979
transform 1 0 14076 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606256979
transform 1 0 13340 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1606256979
transform 1 0 12972 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_137
timestamp 1606256979
transform 1 0 13708 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_145
timestamp 1606256979
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_129
timestamp 1606256979
transform 1 0 12972 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1606256979
transform 1 0 13708 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 15824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 15824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1606256979
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_149
timestamp 1606256979
transform 1 0 14812 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1606256979
transform 1 0 15456 0 1 16864
box -38 -48 130 592
<< labels >>
rlabel metal3 s 16520 16600 17000 16720 6 Test_en_E_in
port 0 nsew default input
rlabel metal3 s 16520 9936 17000 10056 6 Test_en_E_out
port 1 nsew default tristate
rlabel metal2 s 3146 19520 3202 20000 6 Test_en_N_out
port 2 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 Test_en_S_in
port 3 nsew default input
rlabel metal3 s 0 17280 480 17400 6 Test_en_W_in
port 4 nsew default input
rlabel metal3 s 0 18368 480 18488 6 Test_en_W_out
port 5 nsew default tristate
rlabel metal3 s 0 416 480 536 6 ccff_head
port 6 nsew default input
rlabel metal3 s 16520 3272 17000 3392 6 ccff_tail
port 7 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[0]
port 8 nsew default input
rlabel metal2 s 10322 0 10378 480 6 chany_bottom_in[10]
port 9 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[11]
port 10 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[12]
port 11 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[13]
port 12 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_in[14]
port 13 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[15]
port 14 nsew default input
rlabel metal2 s 12346 0 12402 480 6 chany_bottom_in[16]
port 15 nsew default input
rlabel metal2 s 12622 0 12678 480 6 chany_bottom_in[17]
port 16 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[18]
port 17 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[19]
port 18 nsew default input
rlabel metal2 s 7194 0 7250 480 6 chany_bottom_in[1]
port 19 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[2]
port 20 nsew default input
rlabel metal2 s 7930 0 7986 480 6 chany_bottom_in[3]
port 21 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[4]
port 22 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[5]
port 23 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[6]
port 24 nsew default input
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_in[7]
port 25 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_in[8]
port 26 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[9]
port 27 nsew default input
rlabel metal2 s 110 0 166 480 6 chany_bottom_out[0]
port 28 nsew default tristate
rlabel metal2 s 3514 0 3570 480 6 chany_bottom_out[10]
port 29 nsew default tristate
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_out[11]
port 30 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_out[12]
port 31 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_out[13]
port 32 nsew default tristate
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_out[14]
port 33 nsew default tristate
rlabel metal2 s 5170 0 5226 480 6 chany_bottom_out[15]
port 34 nsew default tristate
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_out[16]
port 35 nsew default tristate
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_out[17]
port 36 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_out[18]
port 37 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[19]
port 38 nsew default tristate
rlabel metal2 s 386 0 442 480 6 chany_bottom_out[1]
port 39 nsew default tristate
rlabel metal2 s 754 0 810 480 6 chany_bottom_out[2]
port 40 nsew default tristate
rlabel metal2 s 1122 0 1178 480 6 chany_bottom_out[3]
port 41 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[4]
port 42 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_out[5]
port 43 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_out[6]
port 44 nsew default tristate
rlabel metal2 s 2410 0 2466 480 6 chany_bottom_out[7]
port 45 nsew default tristate
rlabel metal2 s 2778 0 2834 480 6 chany_bottom_out[8]
port 46 nsew default tristate
rlabel metal2 s 3146 0 3202 480 6 chany_bottom_out[9]
port 47 nsew default tristate
rlabel metal2 s 10322 19520 10378 20000 6 chany_top_in[0]
port 48 nsew default input
rlabel metal2 s 13726 19520 13782 20000 6 chany_top_in[10]
port 49 nsew default input
rlabel metal2 s 14002 19520 14058 20000 6 chany_top_in[11]
port 50 nsew default input
rlabel metal2 s 14370 19520 14426 20000 6 chany_top_in[12]
port 51 nsew default input
rlabel metal2 s 14738 19520 14794 20000 6 chany_top_in[13]
port 52 nsew default input
rlabel metal2 s 15014 19520 15070 20000 6 chany_top_in[14]
port 53 nsew default input
rlabel metal2 s 15382 19520 15438 20000 6 chany_top_in[15]
port 54 nsew default input
rlabel metal2 s 15750 19520 15806 20000 6 chany_top_in[16]
port 55 nsew default input
rlabel metal2 s 16026 19520 16082 20000 6 chany_top_in[17]
port 56 nsew default input
rlabel metal2 s 16394 19520 16450 20000 6 chany_top_in[18]
port 57 nsew default input
rlabel metal2 s 16762 19520 16818 20000 6 chany_top_in[19]
port 58 nsew default input
rlabel metal2 s 10598 19520 10654 20000 6 chany_top_in[1]
port 59 nsew default input
rlabel metal2 s 10966 19520 11022 20000 6 chany_top_in[2]
port 60 nsew default input
rlabel metal2 s 11334 19520 11390 20000 6 chany_top_in[3]
port 61 nsew default input
rlabel metal2 s 11610 19520 11666 20000 6 chany_top_in[4]
port 62 nsew default input
rlabel metal2 s 11978 19520 12034 20000 6 chany_top_in[5]
port 63 nsew default input
rlabel metal2 s 12346 19520 12402 20000 6 chany_top_in[6]
port 64 nsew default input
rlabel metal2 s 12622 19520 12678 20000 6 chany_top_in[7]
port 65 nsew default input
rlabel metal2 s 12990 19520 13046 20000 6 chany_top_in[8]
port 66 nsew default input
rlabel metal2 s 13358 19520 13414 20000 6 chany_top_in[9]
port 67 nsew default input
rlabel metal2 s 3514 19520 3570 20000 6 chany_top_out[0]
port 68 nsew default tristate
rlabel metal2 s 6918 19520 6974 20000 6 chany_top_out[10]
port 69 nsew default tristate
rlabel metal2 s 7194 19520 7250 20000 6 chany_top_out[11]
port 70 nsew default tristate
rlabel metal2 s 7562 19520 7618 20000 6 chany_top_out[12]
port 71 nsew default tristate
rlabel metal2 s 7930 19520 7986 20000 6 chany_top_out[13]
port 72 nsew default tristate
rlabel metal2 s 8206 19520 8262 20000 6 chany_top_out[14]
port 73 nsew default tristate
rlabel metal2 s 8574 19520 8630 20000 6 chany_top_out[15]
port 74 nsew default tristate
rlabel metal2 s 8942 19520 8998 20000 6 chany_top_out[16]
port 75 nsew default tristate
rlabel metal2 s 9218 19520 9274 20000 6 chany_top_out[17]
port 76 nsew default tristate
rlabel metal2 s 9586 19520 9642 20000 6 chany_top_out[18]
port 77 nsew default tristate
rlabel metal2 s 9954 19520 10010 20000 6 chany_top_out[19]
port 78 nsew default tristate
rlabel metal2 s 3790 19520 3846 20000 6 chany_top_out[1]
port 79 nsew default tristate
rlabel metal2 s 4158 19520 4214 20000 6 chany_top_out[2]
port 80 nsew default tristate
rlabel metal2 s 4526 19520 4582 20000 6 chany_top_out[3]
port 81 nsew default tristate
rlabel metal2 s 4802 19520 4858 20000 6 chany_top_out[4]
port 82 nsew default tristate
rlabel metal2 s 5170 19520 5226 20000 6 chany_top_out[5]
port 83 nsew default tristate
rlabel metal2 s 5538 19520 5594 20000 6 chany_top_out[6]
port 84 nsew default tristate
rlabel metal2 s 5814 19520 5870 20000 6 chany_top_out[7]
port 85 nsew default tristate
rlabel metal2 s 6182 19520 6238 20000 6 chany_top_out[8]
port 86 nsew default tristate
rlabel metal2 s 6550 19520 6606 20000 6 chany_top_out[9]
port 87 nsew default tristate
rlabel metal2 s 110 19520 166 20000 6 clk_2_N_in
port 88 nsew default input
rlabel metal2 s 1398 19520 1454 20000 6 clk_2_N_out
port 89 nsew default tristate
rlabel metal2 s 14002 0 14058 480 6 clk_2_S_in
port 90 nsew default input
rlabel metal2 s 15382 0 15438 480 6 clk_2_S_out
port 91 nsew default tristate
rlabel metal2 s 386 19520 442 20000 6 clk_3_N_in
port 92 nsew default input
rlabel metal2 s 1766 19520 1822 20000 6 clk_3_N_out
port 93 nsew default tristate
rlabel metal2 s 14370 0 14426 480 6 clk_3_S_in
port 94 nsew default input
rlabel metal2 s 15750 0 15806 480 6 clk_3_S_out
port 95 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 left_grid_pin_16_
port 96 nsew default tristate
rlabel metal3 s 0 2320 480 2440 6 left_grid_pin_17_
port 97 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 left_grid_pin_18_
port 98 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 left_grid_pin_19_
port 99 nsew default tristate
rlabel metal3 s 0 5312 480 5432 6 left_grid_pin_20_
port 100 nsew default tristate
rlabel metal3 s 0 6400 480 6520 6 left_grid_pin_21_
port 101 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 left_grid_pin_22_
port 102 nsew default tristate
rlabel metal3 s 0 8304 480 8424 6 left_grid_pin_23_
port 103 nsew default tristate
rlabel metal3 s 0 9392 480 9512 6 left_grid_pin_24_
port 104 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 left_grid_pin_25_
port 105 nsew default tristate
rlabel metal3 s 0 11296 480 11416 6 left_grid_pin_26_
port 106 nsew default tristate
rlabel metal3 s 0 12384 480 12504 6 left_grid_pin_27_
port 107 nsew default tristate
rlabel metal3 s 0 13336 480 13456 6 left_grid_pin_28_
port 108 nsew default tristate
rlabel metal3 s 0 14288 480 14408 6 left_grid_pin_29_
port 109 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 left_grid_pin_30_
port 110 nsew default tristate
rlabel metal3 s 0 16328 480 16448 6 left_grid_pin_31_
port 111 nsew default tristate
rlabel metal2 s 2134 19520 2190 20000 6 prog_clk_0_N_out
port 112 nsew default tristate
rlabel metal2 s 16026 0 16082 480 6 prog_clk_0_S_out
port 113 nsew default tristate
rlabel metal3 s 0 19320 480 19440 6 prog_clk_0_W_in
port 114 nsew default input
rlabel metal2 s 754 19520 810 20000 6 prog_clk_2_N_in
port 115 nsew default input
rlabel metal2 s 2410 19520 2466 20000 6 prog_clk_2_N_out
port 116 nsew default tristate
rlabel metal2 s 14738 0 14794 480 6 prog_clk_2_S_in
port 117 nsew default input
rlabel metal2 s 16394 0 16450 480 6 prog_clk_2_S_out
port 118 nsew default tristate
rlabel metal2 s 1122 19520 1178 20000 6 prog_clk_3_N_in
port 119 nsew default input
rlabel metal2 s 2778 19520 2834 20000 6 prog_clk_3_N_out
port 120 nsew default tristate
rlabel metal2 s 15014 0 15070 480 6 prog_clk_3_S_in
port 121 nsew default input
rlabel metal2 s 16762 0 16818 480 6 prog_clk_3_S_out
port 122 nsew default tristate
rlabel metal4 s 3409 2128 3729 17456 6 VPWR
port 123 nsew default input
rlabel metal4 s 5875 2128 6195 17456 6 VGND
port 124 nsew default input
<< properties >>
string FIXED_BBOX 0 0 17000 20000
<< end >>
