magic
tech sky130A
magscale 1 2
timestamp 1608157412
<< obsli1 >>
rect 1104 2159 21620 20145
<< obsm1 >>
rect 198 552 22618 20732
<< metal2 >>
rect 202 22000 258 22800
rect 570 22000 626 22800
rect 1030 22000 1086 22800
rect 1490 22000 1546 22800
rect 1950 22000 2006 22800
rect 2410 22000 2466 22800
rect 2870 22000 2926 22800
rect 3330 22000 3386 22800
rect 3790 22000 3846 22800
rect 4250 22000 4306 22800
rect 4710 22000 4766 22800
rect 5170 22000 5226 22800
rect 5630 22000 5686 22800
rect 6090 22000 6146 22800
rect 6550 22000 6606 22800
rect 7010 22000 7066 22800
rect 7470 22000 7526 22800
rect 7930 22000 7986 22800
rect 8390 22000 8446 22800
rect 8850 22000 8906 22800
rect 9310 22000 9366 22800
rect 9770 22000 9826 22800
rect 10230 22000 10286 22800
rect 10690 22000 10746 22800
rect 11150 22000 11206 22800
rect 11610 22000 11666 22800
rect 11978 22000 12034 22800
rect 12438 22000 12494 22800
rect 12898 22000 12954 22800
rect 13358 22000 13414 22800
rect 13818 22000 13874 22800
rect 14278 22000 14334 22800
rect 14738 22000 14794 22800
rect 15198 22000 15254 22800
rect 15658 22000 15714 22800
rect 16118 22000 16174 22800
rect 16578 22000 16634 22800
rect 17038 22000 17094 22800
rect 17498 22000 17554 22800
rect 17958 22000 18014 22800
rect 18418 22000 18474 22800
rect 18878 22000 18934 22800
rect 19338 22000 19394 22800
rect 19798 22000 19854 22800
rect 20258 22000 20314 22800
rect 20718 22000 20774 22800
rect 21178 22000 21234 22800
rect 21638 22000 21694 22800
rect 22098 22000 22154 22800
rect 22558 22000 22614 22800
rect 11426 0 11482 800
<< obsm2 >>
rect 314 21944 514 22545
rect 682 21944 974 22545
rect 1142 21944 1434 22545
rect 1602 21944 1894 22545
rect 2062 21944 2354 22545
rect 2522 21944 2814 22545
rect 2982 21944 3274 22545
rect 3442 21944 3734 22545
rect 3902 21944 4194 22545
rect 4362 21944 4654 22545
rect 4822 21944 5114 22545
rect 5282 21944 5574 22545
rect 5742 21944 6034 22545
rect 6202 21944 6494 22545
rect 6662 21944 6954 22545
rect 7122 21944 7414 22545
rect 7582 21944 7874 22545
rect 8042 21944 8334 22545
rect 8502 21944 8794 22545
rect 8962 21944 9254 22545
rect 9422 21944 9714 22545
rect 9882 21944 10174 22545
rect 10342 21944 10634 22545
rect 10802 21944 11094 22545
rect 11262 21944 11554 22545
rect 11722 21944 11922 22545
rect 12090 21944 12382 22545
rect 12550 21944 12842 22545
rect 13010 21944 13302 22545
rect 13470 21944 13762 22545
rect 13930 21944 14222 22545
rect 14390 21944 14682 22545
rect 14850 21944 15142 22545
rect 15310 21944 15602 22545
rect 15770 21944 16062 22545
rect 16230 21944 16522 22545
rect 16690 21944 16982 22545
rect 17150 21944 17442 22545
rect 17610 21944 17902 22545
rect 18070 21944 18362 22545
rect 18530 21944 18822 22545
rect 18990 21944 19282 22545
rect 19450 21944 19742 22545
rect 19910 21944 20202 22545
rect 20370 21944 20662 22545
rect 20830 21944 21122 22545
rect 21290 21944 21582 22545
rect 21750 21944 22042 22545
rect 22210 21944 22502 22545
rect 204 856 22612 21944
rect 204 167 11370 856
rect 11538 167 22612 856
<< metal3 >>
rect 0 22448 800 22568
rect 0 22040 800 22160
rect 0 21496 800 21616
rect 0 21088 800 21208
rect 0 20544 800 20664
rect 0 20136 800 20256
rect 0 19728 800 19848
rect 0 19184 800 19304
rect 0 18776 800 18896
rect 0 18232 800 18352
rect 0 17824 800 17944
rect 0 17280 800 17400
rect 0 16872 800 16992
rect 0 16464 800 16584
rect 0 15920 800 16040
rect 0 15512 800 15632
rect 0 14968 800 15088
rect 0 14560 800 14680
rect 0 14016 800 14136
rect 0 13608 800 13728
rect 0 13200 800 13320
rect 0 12656 800 12776
rect 0 12248 800 12368
rect 0 11704 800 11824
rect 0 11296 800 11416
rect 22000 11432 22800 11552
rect 0 10752 800 10872
rect 0 10344 800 10464
rect 0 9936 800 10056
rect 0 9392 800 9512
rect 0 8984 800 9104
rect 0 8440 800 8560
rect 0 8032 800 8152
rect 0 7488 800 7608
rect 0 7080 800 7200
rect 0 6672 800 6792
rect 0 6128 800 6248
rect 0 5720 800 5840
rect 0 5176 800 5296
rect 0 4768 800 4888
rect 0 4224 800 4344
rect 0 3816 800 3936
rect 0 3408 800 3528
rect 0 2864 800 2984
rect 0 2456 800 2576
rect 0 1912 800 2032
rect 0 1504 800 1624
rect 0 960 800 1080
rect 0 552 800 672
rect 0 144 800 264
<< obsm3 >>
rect 880 22368 22000 22541
rect 800 22240 22000 22368
rect 880 21960 22000 22240
rect 800 21696 22000 21960
rect 880 21416 22000 21696
rect 800 21288 22000 21416
rect 880 21008 22000 21288
rect 800 20744 22000 21008
rect 880 20464 22000 20744
rect 800 20336 22000 20464
rect 880 20056 22000 20336
rect 800 19928 22000 20056
rect 880 19648 22000 19928
rect 800 19384 22000 19648
rect 880 19104 22000 19384
rect 800 18976 22000 19104
rect 880 18696 22000 18976
rect 800 18432 22000 18696
rect 880 18152 22000 18432
rect 800 18024 22000 18152
rect 880 17744 22000 18024
rect 800 17480 22000 17744
rect 880 17200 22000 17480
rect 800 17072 22000 17200
rect 880 16792 22000 17072
rect 800 16664 22000 16792
rect 880 16384 22000 16664
rect 800 16120 22000 16384
rect 880 15840 22000 16120
rect 800 15712 22000 15840
rect 880 15432 22000 15712
rect 800 15168 22000 15432
rect 880 14888 22000 15168
rect 800 14760 22000 14888
rect 880 14480 22000 14760
rect 800 14216 22000 14480
rect 880 13936 22000 14216
rect 800 13808 22000 13936
rect 880 13528 22000 13808
rect 800 13400 22000 13528
rect 880 13120 22000 13400
rect 800 12856 22000 13120
rect 880 12576 22000 12856
rect 800 12448 22000 12576
rect 880 12168 22000 12448
rect 800 11904 22000 12168
rect 880 11632 22000 11904
rect 880 11624 21920 11632
rect 800 11496 21920 11624
rect 880 11352 21920 11496
rect 880 11216 22000 11352
rect 800 10952 22000 11216
rect 880 10672 22000 10952
rect 800 10544 22000 10672
rect 880 10264 22000 10544
rect 800 10136 22000 10264
rect 880 9856 22000 10136
rect 800 9592 22000 9856
rect 880 9312 22000 9592
rect 800 9184 22000 9312
rect 880 8904 22000 9184
rect 800 8640 22000 8904
rect 880 8360 22000 8640
rect 800 8232 22000 8360
rect 880 7952 22000 8232
rect 800 7688 22000 7952
rect 880 7408 22000 7688
rect 800 7280 22000 7408
rect 880 7000 22000 7280
rect 800 6872 22000 7000
rect 880 6592 22000 6872
rect 800 6328 22000 6592
rect 880 6048 22000 6328
rect 800 5920 22000 6048
rect 880 5640 22000 5920
rect 800 5376 22000 5640
rect 880 5096 22000 5376
rect 800 4968 22000 5096
rect 880 4688 22000 4968
rect 800 4424 22000 4688
rect 880 4144 22000 4424
rect 800 4016 22000 4144
rect 880 3736 22000 4016
rect 800 3608 22000 3736
rect 880 3328 22000 3608
rect 800 3064 22000 3328
rect 880 2784 22000 3064
rect 800 2656 22000 2784
rect 880 2376 22000 2656
rect 800 2112 22000 2376
rect 880 1832 22000 2112
rect 800 1704 22000 1832
rect 880 1424 22000 1704
rect 800 1160 22000 1424
rect 880 880 22000 1160
rect 800 752 22000 880
rect 880 472 22000 752
rect 800 344 22000 472
rect 880 171 22000 344
<< metal4 >>
rect 4376 2128 4696 20176
rect 7808 2128 8128 20176
<< obsm4 >>
rect 11240 2128 18424 20176
<< labels >>
rlabel metal3 s 22000 11432 22800 11552 6 ccff_head
port 1 nsew default input
rlabel metal2 s 11426 0 11482 800 6 ccff_tail
port 2 nsew default output
rlabel metal3 s 0 4224 800 4344 6 chanx_left_in[0]
port 3 nsew default input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[10]
port 4 nsew default input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[11]
port 5 nsew default input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[12]
port 6 nsew default input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[13]
port 7 nsew default input
rlabel metal3 s 0 10752 800 10872 6 chanx_left_in[14]
port 8 nsew default input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[15]
port 9 nsew default input
rlabel metal3 s 0 11704 800 11824 6 chanx_left_in[16]
port 10 nsew default input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 11 nsew default input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[18]
port 12 nsew default input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_in[19]
port 13 nsew default input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[1]
port 14 nsew default input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[2]
port 15 nsew default input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[3]
port 16 nsew default input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[4]
port 17 nsew default input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[5]
port 18 nsew default input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[6]
port 19 nsew default input
rlabel metal3 s 0 7488 800 7608 6 chanx_left_in[7]
port 20 nsew default input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[8]
port 21 nsew default input
rlabel metal3 s 0 8440 800 8560 6 chanx_left_in[9]
port 22 nsew default input
rlabel metal3 s 0 13608 800 13728 6 chanx_left_out[0]
port 23 nsew default output
rlabel metal3 s 0 18232 800 18352 6 chanx_left_out[10]
port 24 nsew default output
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[11]
port 25 nsew default output
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[12]
port 26 nsew default output
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[13]
port 27 nsew default output
rlabel metal3 s 0 20136 800 20256 6 chanx_left_out[14]
port 28 nsew default output
rlabel metal3 s 0 20544 800 20664 6 chanx_left_out[15]
port 29 nsew default output
rlabel metal3 s 0 21088 800 21208 6 chanx_left_out[16]
port 30 nsew default output
rlabel metal3 s 0 21496 800 21616 6 chanx_left_out[17]
port 31 nsew default output
rlabel metal3 s 0 22040 800 22160 6 chanx_left_out[18]
port 32 nsew default output
rlabel metal3 s 0 22448 800 22568 6 chanx_left_out[19]
port 33 nsew default output
rlabel metal3 s 0 14016 800 14136 6 chanx_left_out[1]
port 34 nsew default output
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[2]
port 35 nsew default output
rlabel metal3 s 0 14968 800 15088 6 chanx_left_out[3]
port 36 nsew default output
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[4]
port 37 nsew default output
rlabel metal3 s 0 15920 800 16040 6 chanx_left_out[5]
port 38 nsew default output
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[6]
port 39 nsew default output
rlabel metal3 s 0 16872 800 16992 6 chanx_left_out[7]
port 40 nsew default output
rlabel metal3 s 0 17280 800 17400 6 chanx_left_out[8]
port 41 nsew default output
rlabel metal3 s 0 17824 800 17944 6 chanx_left_out[9]
port 42 nsew default output
rlabel metal2 s 3790 22000 3846 22800 6 chany_top_in[0]
port 43 nsew default input
rlabel metal2 s 8390 22000 8446 22800 6 chany_top_in[10]
port 44 nsew default input
rlabel metal2 s 8850 22000 8906 22800 6 chany_top_in[11]
port 45 nsew default input
rlabel metal2 s 9310 22000 9366 22800 6 chany_top_in[12]
port 46 nsew default input
rlabel metal2 s 9770 22000 9826 22800 6 chany_top_in[13]
port 47 nsew default input
rlabel metal2 s 10230 22000 10286 22800 6 chany_top_in[14]
port 48 nsew default input
rlabel metal2 s 10690 22000 10746 22800 6 chany_top_in[15]
port 49 nsew default input
rlabel metal2 s 11150 22000 11206 22800 6 chany_top_in[16]
port 50 nsew default input
rlabel metal2 s 11610 22000 11666 22800 6 chany_top_in[17]
port 51 nsew default input
rlabel metal2 s 11978 22000 12034 22800 6 chany_top_in[18]
port 52 nsew default input
rlabel metal2 s 12438 22000 12494 22800 6 chany_top_in[19]
port 53 nsew default input
rlabel metal2 s 4250 22000 4306 22800 6 chany_top_in[1]
port 54 nsew default input
rlabel metal2 s 4710 22000 4766 22800 6 chany_top_in[2]
port 55 nsew default input
rlabel metal2 s 5170 22000 5226 22800 6 chany_top_in[3]
port 56 nsew default input
rlabel metal2 s 5630 22000 5686 22800 6 chany_top_in[4]
port 57 nsew default input
rlabel metal2 s 6090 22000 6146 22800 6 chany_top_in[5]
port 58 nsew default input
rlabel metal2 s 6550 22000 6606 22800 6 chany_top_in[6]
port 59 nsew default input
rlabel metal2 s 7010 22000 7066 22800 6 chany_top_in[7]
port 60 nsew default input
rlabel metal2 s 7470 22000 7526 22800 6 chany_top_in[8]
port 61 nsew default input
rlabel metal2 s 7930 22000 7986 22800 6 chany_top_in[9]
port 62 nsew default input
rlabel metal2 s 12898 22000 12954 22800 6 chany_top_out[0]
port 63 nsew default output
rlabel metal2 s 17498 22000 17554 22800 6 chany_top_out[10]
port 64 nsew default output
rlabel metal2 s 17958 22000 18014 22800 6 chany_top_out[11]
port 65 nsew default output
rlabel metal2 s 18418 22000 18474 22800 6 chany_top_out[12]
port 66 nsew default output
rlabel metal2 s 18878 22000 18934 22800 6 chany_top_out[13]
port 67 nsew default output
rlabel metal2 s 19338 22000 19394 22800 6 chany_top_out[14]
port 68 nsew default output
rlabel metal2 s 19798 22000 19854 22800 6 chany_top_out[15]
port 69 nsew default output
rlabel metal2 s 20258 22000 20314 22800 6 chany_top_out[16]
port 70 nsew default output
rlabel metal2 s 20718 22000 20774 22800 6 chany_top_out[17]
port 71 nsew default output
rlabel metal2 s 21178 22000 21234 22800 6 chany_top_out[18]
port 72 nsew default output
rlabel metal2 s 21638 22000 21694 22800 6 chany_top_out[19]
port 73 nsew default output
rlabel metal2 s 13358 22000 13414 22800 6 chany_top_out[1]
port 74 nsew default output
rlabel metal2 s 13818 22000 13874 22800 6 chany_top_out[2]
port 75 nsew default output
rlabel metal2 s 14278 22000 14334 22800 6 chany_top_out[3]
port 76 nsew default output
rlabel metal2 s 14738 22000 14794 22800 6 chany_top_out[4]
port 77 nsew default output
rlabel metal2 s 15198 22000 15254 22800 6 chany_top_out[5]
port 78 nsew default output
rlabel metal2 s 15658 22000 15714 22800 6 chany_top_out[6]
port 79 nsew default output
rlabel metal2 s 16118 22000 16174 22800 6 chany_top_out[7]
port 80 nsew default output
rlabel metal2 s 16578 22000 16634 22800 6 chany_top_out[8]
port 81 nsew default output
rlabel metal2 s 17038 22000 17094 22800 6 chany_top_out[9]
port 82 nsew default output
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_11_
port 83 nsew default input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_13_
port 84 nsew default input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_15_
port 85 nsew default input
rlabel metal3 s 0 3816 800 3936 6 left_bottom_grid_pin_17_
port 86 nsew default input
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_1_
port 87 nsew default input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_3_
port 88 nsew default input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_5_
port 89 nsew default input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_7_
port 90 nsew default input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_9_
port 91 nsew default input
rlabel metal2 s 22098 22000 22154 22800 6 prog_clk_0_N_in
port 92 nsew default input
rlabel metal2 s 202 22000 258 22800 6 top_left_grid_pin_42_
port 93 nsew default input
rlabel metal2 s 570 22000 626 22800 6 top_left_grid_pin_43_
port 94 nsew default input
rlabel metal2 s 1030 22000 1086 22800 6 top_left_grid_pin_44_
port 95 nsew default input
rlabel metal2 s 1490 22000 1546 22800 6 top_left_grid_pin_45_
port 96 nsew default input
rlabel metal2 s 1950 22000 2006 22800 6 top_left_grid_pin_46_
port 97 nsew default input
rlabel metal2 s 2410 22000 2466 22800 6 top_left_grid_pin_47_
port 98 nsew default input
rlabel metal2 s 2870 22000 2926 22800 6 top_left_grid_pin_48_
port 99 nsew default input
rlabel metal2 s 3330 22000 3386 22800 6 top_left_grid_pin_49_
port 100 nsew default input
rlabel metal2 s 22558 22000 22614 22800 6 top_right_grid_pin_1_
port 101 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 102 nsew power input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 103 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22800 22800
string LEFview TRUE
<< end >>
