magic
tech EFS8A
magscale 1 2
timestamp 1603297939
<< locali >>
rect 10051 34153 10057 34187
rect 10051 34085 10085 34153
rect 5215 34017 5250 34051
rect 7205 33371 7239 33609
rect 7107 33065 7113 33099
rect 10051 33065 10057 33099
rect 7107 32997 7141 33065
rect 10051 32997 10085 33065
rect 13035 32929 13070 32963
rect 7199 32215 7233 32283
rect 7199 32181 7205 32215
rect 11287 31841 11322 31875
rect 10235 30039 10269 30107
rect 10235 30005 10241 30039
rect 8027 28713 8033 28747
rect 8027 28645 8061 28713
rect 4847 28577 4882 28611
rect 7849 27931 7883 28101
rect 13599 27081 13737 27115
rect 5267 25449 5273 25483
rect 10419 25449 10425 25483
rect 5267 25381 5301 25449
rect 10419 25381 10453 25449
rect 13587 25313 13622 25347
rect 12667 24225 12702 24259
rect 11897 24055 11931 24157
rect 6561 22491 6595 22729
rect 10419 22185 10425 22219
rect 10419 22117 10453 22185
rect 4203 21437 4295 21471
rect 10609 19295 10643 19465
rect 4623 19159 4657 19227
rect 4623 19125 4629 19159
rect 3111 18921 3249 18955
rect 1995 18785 2030 18819
rect 2915 18785 3042 18819
rect 13587 16609 13622 16643
rect 11471 13345 11506 13379
rect 7199 12631 7233 12699
rect 7199 12597 7205 12631
rect 4623 11305 4629 11339
rect 4623 11237 4657 11305
rect 2881 10081 3042 10115
rect 9631 10081 9758 10115
rect 2881 9911 2915 10081
rect 1501 2975 1535 3145
rect 1501 2941 1662 2975
<< viali >>
rect 9664 36669 9698 36703
rect 10057 36669 10091 36703
rect 9735 36533 9769 36567
rect 8677 36329 8711 36363
rect 7548 36193 7582 36227
rect 8493 36193 8527 36227
rect 9724 36193 9758 36227
rect 7619 35989 7653 36023
rect 8217 35989 8251 36023
rect 9827 35989 9861 36023
rect 10241 35989 10275 36023
rect 7021 35785 7055 35819
rect 7849 35717 7883 35751
rect 8309 35649 8343 35683
rect 9229 35649 9263 35683
rect 9689 35649 9723 35683
rect 10333 35649 10367 35683
rect 6837 35581 6871 35615
rect 7389 35581 7423 35615
rect 8401 35513 8435 35547
rect 8953 35513 8987 35547
rect 10149 35513 10183 35547
rect 10425 35513 10459 35547
rect 10977 35513 11011 35547
rect 7113 35241 7147 35275
rect 9045 35241 9079 35275
rect 10241 35241 10275 35275
rect 13185 35241 13219 35275
rect 6055 35173 6089 35207
rect 8217 35173 8251 35207
rect 10609 35173 10643 35207
rect 5968 35105 6002 35139
rect 6929 35105 6963 35139
rect 12056 35105 12090 35139
rect 13001 35105 13035 35139
rect 8125 35037 8159 35071
rect 8401 35037 8435 35071
rect 10517 35037 10551 35071
rect 11161 35037 11195 35071
rect 7665 34901 7699 34935
rect 12127 34901 12161 34935
rect 5825 34697 5859 34731
rect 9321 34697 9355 34731
rect 12633 34697 12667 34731
rect 12081 34629 12115 34663
rect 8309 34561 8343 34595
rect 10333 34561 10367 34595
rect 10977 34561 11011 34595
rect 13093 34561 13127 34595
rect 5641 34493 5675 34527
rect 6193 34493 6227 34527
rect 9137 34493 9171 34527
rect 9689 34493 9723 34527
rect 12449 34493 12483 34527
rect 13369 34493 13403 34527
rect 7665 34425 7699 34459
rect 7757 34425 7791 34459
rect 8953 34425 8987 34459
rect 10425 34425 10459 34459
rect 6653 34357 6687 34391
rect 7021 34357 7055 34391
rect 7481 34357 7515 34391
rect 8677 34357 8711 34391
rect 10149 34357 10183 34391
rect 11253 34357 11287 34391
rect 5319 34153 5353 34187
rect 10057 34153 10091 34187
rect 13185 34153 13219 34187
rect 6377 34085 6411 34119
rect 7941 34085 7975 34119
rect 8493 34085 8527 34119
rect 11621 34085 11655 34119
rect 5181 34017 5215 34051
rect 10609 34017 10643 34051
rect 13001 34017 13035 34051
rect 6285 33949 6319 33983
rect 7849 33949 7883 33983
rect 9689 33949 9723 33983
rect 11529 33949 11563 33983
rect 11805 33949 11839 33983
rect 6837 33881 6871 33915
rect 7573 33813 7607 33847
rect 10977 33813 11011 33847
rect 4859 33609 4893 33643
rect 6561 33609 6595 33643
rect 7205 33609 7239 33643
rect 7297 33609 7331 33643
rect 10241 33609 10275 33643
rect 10977 33609 11011 33643
rect 11253 33609 11287 33643
rect 13461 33609 13495 33643
rect 5871 33473 5905 33507
rect 4788 33405 4822 33439
rect 5784 33405 5818 33439
rect 12173 33541 12207 33575
rect 7573 33473 7607 33507
rect 8217 33473 8251 33507
rect 8861 33473 8895 33507
rect 12541 33473 12575 33507
rect 12817 33473 12851 33507
rect 9321 33405 9355 33439
rect 11069 33405 11103 33439
rect 7205 33337 7239 33371
rect 7665 33337 7699 33371
rect 9683 33337 9717 33371
rect 10517 33337 10551 33371
rect 11713 33337 11747 33371
rect 12633 33337 12667 33371
rect 5273 33269 5307 33303
rect 5641 33269 5675 33303
rect 6285 33269 6319 33303
rect 9229 33269 9263 33303
rect 5871 33065 5905 33099
rect 6193 33065 6227 33099
rect 7113 33065 7147 33099
rect 7665 33065 7699 33099
rect 7941 33065 7975 33099
rect 10057 33065 10091 33099
rect 10609 33065 10643 33099
rect 12541 33065 12575 33099
rect 8309 32997 8343 33031
rect 8631 32997 8665 33031
rect 11621 32997 11655 33031
rect 12173 32997 12207 33031
rect 5768 32929 5802 32963
rect 8528 32929 8562 32963
rect 13001 32929 13035 32963
rect 6745 32861 6779 32895
rect 9689 32861 9723 32895
rect 11529 32861 11563 32895
rect 8953 32725 8987 32759
rect 9321 32725 9355 32759
rect 11345 32725 11379 32759
rect 13139 32725 13173 32759
rect 5733 32521 5767 32555
rect 7757 32521 7791 32555
rect 8401 32521 8435 32555
rect 9505 32521 9539 32555
rect 11713 32521 11747 32555
rect 12587 32521 12621 32555
rect 12265 32453 12299 32487
rect 6285 32385 6319 32419
rect 6653 32385 6687 32419
rect 8585 32385 8619 32419
rect 6837 32317 6871 32351
rect 10333 32317 10367 32351
rect 10793 32317 10827 32351
rect 12484 32317 12518 32351
rect 8125 32249 8159 32283
rect 8947 32249 8981 32283
rect 10241 32249 10275 32283
rect 7205 32181 7239 32215
rect 9781 32181 9815 32215
rect 10425 32181 10459 32215
rect 11345 32181 11379 32215
rect 13001 32181 13035 32215
rect 9781 31977 9815 32011
rect 11391 31977 11425 32011
rect 11713 31977 11747 32011
rect 6837 31909 6871 31943
rect 7481 31909 7515 31943
rect 8401 31909 8435 31943
rect 6101 31841 6135 31875
rect 6653 31841 6687 31875
rect 7849 31841 7883 31875
rect 8125 31841 8159 31875
rect 9965 31841 9999 31875
rect 10241 31841 10275 31875
rect 11253 31841 11287 31875
rect 10701 31705 10735 31739
rect 7205 31637 7239 31671
rect 8677 31637 8711 31671
rect 9781 31433 9815 31467
rect 10149 31365 10183 31399
rect 7389 31297 7423 31331
rect 9321 31297 9355 31331
rect 10701 31297 10735 31331
rect 6929 31229 6963 31263
rect 7297 31229 7331 31263
rect 8677 31229 8711 31263
rect 9229 31229 9263 31263
rect 8585 31161 8619 31195
rect 10793 31161 10827 31195
rect 11345 31161 11379 31195
rect 5733 31093 5767 31127
rect 6193 31093 6227 31127
rect 6653 31093 6687 31127
rect 7849 31093 7883 31127
rect 10517 31093 10551 31127
rect 11713 31093 11747 31127
rect 7665 30889 7699 30923
rect 9413 30889 9447 30923
rect 10793 30889 10827 30923
rect 8125 30821 8159 30855
rect 8217 30821 8251 30855
rect 9873 30821 9907 30855
rect 11437 30821 11471 30855
rect 7021 30685 7055 30719
rect 8401 30685 8435 30719
rect 9781 30685 9815 30719
rect 10057 30685 10091 30719
rect 11345 30685 11379 30719
rect 11989 30685 12023 30719
rect 6929 30549 6963 30583
rect 8999 30345 9033 30379
rect 10793 30345 10827 30379
rect 11345 30345 11379 30379
rect 8769 30277 8803 30311
rect 11621 30209 11655 30243
rect 7481 30141 7515 30175
rect 7757 30141 7791 30175
rect 8928 30141 8962 30175
rect 9873 30141 9907 30175
rect 7113 30005 7147 30039
rect 7573 30005 7607 30039
rect 8309 30005 8343 30039
rect 9321 30005 9355 30039
rect 9781 30005 9815 30039
rect 10241 30005 10275 30039
rect 7481 29801 7515 29835
rect 7941 29801 7975 29835
rect 10977 29801 11011 29835
rect 10378 29733 10412 29767
rect 11989 29733 12023 29767
rect 6561 29665 6595 29699
rect 6929 29665 6963 29699
rect 8033 29665 8067 29699
rect 8585 29665 8619 29699
rect 7205 29597 7239 29631
rect 8769 29597 8803 29631
rect 9137 29597 9171 29631
rect 10057 29597 10091 29631
rect 11897 29597 11931 29631
rect 12173 29597 12207 29631
rect 5273 29461 5307 29495
rect 9965 29461 9999 29495
rect 8309 29257 8343 29291
rect 8677 29257 8711 29291
rect 10333 29257 10367 29291
rect 11897 29257 11931 29291
rect 5089 29121 5123 29155
rect 5273 29121 5307 29155
rect 5917 29121 5951 29155
rect 7389 29121 7423 29155
rect 9137 29121 9171 29155
rect 10885 29121 10919 29155
rect 7297 29053 7331 29087
rect 8953 29053 8987 29087
rect 10057 29053 10091 29087
rect 12173 29053 12207 29087
rect 5365 28985 5399 29019
rect 7751 28985 7785 29019
rect 9499 28985 9533 29019
rect 6561 28917 6595 28951
rect 10701 28917 10735 28951
rect 7481 28713 7515 28747
rect 8033 28713 8067 28747
rect 8585 28713 8619 28747
rect 9965 28713 9999 28747
rect 11437 28713 11471 28747
rect 4813 28577 4847 28611
rect 6193 28577 6227 28611
rect 6653 28577 6687 28611
rect 7665 28577 7699 28611
rect 9689 28577 9723 28611
rect 10149 28577 10183 28611
rect 11253 28577 11287 28611
rect 6837 28509 6871 28543
rect 8861 28441 8895 28475
rect 4951 28373 4985 28407
rect 5273 28373 5307 28407
rect 5641 28373 5675 28407
rect 7205 28373 7239 28407
rect 4445 28169 4479 28203
rect 4905 28169 4939 28203
rect 6193 28169 6227 28203
rect 8401 28169 8435 28203
rect 9137 28169 9171 28203
rect 10333 28169 10367 28203
rect 11069 28169 11103 28203
rect 7757 28101 7791 28135
rect 7849 28101 7883 28135
rect 8125 28101 8159 28135
rect 5089 28033 5123 28067
rect 6837 28033 6871 28067
rect 4020 27965 4054 27999
rect 8769 28033 8803 28067
rect 10057 28033 10091 28067
rect 9597 27965 9631 27999
rect 9781 27965 9815 27999
rect 10885 27965 10919 27999
rect 11713 27965 11747 27999
rect 5181 27897 5215 27931
rect 5733 27897 5767 27931
rect 6653 27897 6687 27931
rect 7199 27897 7233 27931
rect 7849 27897 7883 27931
rect 11345 27897 11379 27931
rect 4123 27829 4157 27863
rect 4813 27625 4847 27659
rect 5181 27625 5215 27659
rect 6745 27625 6779 27659
rect 4399 27557 4433 27591
rect 5457 27557 5491 27591
rect 7021 27557 7055 27591
rect 9873 27557 9907 27591
rect 11437 27557 11471 27591
rect 4312 27489 4346 27523
rect 8468 27489 8502 27523
rect 12884 27489 12918 27523
rect 5365 27421 5399 27455
rect 6929 27421 6963 27455
rect 9781 27421 9815 27455
rect 10425 27421 10459 27455
rect 11345 27421 11379 27455
rect 11621 27421 11655 27455
rect 5917 27353 5951 27387
rect 7481 27353 7515 27387
rect 6377 27285 6411 27319
rect 8539 27285 8573 27319
rect 9413 27285 9447 27319
rect 12955 27285 12989 27319
rect 3203 27081 3237 27115
rect 6285 27081 6319 27115
rect 7849 27081 7883 27115
rect 8539 27081 8573 27115
rect 13737 27081 13771 27115
rect 4537 27013 4571 27047
rect 7481 27013 7515 27047
rect 10241 27013 10275 27047
rect 5181 26945 5215 26979
rect 5825 26945 5859 26979
rect 6929 26945 6963 26979
rect 10977 26945 11011 26979
rect 3132 26877 3166 26911
rect 4128 26877 4162 26911
rect 6561 26877 6595 26911
rect 8436 26877 8470 26911
rect 9229 26877 9263 26911
rect 11196 26877 11230 26911
rect 11621 26877 11655 26911
rect 12484 26877 12518 26911
rect 12909 26877 12943 26911
rect 13496 26877 13530 26911
rect 4215 26809 4249 26843
rect 5273 26809 5307 26843
rect 7021 26809 7055 26843
rect 9689 26809 9723 26843
rect 9781 26809 9815 26843
rect 10609 26809 10643 26843
rect 13921 26809 13955 26843
rect 3525 26741 3559 26775
rect 4905 26741 4939 26775
rect 8861 26741 8895 26775
rect 11299 26741 11333 26775
rect 11989 26741 12023 26775
rect 12587 26741 12621 26775
rect 13277 26741 13311 26775
rect 5273 26537 5307 26571
rect 5641 26537 5675 26571
rect 5917 26537 5951 26571
rect 7113 26537 7147 26571
rect 12909 26537 12943 26571
rect 4674 26469 4708 26503
rect 6285 26469 6319 26503
rect 9873 26469 9907 26503
rect 11437 26469 11471 26503
rect 7849 26401 7883 26435
rect 8309 26401 8343 26435
rect 13093 26401 13127 26435
rect 13277 26401 13311 26435
rect 4353 26333 4387 26367
rect 6193 26333 6227 26367
rect 8401 26333 8435 26367
rect 9781 26333 9815 26367
rect 11345 26333 11379 26367
rect 6745 26265 6779 26299
rect 9137 26265 9171 26299
rect 10333 26265 10367 26299
rect 11897 26265 11931 26299
rect 7573 26197 7607 26231
rect 9505 26197 9539 26231
rect 10701 26197 10735 26231
rect 11161 26197 11195 26231
rect 12541 26197 12575 26231
rect 5181 25993 5215 26027
rect 6469 25993 6503 26027
rect 7481 25993 7515 26027
rect 9597 25993 9631 26027
rect 10977 25993 11011 26027
rect 11713 25993 11747 26027
rect 13461 25993 13495 26027
rect 7757 25925 7791 25959
rect 8217 25925 8251 25959
rect 9229 25925 9263 25959
rect 6975 25857 7009 25891
rect 8309 25857 8343 25891
rect 9965 25857 9999 25891
rect 12541 25857 12575 25891
rect 12817 25857 12851 25891
rect 3801 25789 3835 25823
rect 4261 25789 4295 25823
rect 6888 25789 6922 25823
rect 10057 25789 10091 25823
rect 4169 25721 4203 25755
rect 4582 25721 4616 25755
rect 8630 25721 8664 25755
rect 10378 25721 10412 25755
rect 11345 25721 11379 25755
rect 12633 25721 12667 25755
rect 5457 25653 5491 25687
rect 6101 25653 6135 25687
rect 12265 25653 12299 25687
rect 4353 25449 4387 25483
rect 5273 25449 5307 25483
rect 5825 25449 5859 25483
rect 8401 25449 8435 25483
rect 8953 25449 8987 25483
rect 9965 25449 9999 25483
rect 10425 25449 10459 25483
rect 10977 25449 11011 25483
rect 13001 25449 13035 25483
rect 7107 25381 7141 25415
rect 12126 25381 12160 25415
rect 2697 25313 2731 25347
rect 2881 25313 2915 25347
rect 3157 25313 3191 25347
rect 10057 25313 10091 25347
rect 12725 25313 12759 25347
rect 13553 25313 13587 25347
rect 4905 25245 4939 25279
rect 6745 25245 6779 25279
rect 8493 25245 8527 25279
rect 11805 25245 11839 25279
rect 13691 25177 13725 25211
rect 4721 25109 4755 25143
rect 6561 25109 6595 25143
rect 7665 25109 7699 25143
rect 7941 25109 7975 25143
rect 2513 24905 2547 24939
rect 2881 24905 2915 24939
rect 4997 24905 5031 24939
rect 6653 24905 6687 24939
rect 8217 24905 8251 24939
rect 10057 24905 10091 24939
rect 10425 24905 10459 24939
rect 11805 24905 11839 24939
rect 13553 24905 13587 24939
rect 4169 24769 4203 24803
rect 5917 24769 5951 24803
rect 7205 24769 7239 24803
rect 8861 24769 8895 24803
rect 9505 24769 9539 24803
rect 3617 24701 3651 24735
rect 4077 24701 4111 24735
rect 5457 24701 5491 24735
rect 5641 24701 5675 24735
rect 10517 24701 10551 24735
rect 12265 24701 12299 24735
rect 12725 24701 12759 24735
rect 12909 24701 12943 24735
rect 6285 24633 6319 24667
rect 7297 24633 7331 24667
rect 7849 24633 7883 24667
rect 8677 24633 8711 24667
rect 8953 24633 8987 24667
rect 10838 24633 10872 24667
rect 3433 24565 3467 24599
rect 11437 24565 11471 24599
rect 12541 24565 12575 24599
rect 10149 24361 10183 24395
rect 10977 24361 11011 24395
rect 4813 24293 4847 24327
rect 6561 24293 6595 24327
rect 7205 24293 7239 24327
rect 11253 24293 11287 24327
rect 2973 24225 3007 24259
rect 4077 24225 4111 24259
rect 4537 24225 4571 24259
rect 6009 24225 6043 24259
rect 8585 24225 8619 24259
rect 9689 24225 9723 24259
rect 10517 24225 10551 24259
rect 12633 24225 12667 24259
rect 7113 24157 7147 24191
rect 11161 24157 11195 24191
rect 11805 24157 11839 24191
rect 11897 24157 11931 24191
rect 12541 24157 12575 24191
rect 6193 24089 6227 24123
rect 7665 24089 7699 24123
rect 12771 24089 12805 24123
rect 3157 24021 3191 24055
rect 3709 24021 3743 24055
rect 5273 24021 5307 24055
rect 5641 24021 5675 24055
rect 6837 24021 6871 24055
rect 8769 24021 8803 24055
rect 9045 24021 9079 24055
rect 9873 24021 9907 24055
rect 11897 24021 11931 24055
rect 12081 24021 12115 24055
rect 2789 23817 2823 23851
rect 8493 23817 8527 23851
rect 11253 23817 11287 23851
rect 2513 23749 2547 23783
rect 6653 23749 6687 23783
rect 12633 23749 12667 23783
rect 4353 23681 4387 23715
rect 6837 23681 6871 23715
rect 8677 23681 8711 23715
rect 8953 23681 8987 23715
rect 10885 23681 10919 23715
rect 2605 23613 2639 23647
rect 3525 23613 3559 23647
rect 3617 23613 3651 23647
rect 4169 23613 4203 23647
rect 5181 23613 5215 23647
rect 5733 23613 5767 23647
rect 10057 23613 10091 23647
rect 10425 23613 10459 23647
rect 10609 23613 10643 23647
rect 11529 23613 11563 23647
rect 4997 23545 5031 23579
rect 5917 23545 5951 23579
rect 6285 23545 6319 23579
rect 7158 23545 7192 23579
rect 8769 23545 8803 23579
rect 3157 23477 3191 23511
rect 4721 23477 4755 23511
rect 7757 23477 7791 23511
rect 8033 23477 8067 23511
rect 9689 23477 9723 23511
rect 4353 23273 4387 23307
rect 6193 23273 6227 23307
rect 7297 23273 7331 23307
rect 7941 23273 7975 23307
rect 9873 23273 9907 23307
rect 4997 23205 5031 23239
rect 6739 23205 6773 23239
rect 11253 23205 11287 23239
rect 11805 23205 11839 23239
rect 2973 23137 3007 23171
rect 6377 23137 6411 23171
rect 8125 23137 8159 23171
rect 9689 23137 9723 23171
rect 10149 23137 10183 23171
rect 4905 23069 4939 23103
rect 5549 23069 5583 23103
rect 11161 23069 11195 23103
rect 12633 23069 12667 23103
rect 3157 22933 3191 22967
rect 3709 22933 3743 22967
rect 4721 22933 4755 22967
rect 7573 22933 7607 22967
rect 8309 22933 8343 22967
rect 8585 22933 8619 22967
rect 9045 22933 9079 22967
rect 2973 22729 3007 22763
rect 3525 22729 3559 22763
rect 4077 22729 4111 22763
rect 5825 22729 5859 22763
rect 6469 22729 6503 22763
rect 6561 22729 6595 22763
rect 11437 22729 11471 22763
rect 12633 22729 12667 22763
rect 3801 22661 3835 22695
rect 5549 22661 5583 22695
rect 3617 22525 3651 22559
rect 4629 22525 4663 22559
rect 13645 22661 13679 22695
rect 6929 22593 6963 22627
rect 7205 22593 7239 22627
rect 8217 22593 8251 22627
rect 10425 22593 10459 22627
rect 8401 22525 8435 22559
rect 8953 22525 8987 22559
rect 9965 22525 9999 22559
rect 10057 22525 10091 22559
rect 10241 22525 10275 22559
rect 10977 22525 11011 22559
rect 12449 22525 12483 22559
rect 12909 22525 12943 22559
rect 13461 22525 13495 22559
rect 13921 22525 13955 22559
rect 4537 22457 4571 22491
rect 4991 22457 5025 22491
rect 6561 22457 6595 22491
rect 7021 22457 7055 22491
rect 9137 22457 9171 22491
rect 9505 22389 9539 22423
rect 9781 22389 9815 22423
rect 11713 22389 11747 22423
rect 4353 22185 4387 22219
rect 5457 22185 5491 22219
rect 7665 22185 7699 22219
rect 9413 22185 9447 22219
rect 10425 22185 10459 22219
rect 10977 22185 11011 22219
rect 4899 22117 4933 22151
rect 12541 22117 12575 22151
rect 6285 22049 6319 22083
rect 6745 22049 6779 22083
rect 8677 22049 8711 22083
rect 10057 22049 10091 22083
rect 11805 22049 11839 22083
rect 12081 22049 12115 22083
rect 4537 21981 4571 22015
rect 6837 21981 6871 22015
rect 7389 21981 7423 22015
rect 8769 21981 8803 22015
rect 11897 21913 11931 21947
rect 9873 21845 9907 21879
rect 5273 21641 5307 21675
rect 5917 21641 5951 21675
rect 7941 21641 7975 21675
rect 10977 21641 11011 21675
rect 12633 21641 12667 21675
rect 6929 21573 6963 21607
rect 8493 21573 8527 21607
rect 10057 21573 10091 21607
rect 11345 21573 11379 21607
rect 4813 21505 4847 21539
rect 6285 21505 6319 21539
rect 7573 21505 7607 21539
rect 4169 21437 4203 21471
rect 4721 21437 4755 21471
rect 6837 21437 6871 21471
rect 7113 21437 7147 21471
rect 8401 21437 8435 21471
rect 8677 21437 8711 21471
rect 9965 21437 9999 21471
rect 10241 21437 10275 21471
rect 10701 21437 10735 21471
rect 12449 21437 12483 21471
rect 12909 21437 12943 21471
rect 4077 21369 4111 21403
rect 6653 21369 6687 21403
rect 9137 21369 9171 21403
rect 3801 21301 3835 21335
rect 8309 21301 8343 21335
rect 9505 21301 9539 21335
rect 9873 21301 9907 21335
rect 11805 21301 11839 21335
rect 12173 21301 12207 21335
rect 4261 21097 4295 21131
rect 6285 21097 6319 21131
rect 10149 21097 10183 21131
rect 10793 21097 10827 21131
rect 12265 21097 12299 21131
rect 6745 21029 6779 21063
rect 7297 21029 7331 21063
rect 4261 20961 4295 20995
rect 4629 20961 4663 20995
rect 8160 20961 8194 20995
rect 9781 20961 9815 20995
rect 11253 20961 11287 20995
rect 11529 20961 11563 20995
rect 6653 20893 6687 20927
rect 8263 20893 8297 20927
rect 11713 20893 11747 20927
rect 8677 20825 8711 20859
rect 11345 20825 11379 20859
rect 7573 20757 7607 20791
rect 9505 20757 9539 20791
rect 3617 20553 3651 20587
rect 4629 20553 4663 20587
rect 6285 20553 6319 20587
rect 9781 20553 9815 20587
rect 11989 20553 12023 20587
rect 7481 20485 7515 20519
rect 10057 20485 10091 20519
rect 3847 20417 3881 20451
rect 5457 20417 5491 20451
rect 7849 20417 7883 20451
rect 9137 20417 9171 20451
rect 3760 20349 3794 20383
rect 8309 20349 8343 20383
rect 8769 20349 8803 20383
rect 9965 20349 9999 20383
rect 10241 20349 10275 20383
rect 4813 20281 4847 20315
rect 4905 20281 4939 20315
rect 6929 20281 6963 20315
rect 7021 20281 7055 20315
rect 10701 20281 10735 20315
rect 11345 20281 11379 20315
rect 4261 20213 4295 20247
rect 6653 20213 6687 20247
rect 11713 20213 11747 20247
rect 4813 20009 4847 20043
rect 5089 20009 5123 20043
rect 6469 20009 6503 20043
rect 9505 20009 9539 20043
rect 11621 20009 11655 20043
rect 2973 19941 3007 19975
rect 5870 19941 5904 19975
rect 7481 19941 7515 19975
rect 10609 19941 10643 19975
rect 4307 19873 4341 19907
rect 9873 19873 9907 19907
rect 10149 19873 10183 19907
rect 11437 19873 11471 19907
rect 4399 19805 4433 19839
rect 5549 19805 5583 19839
rect 7389 19805 7423 19839
rect 7941 19737 7975 19771
rect 9965 19737 9999 19771
rect 6929 19669 6963 19703
rect 8309 19669 8343 19703
rect 3801 19465 3835 19499
rect 5181 19465 5215 19499
rect 7849 19465 7883 19499
rect 9689 19465 9723 19499
rect 10609 19465 10643 19499
rect 10885 19465 10919 19499
rect 11529 19465 11563 19499
rect 9321 19397 9355 19431
rect 4077 19329 4111 19363
rect 7573 19329 7607 19363
rect 8953 19329 8987 19363
rect 2697 19261 2731 19295
rect 3249 19261 3283 19295
rect 4261 19261 4295 19295
rect 5917 19261 5951 19295
rect 8585 19261 8619 19295
rect 10425 19261 10459 19295
rect 10609 19261 10643 19295
rect 3433 19193 3467 19227
rect 6929 19193 6963 19227
rect 7021 19193 7055 19227
rect 8309 19193 8343 19227
rect 8401 19193 8435 19227
rect 10517 19193 10551 19227
rect 11161 19193 11195 19227
rect 2513 19125 2547 19159
rect 4629 19125 4663 19159
rect 5549 19125 5583 19159
rect 6653 19125 6687 19159
rect 3249 18921 3283 18955
rect 4261 18921 4295 18955
rect 5457 18921 5491 18955
rect 6469 18921 6503 18955
rect 8309 18921 8343 18955
rect 9413 18921 9447 18955
rect 10701 18921 10735 18955
rect 2789 18853 2823 18887
rect 5911 18853 5945 18887
rect 7481 18853 7515 18887
rect 1961 18785 1995 18819
rect 2881 18785 2915 18819
rect 4604 18785 4638 18819
rect 9045 18785 9079 18819
rect 9677 18785 9711 18819
rect 9965 18785 9999 18819
rect 11897 18785 11931 18819
rect 3525 18717 3559 18751
rect 5549 18717 5583 18751
rect 7389 18717 7423 18751
rect 9781 18717 9815 18751
rect 10425 18717 10459 18751
rect 11253 18717 11287 18751
rect 4675 18649 4709 18683
rect 7941 18649 7975 18683
rect 2099 18581 2133 18615
rect 4997 18581 5031 18615
rect 6837 18581 6871 18615
rect 2053 18377 2087 18411
rect 4629 18377 4663 18411
rect 6009 18377 6043 18411
rect 6561 18377 6595 18411
rect 8033 18377 8067 18411
rect 8493 18377 8527 18411
rect 9597 18377 9631 18411
rect 10333 18377 10367 18411
rect 11437 18377 11471 18411
rect 2605 18309 2639 18343
rect 2973 18309 3007 18343
rect 7757 18309 7791 18343
rect 8861 18309 8895 18343
rect 4169 18241 4203 18275
rect 9468 18241 9502 18275
rect 9689 18241 9723 18275
rect 2421 18173 2455 18207
rect 3433 18173 3467 18207
rect 3893 18173 3927 18207
rect 4997 18173 5031 18207
rect 5549 18173 5583 18207
rect 6837 18173 6871 18207
rect 10057 18173 10091 18207
rect 10885 18173 10919 18207
rect 11713 18173 11747 18207
rect 12449 18173 12483 18207
rect 12909 18173 12943 18207
rect 5733 18105 5767 18139
rect 7158 18105 7192 18139
rect 9321 18105 9355 18139
rect 9229 18037 9263 18071
rect 10793 18037 10827 18071
rect 11069 18037 11103 18071
rect 12633 18037 12667 18071
rect 3157 17833 3191 17867
rect 3525 17833 3559 17867
rect 4215 17833 4249 17867
rect 6101 17833 6135 17867
rect 6561 17833 6595 17867
rect 9321 17833 9355 17867
rect 13277 17833 13311 17867
rect 5825 17765 5859 17799
rect 6745 17765 6779 17799
rect 6837 17765 6871 17799
rect 7389 17765 7423 17799
rect 8125 17765 8159 17799
rect 8217 17765 8251 17799
rect 10793 17765 10827 17799
rect 2973 17697 3007 17731
rect 4144 17697 4178 17731
rect 5273 17697 5307 17731
rect 5549 17697 5583 17731
rect 8401 17697 8435 17731
rect 9677 17697 9711 17731
rect 9781 17697 9815 17731
rect 9965 17697 9999 17731
rect 11529 17697 11563 17731
rect 12817 17697 12851 17731
rect 13093 17697 13127 17731
rect 4997 17629 5031 17663
rect 10149 17629 10183 17663
rect 11253 17629 11287 17663
rect 2513 17561 2547 17595
rect 7757 17561 7791 17595
rect 12909 17561 12943 17595
rect 4629 17493 4663 17527
rect 8493 17493 8527 17527
rect 5273 17289 5307 17323
rect 5641 17289 5675 17323
rect 8309 17289 8343 17323
rect 10057 17289 10091 17323
rect 10425 17289 10459 17323
rect 11621 17289 11655 17323
rect 13553 17289 13587 17323
rect 6285 17221 6319 17255
rect 10701 17221 10735 17255
rect 13185 17221 13219 17255
rect 3065 17153 3099 17187
rect 7573 17153 7607 17187
rect 3801 17085 3835 17119
rect 4261 17085 4295 17119
rect 4721 17085 4755 17119
rect 7113 17085 7147 17119
rect 7205 17085 7239 17119
rect 7389 17085 7423 17119
rect 8953 17085 8987 17119
rect 9321 17085 9355 17119
rect 9505 17085 9539 17119
rect 10609 17085 10643 17119
rect 10885 17085 10919 17119
rect 4997 17017 5031 17051
rect 6653 17017 6687 17051
rect 12909 17017 12943 17051
rect 4169 16949 4203 16983
rect 9781 16949 9815 16983
rect 11069 16949 11103 16983
rect 5273 16745 5307 16779
rect 5917 16745 5951 16779
rect 8033 16745 8067 16779
rect 8769 16745 8803 16779
rect 9137 16745 9171 16779
rect 9505 16745 9539 16779
rect 10793 16745 10827 16779
rect 13691 16745 13725 16779
rect 11989 16677 12023 16711
rect 4261 16609 4295 16643
rect 4721 16609 4755 16643
rect 6653 16609 6687 16643
rect 7573 16609 7607 16643
rect 7665 16609 7699 16643
rect 7849 16609 7883 16643
rect 9689 16609 9723 16643
rect 9965 16609 9999 16643
rect 11897 16609 11931 16643
rect 13553 16609 13587 16643
rect 4813 16541 4847 16575
rect 6745 16541 6779 16575
rect 10149 16541 10183 16575
rect 11069 16541 11103 16575
rect 7205 16473 7239 16507
rect 9781 16473 9815 16507
rect 3755 16201 3789 16235
rect 4537 16201 4571 16235
rect 6101 16201 6135 16235
rect 7849 16201 7883 16235
rect 10057 16201 10091 16235
rect 6561 16133 6595 16167
rect 4629 16065 4663 16099
rect 8585 16065 8619 16099
rect 10885 16065 10919 16099
rect 12449 16065 12483 16099
rect 3525 15997 3559 16031
rect 3652 15997 3686 16031
rect 6837 15997 6871 16031
rect 7389 15997 7423 16031
rect 8861 15997 8895 16031
rect 9321 15997 9355 16031
rect 9505 15997 9539 16031
rect 4950 15929 4984 15963
rect 10977 15929 11011 15963
rect 11529 15929 11563 15963
rect 13553 15929 13587 15963
rect 4169 15861 4203 15895
rect 5549 15861 5583 15895
rect 7113 15861 7147 15895
rect 9597 15861 9631 15895
rect 10701 15861 10735 15895
rect 11897 15861 11931 15895
rect 7757 15657 7791 15691
rect 9045 15657 9079 15691
rect 9505 15657 9539 15691
rect 11161 15657 11195 15691
rect 4950 15589 4984 15623
rect 6561 15589 6595 15623
rect 7113 15589 7147 15623
rect 10194 15589 10228 15623
rect 11805 15589 11839 15623
rect 4629 15521 4663 15555
rect 7941 15521 7975 15555
rect 8217 15521 8251 15555
rect 9873 15521 9907 15555
rect 10793 15521 10827 15555
rect 2973 15453 3007 15487
rect 6469 15453 6503 15487
rect 8033 15453 8067 15487
rect 8401 15453 8435 15487
rect 11713 15453 11747 15487
rect 11989 15453 12023 15487
rect 4261 15317 4295 15351
rect 5549 15317 5583 15351
rect 6193 15317 6227 15351
rect 7481 15317 7515 15351
rect 5549 15113 5583 15147
rect 6561 15113 6595 15147
rect 7849 15113 7883 15147
rect 9413 15113 9447 15147
rect 10333 15113 10367 15147
rect 11069 15113 11103 15147
rect 11805 15113 11839 15147
rect 3893 15045 3927 15079
rect 5181 15045 5215 15079
rect 5917 15045 5951 15079
rect 6285 15045 6319 15079
rect 2329 14977 2363 15011
rect 7205 14977 7239 15011
rect 2697 14909 2731 14943
rect 2973 14909 3007 14943
rect 3985 14909 4019 14943
rect 5733 14909 5767 14943
rect 8401 14909 8435 14943
rect 8861 14909 8895 14943
rect 10701 14909 10735 14943
rect 11437 14909 11471 14943
rect 3157 14841 3191 14875
rect 3433 14841 3467 14875
rect 4347 14841 4381 14875
rect 6929 14841 6963 14875
rect 7021 14841 7055 14875
rect 4905 14773 4939 14807
rect 8217 14773 8251 14807
rect 8493 14773 8527 14807
rect 9873 14773 9907 14807
rect 12173 14773 12207 14807
rect 2513 14569 2547 14603
rect 6193 14569 6227 14603
rect 7205 14569 7239 14603
rect 8861 14569 8895 14603
rect 9505 14569 9539 14603
rect 4721 14501 4755 14535
rect 6745 14501 6779 14535
rect 7618 14501 7652 14535
rect 10010 14501 10044 14535
rect 6285 14433 6319 14467
rect 7297 14433 7331 14467
rect 9689 14433 9723 14467
rect 11472 14433 11506 14467
rect 4629 14365 4663 14399
rect 5089 14365 5123 14399
rect 6469 14297 6503 14331
rect 5549 14229 5583 14263
rect 8217 14229 8251 14263
rect 8585 14229 8619 14263
rect 10609 14229 10643 14263
rect 11575 14229 11609 14263
rect 4629 14025 4663 14059
rect 6377 14025 6411 14059
rect 7113 14025 7147 14059
rect 9045 14025 9079 14059
rect 9781 14025 9815 14059
rect 10977 14025 11011 14059
rect 3525 13889 3559 13923
rect 7297 13889 7331 13923
rect 8493 13889 8527 13923
rect 9965 13889 9999 13923
rect 3617 13821 3651 13855
rect 4169 13821 4203 13855
rect 4353 13821 4387 13855
rect 5273 13753 5307 13787
rect 5365 13753 5399 13787
rect 5917 13753 5951 13787
rect 7618 13753 7652 13787
rect 9413 13753 9447 13787
rect 10057 13753 10091 13787
rect 10609 13753 10643 13787
rect 5089 13685 5123 13719
rect 8217 13685 8251 13719
rect 11437 13685 11471 13719
rect 3617 13481 3651 13515
rect 4629 13481 4663 13515
rect 7297 13481 7331 13515
rect 7757 13481 7791 13515
rect 3111 13413 3145 13447
rect 5451 13413 5485 13447
rect 8217 13413 8251 13447
rect 10057 13413 10091 13447
rect 10609 13413 10643 13447
rect 3024 13345 3058 13379
rect 4144 13345 4178 13379
rect 11437 13345 11471 13379
rect 5089 13277 5123 13311
rect 6837 13277 6871 13311
rect 8125 13277 8159 13311
rect 9965 13277 9999 13311
rect 11575 13277 11609 13311
rect 8677 13209 8711 13243
rect 4215 13141 4249 13175
rect 4905 13141 4939 13175
rect 6009 13141 6043 13175
rect 9045 13141 9079 13175
rect 6193 12937 6227 12971
rect 6653 12937 6687 12971
rect 8125 12937 8159 12971
rect 8401 12937 8435 12971
rect 11437 12937 11471 12971
rect 4721 12869 4755 12903
rect 4353 12801 4387 12835
rect 5641 12801 5675 12835
rect 6837 12801 6871 12835
rect 8953 12801 8987 12835
rect 9965 12801 9999 12835
rect 10149 12801 10183 12835
rect 3893 12733 3927 12767
rect 4169 12733 4203 12767
rect 4997 12733 5031 12767
rect 10701 12733 10735 12767
rect 3525 12665 3559 12699
rect 5273 12665 5307 12699
rect 5365 12665 5399 12699
rect 8677 12665 8711 12699
rect 8769 12665 8803 12699
rect 3065 12597 3099 12631
rect 7205 12597 7239 12631
rect 7757 12597 7791 12631
rect 3709 12393 3743 12427
rect 4721 12393 4755 12427
rect 6009 12393 6043 12427
rect 7665 12393 7699 12427
rect 9781 12393 9815 12427
rect 10701 12393 10735 12427
rect 3111 12325 3145 12359
rect 5089 12325 5123 12359
rect 6653 12325 6687 12359
rect 8217 12325 8251 12359
rect 9045 12325 9079 12359
rect 9505 12325 9539 12359
rect 3024 12257 3058 12291
rect 9965 12257 9999 12291
rect 10149 12257 10183 12291
rect 11320 12257 11354 12291
rect 4997 12189 5031 12223
rect 5641 12189 5675 12223
rect 6561 12189 6595 12223
rect 8125 12189 8159 12223
rect 7113 12121 7147 12155
rect 8677 12121 8711 12155
rect 11391 12121 11425 12155
rect 2973 11849 3007 11883
rect 4629 11849 4663 11883
rect 4997 11849 5031 11883
rect 6561 11849 6595 11883
rect 7021 11849 7055 11883
rect 7481 11849 7515 11883
rect 8585 11849 8619 11883
rect 8861 11849 8895 11883
rect 10057 11781 10091 11815
rect 6101 11713 6135 11747
rect 7665 11713 7699 11747
rect 9505 11713 9539 11747
rect 10793 11713 10827 11747
rect 11115 11713 11149 11747
rect 3433 11645 3467 11679
rect 3525 11645 3559 11679
rect 4077 11645 4111 11679
rect 11028 11645 11062 11679
rect 11805 11645 11839 11679
rect 4261 11577 4295 11611
rect 5181 11577 5215 11611
rect 5273 11577 5307 11611
rect 5825 11577 5859 11611
rect 7986 11577 8020 11611
rect 9597 11577 9631 11611
rect 10425 11577 10459 11611
rect 9229 11509 9263 11543
rect 11437 11509 11471 11543
rect 3617 11305 3651 11339
rect 4629 11305 4663 11339
rect 5181 11305 5215 11339
rect 8585 11305 8619 11339
rect 9505 11305 9539 11339
rect 7618 11237 7652 11271
rect 9873 11237 9907 11271
rect 10425 11237 10459 11271
rect 11437 11237 11471 11271
rect 2421 11169 2455 11203
rect 2973 11169 3007 11203
rect 6352 11169 6386 11203
rect 3157 11101 3191 11135
rect 4261 11101 4295 11135
rect 7297 11101 7331 11135
rect 9781 11101 9815 11135
rect 11345 11101 11379 11135
rect 11897 11033 11931 11067
rect 5457 10965 5491 10999
rect 6423 10965 6457 10999
rect 8217 10965 8251 10999
rect 2421 10761 2455 10795
rect 2881 10761 2915 10795
rect 3571 10761 3605 10795
rect 5641 10761 5675 10795
rect 6377 10761 6411 10795
rect 7297 10761 7331 10795
rect 10241 10761 10275 10795
rect 10609 10761 10643 10795
rect 10931 10761 10965 10795
rect 11621 10761 11655 10795
rect 8401 10693 8435 10727
rect 9137 10693 9171 10727
rect 8677 10625 8711 10659
rect 9965 10625 9999 10659
rect 3500 10557 3534 10591
rect 4445 10557 4479 10591
rect 7481 10557 7515 10591
rect 10860 10557 10894 10591
rect 11253 10557 11287 10591
rect 4353 10489 4387 10523
rect 4766 10489 4800 10523
rect 7802 10489 7836 10523
rect 9321 10489 9355 10523
rect 9413 10489 9447 10523
rect 3985 10421 4019 10455
rect 5365 10421 5399 10455
rect 11989 10421 12023 10455
rect 3111 10217 3145 10251
rect 5089 10217 5123 10251
rect 7481 10217 7515 10251
rect 9321 10217 9355 10251
rect 9827 10217 9861 10251
rect 5457 10149 5491 10183
rect 8217 10149 8251 10183
rect 8769 10149 8803 10183
rect 4312 10081 4346 10115
rect 9597 10081 9631 10115
rect 4399 10013 4433 10047
rect 5365 10013 5399 10047
rect 5641 10013 5675 10047
rect 6837 10013 6871 10047
rect 8125 10013 8159 10047
rect 2881 9877 2915 9911
rect 4721 9877 4755 9911
rect 7849 9877 7883 9911
rect 3985 9673 4019 9707
rect 4721 9673 4755 9707
rect 8125 9673 8159 9707
rect 8539 9673 8573 9707
rect 5825 9605 5859 9639
rect 9229 9605 9263 9639
rect 7573 9537 7607 9571
rect 4220 9469 4254 9503
rect 6837 9469 6871 9503
rect 7297 9469 7331 9503
rect 8468 9469 8502 9503
rect 3709 9401 3743 9435
rect 4307 9401 4341 9435
rect 5273 9401 5307 9435
rect 5365 9401 5399 9435
rect 6561 9401 6595 9435
rect 2973 9333 3007 9367
rect 5089 9333 5123 9367
rect 6285 9333 6319 9367
rect 8861 9333 8895 9367
rect 9689 9333 9723 9367
rect 5641 9129 5675 9163
rect 6009 9129 6043 9163
rect 8953 9129 8987 9163
rect 7297 9061 7331 9095
rect 4445 8993 4479 9027
rect 4721 8993 4755 9027
rect 6561 8993 6595 9027
rect 7113 8993 7147 9027
rect 8125 8993 8159 9027
rect 4813 8925 4847 8959
rect 6469 8925 6503 8959
rect 8309 8857 8343 8891
rect 8585 8857 8619 8891
rect 5365 8789 5399 8823
rect 7665 8789 7699 8823
rect 4997 8585 5031 8619
rect 6193 8585 6227 8619
rect 8217 8585 8251 8619
rect 3525 8449 3559 8483
rect 6837 8449 6871 8483
rect 3893 8381 3927 8415
rect 4169 8381 4203 8415
rect 5181 8381 5215 8415
rect 5641 8381 5675 8415
rect 6653 8381 6687 8415
rect 8585 8381 8619 8415
rect 9045 8381 9079 8415
rect 4353 8313 4387 8347
rect 5917 8313 5951 8347
rect 7158 8313 7192 8347
rect 4721 8245 4755 8279
rect 7757 8245 7791 8279
rect 8677 8245 8711 8279
rect 3249 8041 3283 8075
rect 3709 8041 3743 8075
rect 4261 8041 4295 8075
rect 4813 8041 4847 8075
rect 7757 8041 7791 8075
rect 9781 8041 9815 8075
rect 6653 7973 6687 8007
rect 8217 7973 8251 8007
rect 5181 7905 5215 7939
rect 5365 7905 5399 7939
rect 9965 7905 9999 7939
rect 10149 7905 10183 7939
rect 5641 7837 5675 7871
rect 6561 7837 6595 7871
rect 8125 7837 8159 7871
rect 8769 7837 8803 7871
rect 7113 7769 7147 7803
rect 9505 7701 9539 7735
rect 7021 7497 7055 7531
rect 8585 7497 8619 7531
rect 8861 7497 8895 7531
rect 10425 7497 10459 7531
rect 6561 7429 6595 7463
rect 9229 7429 9263 7463
rect 11437 7429 11471 7463
rect 3065 7361 3099 7395
rect 4721 7361 4755 7395
rect 7665 7361 7699 7395
rect 9505 7361 9539 7395
rect 11115 7361 11149 7395
rect 3433 7293 3467 7327
rect 3709 7293 3743 7327
rect 4629 7293 4663 7327
rect 11028 7293 11062 7327
rect 3893 7225 3927 7259
rect 5083 7225 5117 7259
rect 7986 7225 8020 7259
rect 9597 7225 9631 7259
rect 10149 7225 10183 7259
rect 4261 7157 4295 7191
rect 5641 7157 5675 7191
rect 7481 7157 7515 7191
rect 6469 6953 6503 6987
rect 9505 6953 9539 6987
rect 4997 6885 5031 6919
rect 5594 6885 5628 6919
rect 7802 6885 7836 6919
rect 9873 6885 9907 6919
rect 2421 6817 2455 6851
rect 2973 6817 3007 6851
rect 4261 6817 4295 6851
rect 5273 6817 5307 6851
rect 7481 6817 7515 6851
rect 3157 6749 3191 6783
rect 9781 6749 9815 6783
rect 10057 6749 10091 6783
rect 4445 6681 4479 6715
rect 6193 6613 6227 6647
rect 8401 6613 8435 6647
rect 8769 6613 8803 6647
rect 2329 6409 2363 6443
rect 2881 6409 2915 6443
rect 3249 6409 3283 6443
rect 4537 6409 4571 6443
rect 6193 6409 6227 6443
rect 9045 6409 9079 6443
rect 9873 6341 9907 6375
rect 2559 6273 2593 6307
rect 4997 6273 5031 6307
rect 7481 6273 7515 6307
rect 8677 6273 8711 6307
rect 10241 6273 10275 6307
rect 2472 6205 2506 6239
rect 3433 6205 3467 6239
rect 3985 6205 4019 6239
rect 8401 6205 8435 6239
rect 4169 6137 4203 6171
rect 5318 6137 5352 6171
rect 6561 6137 6595 6171
rect 7297 6137 7331 6171
rect 7802 6137 7836 6171
rect 9321 6137 9355 6171
rect 9413 6137 9447 6171
rect 4905 6069 4939 6103
rect 5917 6069 5951 6103
rect 10609 6069 10643 6103
rect 2421 5865 2455 5899
rect 3525 5865 3559 5899
rect 7297 5865 7331 5899
rect 8217 5865 8251 5899
rect 9321 5865 9355 5899
rect 9827 5865 9861 5899
rect 5825 5797 5859 5831
rect 4077 5729 4111 5763
rect 4537 5729 4571 5763
rect 7205 5729 7239 5763
rect 7665 5729 7699 5763
rect 9724 5729 9758 5763
rect 4813 5661 4847 5695
rect 5733 5661 5767 5695
rect 6009 5661 6043 5695
rect 5273 5525 5307 5559
rect 4629 5321 4663 5355
rect 5089 5321 5123 5355
rect 6193 5321 6227 5355
rect 7757 5321 7791 5355
rect 9689 5321 9723 5355
rect 6561 5253 6595 5287
rect 10011 5253 10045 5287
rect 5273 5185 5307 5219
rect 5733 5185 5767 5219
rect 9045 5185 9079 5219
rect 3525 5117 3559 5151
rect 3893 5117 3927 5151
rect 4077 5117 4111 5151
rect 6837 5117 6871 5151
rect 7389 5117 7423 5151
rect 9940 5117 9974 5151
rect 10333 5117 10367 5151
rect 4353 5049 4387 5083
rect 5374 5049 5408 5083
rect 8401 5049 8435 5083
rect 8493 5049 8527 5083
rect 7021 4981 7055 5015
rect 8217 4981 8251 5015
rect 3709 4777 3743 4811
rect 4353 4777 4387 4811
rect 6285 4777 6319 4811
rect 8217 4777 8251 4811
rect 5042 4709 5076 4743
rect 7113 4709 7147 4743
rect 7618 4709 7652 4743
rect 8585 4709 8619 4743
rect 9827 4709 9861 4743
rect 3040 4641 3074 4675
rect 5917 4641 5951 4675
rect 7297 4641 7331 4675
rect 9740 4641 9774 4675
rect 10736 4641 10770 4675
rect 4721 4573 4755 4607
rect 5641 4505 5675 4539
rect 3111 4437 3145 4471
rect 8953 4437 8987 4471
rect 10839 4437 10873 4471
rect 6193 4233 6227 4267
rect 6653 4233 6687 4267
rect 8677 4233 8711 4267
rect 9965 4233 9999 4267
rect 10333 4233 10367 4267
rect 10977 4233 11011 4267
rect 2145 4165 2179 4199
rect 4261 4165 4295 4199
rect 2743 4097 2777 4131
rect 5273 4097 5307 4131
rect 7113 4097 7147 4131
rect 8953 4097 8987 4131
rect 9229 4097 9263 4131
rect 1660 4029 1694 4063
rect 2656 4029 2690 4063
rect 3065 4029 3099 4063
rect 4813 4029 4847 4063
rect 10425 4029 10459 4063
rect 2513 3961 2547 3995
rect 3709 3961 3743 3995
rect 3801 3961 3835 3995
rect 5365 3961 5399 3995
rect 5917 3961 5951 3995
rect 7475 3961 7509 3995
rect 9045 3961 9079 3995
rect 1731 3893 1765 3927
rect 3525 3893 3559 3927
rect 8033 3893 8067 3927
rect 10609 3893 10643 3927
rect 3709 3689 3743 3723
rect 5365 3689 5399 3723
rect 5641 3689 5675 3723
rect 7205 3689 7239 3723
rect 7573 3689 7607 3723
rect 7941 3689 7975 3723
rect 10931 3689 10965 3723
rect 1869 3621 1903 3655
rect 4439 3621 4473 3655
rect 6009 3621 6043 3655
rect 6561 3621 6595 3655
rect 8217 3621 8251 3655
rect 8769 3621 8803 3655
rect 2028 3553 2062 3587
rect 4077 3553 4111 3587
rect 9689 3553 9723 3587
rect 10828 3553 10862 3587
rect 2973 3485 3007 3519
rect 5917 3485 5951 3519
rect 8125 3485 8159 3519
rect 2099 3417 2133 3451
rect 2697 3349 2731 3383
rect 4997 3349 5031 3383
rect 9873 3349 9907 3383
rect 1501 3145 1535 3179
rect 2145 3145 2179 3179
rect 2513 3145 2547 3179
rect 5365 3145 5399 3179
rect 5917 3145 5951 3179
rect 6193 3145 6227 3179
rect 8033 3145 8067 3179
rect 9229 3145 9263 3179
rect 9597 3145 9631 3179
rect 10241 3145 10275 3179
rect 11621 3145 11655 3179
rect 1731 3077 1765 3111
rect 8769 3077 8803 3111
rect 2697 3009 2731 3043
rect 4169 3009 4203 3043
rect 8217 3009 8251 3043
rect 3341 2941 3375 2975
rect 6837 2941 6871 2975
rect 7389 2941 7423 2975
rect 9689 2941 9723 2975
rect 10828 2941 10862 2975
rect 11253 2941 11287 2975
rect 2789 2873 2823 2907
rect 4531 2873 4565 2907
rect 8309 2873 8343 2907
rect 3709 2805 3743 2839
rect 3985 2805 4019 2839
rect 5089 2805 5123 2839
rect 7021 2805 7055 2839
rect 9873 2805 9907 2839
rect 10931 2805 10965 2839
rect 3525 2601 3559 2635
rect 4261 2601 4295 2635
rect 6653 2601 6687 2635
rect 8125 2601 8159 2635
rect 11621 2601 11655 2635
rect 2329 2533 2363 2567
rect 2513 2533 2547 2567
rect 2605 2533 2639 2567
rect 3157 2533 3191 2567
rect 4813 2533 4847 2567
rect 5089 2533 5123 2567
rect 5641 2533 5675 2567
rect 7113 2533 7147 2567
rect 10885 2533 10919 2567
rect 1476 2465 1510 2499
rect 8493 2465 8527 2499
rect 9045 2465 9079 2499
rect 10333 2465 10367 2499
rect 11437 2465 11471 2499
rect 11989 2465 12023 2499
rect 13185 2465 13219 2499
rect 13737 2465 13771 2499
rect 4997 2397 5031 2431
rect 5917 2397 5951 2431
rect 6377 2397 6411 2431
rect 7021 2397 7055 2431
rect 1961 2329 1995 2363
rect 7573 2329 7607 2363
rect 10517 2329 10551 2363
rect 13369 2329 13403 2363
rect 1547 2261 1581 2295
rect 8677 2261 8711 2295
<< metal1 >>
rect 1210 39652 1216 39704
rect 1268 39692 1274 39704
rect 3234 39692 3240 39704
rect 1268 39664 3240 39692
rect 1268 39652 1274 39664
rect 3234 39652 3240 39664
rect 3292 39652 3298 39704
rect 1394 39584 1400 39636
rect 1452 39624 1458 39636
rect 2130 39624 2136 39636
rect 1452 39596 2136 39624
rect 1452 39584 1458 39596
rect 2130 39584 2136 39596
rect 2188 39584 2194 39636
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 9652 36703 9710 36709
rect 9652 36669 9664 36703
rect 9698 36700 9710 36703
rect 10045 36703 10103 36709
rect 10045 36700 10057 36703
rect 9698 36672 10057 36700
rect 9698 36669 9710 36672
rect 9652 36663 9710 36669
rect 10045 36669 10057 36672
rect 10091 36700 10103 36703
rect 12434 36700 12440 36712
rect 10091 36672 12440 36700
rect 10091 36669 10103 36672
rect 10045 36663 10103 36669
rect 12434 36660 12440 36672
rect 12492 36660 12498 36712
rect 9723 36567 9781 36573
rect 9723 36533 9735 36567
rect 9769 36564 9781 36567
rect 9950 36564 9956 36576
rect 9769 36536 9956 36564
rect 9769 36533 9781 36536
rect 9723 36527 9781 36533
rect 9950 36524 9956 36536
rect 10008 36524 10014 36576
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 8665 36363 8723 36369
rect 8665 36329 8677 36363
rect 8711 36360 8723 36363
rect 8846 36360 8852 36372
rect 8711 36332 8852 36360
rect 8711 36329 8723 36332
rect 8665 36323 8723 36329
rect 8846 36320 8852 36332
rect 8904 36320 8910 36372
rect 2958 36252 2964 36304
rect 3016 36292 3022 36304
rect 3016 36264 9628 36292
rect 3016 36252 3022 36264
rect 7558 36233 7564 36236
rect 7536 36227 7564 36233
rect 7536 36224 7548 36227
rect 7471 36196 7548 36224
rect 7536 36193 7548 36196
rect 7616 36224 7622 36236
rect 7834 36224 7840 36236
rect 7616 36196 7840 36224
rect 7536 36187 7564 36193
rect 7558 36184 7564 36187
rect 7616 36184 7622 36196
rect 7834 36184 7840 36196
rect 7892 36184 7898 36236
rect 8386 36184 8392 36236
rect 8444 36224 8450 36236
rect 8481 36227 8539 36233
rect 8481 36224 8493 36227
rect 8444 36196 8493 36224
rect 8444 36184 8450 36196
rect 8481 36193 8493 36196
rect 8527 36193 8539 36227
rect 9600 36224 9628 36264
rect 9674 36224 9680 36236
rect 9732 36233 9738 36236
rect 9732 36227 9770 36233
rect 9587 36196 9680 36224
rect 8481 36187 8539 36193
rect 9674 36184 9680 36196
rect 9758 36193 9770 36227
rect 9732 36187 9770 36193
rect 9732 36184 9738 36187
rect 7607 36023 7665 36029
rect 7607 35989 7619 36023
rect 7653 36020 7665 36023
rect 8110 36020 8116 36032
rect 7653 35992 8116 36020
rect 7653 35989 7665 35992
rect 7607 35983 7665 35989
rect 8110 35980 8116 35992
rect 8168 35980 8174 36032
rect 8202 35980 8208 36032
rect 8260 36020 8266 36032
rect 9815 36023 9873 36029
rect 8260 35992 8305 36020
rect 8260 35980 8266 35992
rect 9815 35989 9827 36023
rect 9861 36020 9873 36023
rect 10229 36023 10287 36029
rect 10229 36020 10241 36023
rect 9861 35992 10241 36020
rect 9861 35989 9873 35992
rect 9815 35983 9873 35989
rect 10229 35989 10241 35992
rect 10275 36020 10287 36023
rect 10318 36020 10324 36032
rect 10275 35992 10324 36020
rect 10275 35989 10287 35992
rect 10229 35983 10287 35989
rect 10318 35980 10324 35992
rect 10376 35980 10382 36032
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 7009 35819 7067 35825
rect 7009 35785 7021 35819
rect 7055 35816 7067 35819
rect 13446 35816 13452 35828
rect 7055 35788 13452 35816
rect 7055 35785 7067 35788
rect 7009 35779 7067 35785
rect 13446 35776 13452 35788
rect 13504 35776 13510 35828
rect 7834 35748 7840 35760
rect 7747 35720 7840 35748
rect 7834 35708 7840 35720
rect 7892 35748 7898 35760
rect 11238 35748 11244 35760
rect 7892 35720 11244 35748
rect 7892 35708 7898 35720
rect 11238 35708 11244 35720
rect 11296 35708 11302 35760
rect 8110 35640 8116 35692
rect 8168 35680 8174 35692
rect 8297 35683 8355 35689
rect 8297 35680 8309 35683
rect 8168 35652 8309 35680
rect 8168 35640 8174 35652
rect 8297 35649 8309 35652
rect 8343 35649 8355 35683
rect 8297 35643 8355 35649
rect 8386 35640 8392 35692
rect 8444 35680 8450 35692
rect 9217 35683 9275 35689
rect 9217 35680 9229 35683
rect 8444 35652 9229 35680
rect 8444 35640 8450 35652
rect 9217 35649 9229 35652
rect 9263 35649 9275 35683
rect 9674 35680 9680 35692
rect 9635 35652 9680 35680
rect 9217 35643 9275 35649
rect 9674 35640 9680 35652
rect 9732 35640 9738 35692
rect 10318 35680 10324 35692
rect 10279 35652 10324 35680
rect 10318 35640 10324 35652
rect 10376 35640 10382 35692
rect 4430 35572 4436 35624
rect 4488 35612 4494 35624
rect 6825 35615 6883 35621
rect 6825 35612 6837 35615
rect 4488 35584 6837 35612
rect 4488 35572 4494 35584
rect 6825 35581 6837 35584
rect 6871 35612 6883 35615
rect 7377 35615 7435 35621
rect 7377 35612 7389 35615
rect 6871 35584 7389 35612
rect 6871 35581 6883 35584
rect 6825 35575 6883 35581
rect 7377 35581 7389 35584
rect 7423 35581 7435 35615
rect 7377 35575 7435 35581
rect 8389 35547 8447 35553
rect 8389 35513 8401 35547
rect 8435 35513 8447 35547
rect 8389 35507 8447 35513
rect 8202 35436 8208 35488
rect 8260 35476 8266 35488
rect 8404 35476 8432 35507
rect 8478 35504 8484 35556
rect 8536 35544 8542 35556
rect 8941 35547 8999 35553
rect 8941 35544 8953 35547
rect 8536 35516 8953 35544
rect 8536 35504 8542 35516
rect 8941 35513 8953 35516
rect 8987 35513 8999 35547
rect 8941 35507 8999 35513
rect 10137 35547 10195 35553
rect 10137 35513 10149 35547
rect 10183 35544 10195 35547
rect 10410 35544 10416 35556
rect 10183 35516 10416 35544
rect 10183 35513 10195 35516
rect 10137 35507 10195 35513
rect 10410 35504 10416 35516
rect 10468 35504 10474 35556
rect 10962 35544 10968 35556
rect 10923 35516 10968 35544
rect 10962 35504 10968 35516
rect 11020 35504 11026 35556
rect 8260 35448 8432 35476
rect 8260 35436 8266 35448
rect 9674 35436 9680 35488
rect 9732 35476 9738 35488
rect 10870 35476 10876 35488
rect 9732 35448 10876 35476
rect 9732 35436 9738 35448
rect 10870 35436 10876 35448
rect 10928 35436 10934 35488
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 7101 35275 7159 35281
rect 7101 35241 7113 35275
rect 7147 35272 7159 35275
rect 8018 35272 8024 35284
rect 7147 35244 8024 35272
rect 7147 35241 7159 35244
rect 7101 35235 7159 35241
rect 8018 35232 8024 35244
rect 8076 35232 8082 35284
rect 8110 35232 8116 35284
rect 8168 35272 8174 35284
rect 9033 35275 9091 35281
rect 9033 35272 9045 35275
rect 8168 35244 9045 35272
rect 8168 35232 8174 35244
rect 9033 35241 9045 35244
rect 9079 35241 9091 35275
rect 9033 35235 9091 35241
rect 9950 35232 9956 35284
rect 10008 35272 10014 35284
rect 10229 35275 10287 35281
rect 10229 35272 10241 35275
rect 10008 35244 10241 35272
rect 10008 35232 10014 35244
rect 10229 35241 10241 35244
rect 10275 35241 10287 35275
rect 10229 35235 10287 35241
rect 13173 35275 13231 35281
rect 13173 35241 13185 35275
rect 13219 35272 13231 35275
rect 14642 35272 14648 35284
rect 13219 35244 14648 35272
rect 13219 35241 13231 35244
rect 13173 35235 13231 35241
rect 14642 35232 14648 35244
rect 14700 35232 14706 35284
rect 5810 35164 5816 35216
rect 5868 35204 5874 35216
rect 6043 35207 6101 35213
rect 6043 35204 6055 35207
rect 5868 35176 6055 35204
rect 5868 35164 5874 35176
rect 6043 35173 6055 35176
rect 6089 35173 6101 35207
rect 8202 35204 8208 35216
rect 8163 35176 8208 35204
rect 6043 35167 6101 35173
rect 8202 35164 8208 35176
rect 8260 35164 8266 35216
rect 10594 35204 10600 35216
rect 10555 35176 10600 35204
rect 10594 35164 10600 35176
rect 10652 35164 10658 35216
rect 5956 35139 6014 35145
rect 5956 35105 5968 35139
rect 6002 35136 6014 35139
rect 6730 35136 6736 35148
rect 6002 35108 6736 35136
rect 6002 35105 6014 35108
rect 5956 35099 6014 35105
rect 6730 35096 6736 35108
rect 6788 35096 6794 35148
rect 6917 35139 6975 35145
rect 6917 35105 6929 35139
rect 6963 35136 6975 35139
rect 7006 35136 7012 35148
rect 6963 35108 7012 35136
rect 6963 35105 6975 35108
rect 6917 35099 6975 35105
rect 7006 35096 7012 35108
rect 7064 35096 7070 35148
rect 12044 35139 12102 35145
rect 12044 35105 12056 35139
rect 12090 35136 12102 35139
rect 12158 35136 12164 35148
rect 12090 35108 12164 35136
rect 12090 35105 12102 35108
rect 12044 35099 12102 35105
rect 12158 35096 12164 35108
rect 12216 35096 12222 35148
rect 12986 35136 12992 35148
rect 12947 35108 12992 35136
rect 12986 35096 12992 35108
rect 13044 35096 13050 35148
rect 8110 35068 8116 35080
rect 8071 35040 8116 35068
rect 8110 35028 8116 35040
rect 8168 35028 8174 35080
rect 8294 35028 8300 35080
rect 8352 35068 8358 35080
rect 8389 35071 8447 35077
rect 8389 35068 8401 35071
rect 8352 35040 8401 35068
rect 8352 35028 8358 35040
rect 8389 35037 8401 35040
rect 8435 35037 8447 35071
rect 10502 35068 10508 35080
rect 10463 35040 10508 35068
rect 8389 35031 8447 35037
rect 10502 35028 10508 35040
rect 10560 35028 10566 35080
rect 11149 35071 11207 35077
rect 11149 35037 11161 35071
rect 11195 35068 11207 35071
rect 11422 35068 11428 35080
rect 11195 35040 11428 35068
rect 11195 35037 11207 35040
rect 11149 35031 11207 35037
rect 11422 35028 11428 35040
rect 11480 35028 11486 35080
rect 5810 34960 5816 35012
rect 5868 35000 5874 35012
rect 12618 35000 12624 35012
rect 5868 34972 12624 35000
rect 5868 34960 5874 34972
rect 12618 34960 12624 34972
rect 12676 34960 12682 35012
rect 7650 34932 7656 34944
rect 7611 34904 7656 34932
rect 7650 34892 7656 34904
rect 7708 34892 7714 34944
rect 12115 34935 12173 34941
rect 12115 34901 12127 34935
rect 12161 34932 12173 34935
rect 12526 34932 12532 34944
rect 12161 34904 12532 34932
rect 12161 34901 12173 34904
rect 12115 34895 12173 34901
rect 12526 34892 12532 34904
rect 12584 34892 12590 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 5810 34728 5816 34740
rect 5771 34700 5816 34728
rect 5810 34688 5816 34700
rect 5868 34688 5874 34740
rect 9309 34731 9367 34737
rect 9309 34697 9321 34731
rect 9355 34728 9367 34731
rect 9766 34728 9772 34740
rect 9355 34700 9772 34728
rect 9355 34697 9367 34700
rect 9309 34691 9367 34697
rect 9766 34688 9772 34700
rect 9824 34688 9830 34740
rect 11330 34688 11336 34740
rect 11388 34728 11394 34740
rect 12621 34731 12679 34737
rect 12621 34728 12633 34731
rect 11388 34700 12633 34728
rect 11388 34688 11394 34700
rect 12621 34697 12633 34700
rect 12667 34697 12679 34731
rect 12621 34691 12679 34697
rect 7742 34620 7748 34672
rect 7800 34660 7806 34672
rect 12069 34663 12127 34669
rect 7800 34632 9168 34660
rect 7800 34620 7806 34632
rect 8294 34592 8300 34604
rect 8255 34564 8300 34592
rect 8294 34552 8300 34564
rect 8352 34552 8358 34604
rect 4154 34484 4160 34536
rect 4212 34524 4218 34536
rect 9140 34533 9168 34632
rect 12069 34629 12081 34663
rect 12115 34660 12127 34663
rect 12158 34660 12164 34672
rect 12115 34632 12164 34660
rect 12115 34629 12127 34632
rect 12069 34623 12127 34629
rect 12158 34620 12164 34632
rect 12216 34620 12222 34672
rect 9950 34552 9956 34604
rect 10008 34592 10014 34604
rect 10321 34595 10379 34601
rect 10321 34592 10333 34595
rect 10008 34564 10333 34592
rect 10008 34552 10014 34564
rect 10321 34561 10333 34564
rect 10367 34561 10379 34595
rect 10962 34592 10968 34604
rect 10923 34564 10968 34592
rect 10321 34555 10379 34561
rect 10962 34552 10968 34564
rect 11020 34552 11026 34604
rect 13081 34595 13139 34601
rect 13081 34592 13093 34595
rect 12452 34564 13093 34592
rect 12452 34536 12480 34564
rect 13081 34561 13093 34564
rect 13127 34561 13139 34595
rect 13081 34555 13139 34561
rect 5629 34527 5687 34533
rect 5629 34524 5641 34527
rect 4212 34496 5641 34524
rect 4212 34484 4218 34496
rect 5629 34493 5641 34496
rect 5675 34524 5687 34527
rect 6181 34527 6239 34533
rect 6181 34524 6193 34527
rect 5675 34496 6193 34524
rect 5675 34493 5687 34496
rect 5629 34487 5687 34493
rect 6181 34493 6193 34496
rect 6227 34493 6239 34527
rect 6181 34487 6239 34493
rect 9125 34527 9183 34533
rect 9125 34493 9137 34527
rect 9171 34524 9183 34527
rect 9677 34527 9735 34533
rect 9677 34524 9689 34527
rect 9171 34496 9689 34524
rect 9171 34493 9183 34496
rect 9125 34487 9183 34493
rect 9677 34493 9689 34496
rect 9723 34493 9735 34527
rect 12434 34524 12440 34536
rect 12395 34496 12440 34524
rect 9677 34487 9735 34493
rect 12434 34484 12440 34496
rect 12492 34484 12498 34536
rect 12986 34484 12992 34536
rect 13044 34524 13050 34536
rect 13357 34527 13415 34533
rect 13357 34524 13369 34527
rect 13044 34496 13369 34524
rect 13044 34484 13050 34496
rect 13357 34493 13369 34496
rect 13403 34493 13415 34527
rect 13357 34487 13415 34493
rect 6086 34416 6092 34468
rect 6144 34456 6150 34468
rect 7650 34456 7656 34468
rect 6144 34428 7656 34456
rect 6144 34416 6150 34428
rect 7650 34416 7656 34428
rect 7708 34416 7714 34468
rect 7745 34459 7803 34465
rect 7745 34425 7757 34459
rect 7791 34456 7803 34459
rect 7926 34456 7932 34468
rect 7791 34428 7932 34456
rect 7791 34425 7803 34428
rect 7745 34419 7803 34425
rect 6641 34391 6699 34397
rect 6641 34357 6653 34391
rect 6687 34388 6699 34391
rect 6730 34388 6736 34400
rect 6687 34360 6736 34388
rect 6687 34357 6699 34360
rect 6641 34351 6699 34357
rect 6730 34348 6736 34360
rect 6788 34348 6794 34400
rect 7006 34388 7012 34400
rect 6967 34360 7012 34388
rect 7006 34348 7012 34360
rect 7064 34348 7070 34400
rect 7469 34391 7527 34397
rect 7469 34357 7481 34391
rect 7515 34388 7527 34391
rect 7760 34388 7788 34419
rect 7926 34416 7932 34428
rect 7984 34416 7990 34468
rect 8110 34416 8116 34468
rect 8168 34456 8174 34468
rect 8941 34459 8999 34465
rect 8941 34456 8953 34459
rect 8168 34428 8953 34456
rect 8168 34416 8174 34428
rect 8941 34425 8953 34428
rect 8987 34425 8999 34459
rect 8941 34419 8999 34425
rect 10413 34459 10471 34465
rect 10413 34425 10425 34459
rect 10459 34425 10471 34459
rect 10413 34419 10471 34425
rect 7515 34360 7788 34388
rect 7515 34357 7527 34360
rect 7469 34351 7527 34357
rect 8202 34348 8208 34400
rect 8260 34388 8266 34400
rect 8665 34391 8723 34397
rect 8665 34388 8677 34391
rect 8260 34360 8677 34388
rect 8260 34348 8266 34360
rect 8665 34357 8677 34360
rect 8711 34388 8723 34391
rect 9490 34388 9496 34400
rect 8711 34360 9496 34388
rect 8711 34357 8723 34360
rect 8665 34351 8723 34357
rect 9490 34348 9496 34360
rect 9548 34348 9554 34400
rect 10137 34391 10195 34397
rect 10137 34357 10149 34391
rect 10183 34388 10195 34391
rect 10226 34388 10232 34400
rect 10183 34360 10232 34388
rect 10183 34357 10195 34360
rect 10137 34351 10195 34357
rect 10226 34348 10232 34360
rect 10284 34388 10290 34400
rect 10428 34388 10456 34419
rect 10686 34416 10692 34468
rect 10744 34456 10750 34468
rect 12452 34456 12480 34484
rect 10744 34428 12480 34456
rect 10744 34416 10750 34428
rect 10594 34388 10600 34400
rect 10284 34360 10600 34388
rect 10284 34348 10290 34360
rect 10594 34348 10600 34360
rect 10652 34388 10658 34400
rect 11241 34391 11299 34397
rect 11241 34388 11253 34391
rect 10652 34360 11253 34388
rect 10652 34348 10658 34360
rect 11241 34357 11253 34360
rect 11287 34357 11299 34391
rect 11241 34351 11299 34357
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 5307 34187 5365 34193
rect 5307 34153 5319 34187
rect 5353 34184 5365 34187
rect 8110 34184 8116 34196
rect 5353 34156 8116 34184
rect 5353 34153 5365 34156
rect 5307 34147 5365 34153
rect 8110 34144 8116 34156
rect 8168 34144 8174 34196
rect 9950 34144 9956 34196
rect 10008 34184 10014 34196
rect 10045 34187 10103 34193
rect 10045 34184 10057 34187
rect 10008 34156 10057 34184
rect 10008 34144 10014 34156
rect 10045 34153 10057 34156
rect 10091 34153 10103 34187
rect 10045 34147 10103 34153
rect 13173 34187 13231 34193
rect 13173 34153 13185 34187
rect 13219 34184 13231 34187
rect 15562 34184 15568 34196
rect 13219 34156 15568 34184
rect 13219 34153 13231 34156
rect 13173 34147 13231 34153
rect 15562 34144 15568 34156
rect 15620 34144 15626 34196
rect 6362 34116 6368 34128
rect 6323 34088 6368 34116
rect 6362 34076 6368 34088
rect 6420 34076 6426 34128
rect 7926 34116 7932 34128
rect 7887 34088 7932 34116
rect 7926 34076 7932 34088
rect 7984 34076 7990 34128
rect 8478 34116 8484 34128
rect 8439 34088 8484 34116
rect 8478 34076 8484 34088
rect 8536 34076 8542 34128
rect 10962 34116 10968 34128
rect 10612 34088 10968 34116
rect 5169 34051 5227 34057
rect 5169 34017 5181 34051
rect 5215 34048 5227 34051
rect 5258 34048 5264 34060
rect 5215 34020 5264 34048
rect 5215 34017 5227 34020
rect 5169 34011 5227 34017
rect 5258 34008 5264 34020
rect 5316 34008 5322 34060
rect 10612 34057 10640 34088
rect 10962 34076 10968 34088
rect 11020 34116 11026 34128
rect 11609 34119 11667 34125
rect 11609 34116 11621 34119
rect 11020 34088 11621 34116
rect 11020 34076 11026 34088
rect 11609 34085 11621 34088
rect 11655 34085 11667 34119
rect 11609 34079 11667 34085
rect 10597 34051 10655 34057
rect 10597 34017 10609 34051
rect 10643 34017 10655 34051
rect 10597 34011 10655 34017
rect 12158 34008 12164 34060
rect 12216 34048 12222 34060
rect 12434 34048 12440 34060
rect 12216 34020 12440 34048
rect 12216 34008 12222 34020
rect 12434 34008 12440 34020
rect 12492 34048 12498 34060
rect 12989 34051 13047 34057
rect 12989 34048 13001 34051
rect 12492 34020 13001 34048
rect 12492 34008 12498 34020
rect 12989 34017 13001 34020
rect 13035 34048 13047 34051
rect 13446 34048 13452 34060
rect 13035 34020 13452 34048
rect 13035 34017 13047 34020
rect 12989 34011 13047 34017
rect 13446 34008 13452 34020
rect 13504 34008 13510 34060
rect 6273 33983 6331 33989
rect 6273 33980 6285 33983
rect 6196 33952 6285 33980
rect 6196 33924 6224 33952
rect 6273 33949 6285 33952
rect 6319 33949 6331 33983
rect 7834 33980 7840 33992
rect 7795 33952 7840 33980
rect 6273 33943 6331 33949
rect 7834 33940 7840 33952
rect 7892 33940 7898 33992
rect 9677 33983 9735 33989
rect 9677 33949 9689 33983
rect 9723 33980 9735 33983
rect 9766 33980 9772 33992
rect 9723 33952 9772 33980
rect 9723 33949 9735 33952
rect 9677 33943 9735 33949
rect 9766 33940 9772 33952
rect 9824 33940 9830 33992
rect 11330 33940 11336 33992
rect 11388 33980 11394 33992
rect 11517 33983 11575 33989
rect 11517 33980 11529 33983
rect 11388 33952 11529 33980
rect 11388 33940 11394 33952
rect 11517 33949 11529 33952
rect 11563 33949 11575 33983
rect 11517 33943 11575 33949
rect 11793 33983 11851 33989
rect 11793 33949 11805 33983
rect 11839 33949 11851 33983
rect 11793 33943 11851 33949
rect 6178 33872 6184 33924
rect 6236 33872 6242 33924
rect 6825 33915 6883 33921
rect 6825 33881 6837 33915
rect 6871 33912 6883 33915
rect 8478 33912 8484 33924
rect 6871 33884 8484 33912
rect 6871 33881 6883 33884
rect 6825 33875 6883 33881
rect 8478 33872 8484 33884
rect 8536 33872 8542 33924
rect 11054 33872 11060 33924
rect 11112 33912 11118 33924
rect 11808 33912 11836 33943
rect 11112 33884 11836 33912
rect 11112 33872 11118 33884
rect 7558 33844 7564 33856
rect 7519 33816 7564 33844
rect 7558 33804 7564 33816
rect 7616 33804 7622 33856
rect 10502 33804 10508 33856
rect 10560 33844 10566 33856
rect 10965 33847 11023 33853
rect 10965 33844 10977 33847
rect 10560 33816 10977 33844
rect 10560 33804 10566 33816
rect 10965 33813 10977 33816
rect 11011 33844 11023 33847
rect 12158 33844 12164 33856
rect 11011 33816 12164 33844
rect 11011 33813 11023 33816
rect 10965 33807 11023 33813
rect 12158 33804 12164 33816
rect 12216 33804 12222 33856
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 4847 33643 4905 33649
rect 4847 33609 4859 33643
rect 4893 33640 4905 33643
rect 6086 33640 6092 33652
rect 4893 33612 6092 33640
rect 4893 33609 4905 33612
rect 4847 33603 4905 33609
rect 6086 33600 6092 33612
rect 6144 33600 6150 33652
rect 6362 33600 6368 33652
rect 6420 33640 6426 33652
rect 6549 33643 6607 33649
rect 6549 33640 6561 33643
rect 6420 33612 6561 33640
rect 6420 33600 6426 33612
rect 6549 33609 6561 33612
rect 6595 33640 6607 33643
rect 7193 33643 7251 33649
rect 7193 33640 7205 33643
rect 6595 33612 7205 33640
rect 6595 33609 6607 33612
rect 6549 33603 6607 33609
rect 7193 33609 7205 33612
rect 7239 33640 7251 33643
rect 7285 33643 7343 33649
rect 7285 33640 7297 33643
rect 7239 33612 7297 33640
rect 7239 33609 7251 33612
rect 7193 33603 7251 33609
rect 7285 33609 7297 33612
rect 7331 33609 7343 33643
rect 10226 33640 10232 33652
rect 10187 33612 10232 33640
rect 7285 33603 7343 33609
rect 10226 33600 10232 33612
rect 10284 33600 10290 33652
rect 10962 33640 10968 33652
rect 10923 33612 10968 33640
rect 10962 33600 10968 33612
rect 11020 33600 11026 33652
rect 11241 33643 11299 33649
rect 11241 33609 11253 33643
rect 11287 33640 11299 33643
rect 11514 33640 11520 33652
rect 11287 33612 11520 33640
rect 11287 33609 11299 33612
rect 11241 33603 11299 33609
rect 11514 33600 11520 33612
rect 11572 33600 11578 33652
rect 13446 33640 13452 33652
rect 13407 33612 13452 33640
rect 13446 33600 13452 33612
rect 13504 33600 13510 33652
rect 10410 33532 10416 33584
rect 10468 33572 10474 33584
rect 12161 33575 12219 33581
rect 12161 33572 12173 33575
rect 10468 33544 12173 33572
rect 10468 33532 10474 33544
rect 12161 33541 12173 33544
rect 12207 33541 12219 33575
rect 12161 33535 12219 33541
rect 5859 33507 5917 33513
rect 5859 33473 5871 33507
rect 5905 33504 5917 33507
rect 7558 33504 7564 33516
rect 5905 33476 7564 33504
rect 5905 33473 5917 33476
rect 5859 33467 5917 33473
rect 7558 33464 7564 33476
rect 7616 33464 7622 33516
rect 8018 33464 8024 33516
rect 8076 33504 8082 33516
rect 8205 33507 8263 33513
rect 8205 33504 8217 33507
rect 8076 33476 8217 33504
rect 8076 33464 8082 33476
rect 8205 33473 8217 33476
rect 8251 33504 8263 33507
rect 8294 33504 8300 33516
rect 8251 33476 8300 33504
rect 8251 33473 8263 33476
rect 8205 33467 8263 33473
rect 8294 33464 8300 33476
rect 8352 33464 8358 33516
rect 8849 33507 8907 33513
rect 8849 33473 8861 33507
rect 8895 33504 8907 33507
rect 9766 33504 9772 33516
rect 8895 33476 9772 33504
rect 8895 33473 8907 33476
rect 8849 33467 8907 33473
rect 9766 33464 9772 33476
rect 9824 33464 9830 33516
rect 658 33396 664 33448
rect 716 33436 722 33448
rect 4776 33439 4834 33445
rect 4776 33436 4788 33439
rect 716 33408 4788 33436
rect 716 33396 722 33408
rect 4776 33405 4788 33408
rect 4822 33436 4834 33439
rect 5772 33439 5830 33445
rect 4822 33408 5672 33436
rect 4822 33405 4834 33408
rect 4776 33399 4834 33405
rect 5258 33300 5264 33312
rect 5219 33272 5264 33300
rect 5258 33260 5264 33272
rect 5316 33260 5322 33312
rect 5644 33309 5672 33408
rect 5772 33405 5784 33439
rect 5818 33436 5830 33439
rect 9306 33436 9312 33448
rect 5818 33408 6316 33436
rect 9267 33408 9312 33436
rect 5818 33405 5830 33408
rect 5772 33399 5830 33405
rect 5629 33303 5687 33309
rect 5629 33269 5641 33303
rect 5675 33300 5687 33303
rect 5994 33300 6000 33312
rect 5675 33272 6000 33300
rect 5675 33269 5687 33272
rect 5629 33263 5687 33269
rect 5994 33260 6000 33272
rect 6052 33260 6058 33312
rect 6288 33309 6316 33408
rect 9306 33396 9312 33408
rect 9364 33396 9370 33448
rect 11057 33439 11115 33445
rect 11057 33405 11069 33439
rect 11103 33405 11115 33439
rect 12176 33436 12204 33535
rect 12526 33504 12532 33516
rect 12487 33476 12532 33504
rect 12526 33464 12532 33476
rect 12584 33464 12590 33516
rect 12802 33504 12808 33516
rect 12763 33476 12808 33504
rect 12802 33464 12808 33476
rect 12860 33464 12866 33516
rect 12176 33408 12388 33436
rect 11057 33399 11115 33405
rect 7193 33371 7251 33377
rect 7193 33337 7205 33371
rect 7239 33368 7251 33371
rect 7650 33368 7656 33380
rect 7239 33340 7656 33368
rect 7239 33337 7251 33340
rect 7193 33331 7251 33337
rect 7650 33328 7656 33340
rect 7708 33328 7714 33380
rect 9671 33371 9729 33377
rect 9671 33368 9683 33371
rect 9646 33337 9683 33368
rect 9717 33368 9729 33371
rect 9950 33368 9956 33380
rect 9717 33340 9956 33368
rect 9717 33337 9729 33340
rect 9646 33331 9729 33337
rect 9646 33312 9674 33331
rect 9950 33328 9956 33340
rect 10008 33368 10014 33380
rect 10505 33371 10563 33377
rect 10505 33368 10517 33371
rect 10008 33340 10517 33368
rect 10008 33328 10014 33340
rect 10505 33337 10517 33340
rect 10551 33337 10563 33371
rect 10505 33331 10563 33337
rect 10778 33328 10784 33380
rect 10836 33368 10842 33380
rect 11072 33368 11100 33399
rect 11701 33371 11759 33377
rect 11701 33368 11713 33371
rect 10836 33340 11713 33368
rect 10836 33328 10842 33340
rect 11701 33337 11713 33340
rect 11747 33368 11759 33371
rect 12250 33368 12256 33380
rect 11747 33340 12256 33368
rect 11747 33337 11759 33340
rect 11701 33331 11759 33337
rect 12250 33328 12256 33340
rect 12308 33328 12314 33380
rect 12360 33368 12388 33408
rect 12621 33371 12679 33377
rect 12621 33368 12633 33371
rect 12360 33340 12633 33368
rect 12621 33337 12633 33340
rect 12667 33337 12679 33371
rect 12621 33331 12679 33337
rect 6273 33303 6331 33309
rect 6273 33269 6285 33303
rect 6319 33300 6331 33303
rect 7006 33300 7012 33312
rect 6319 33272 7012 33300
rect 6319 33269 6331 33272
rect 6273 33263 6331 33269
rect 7006 33260 7012 33272
rect 7064 33300 7070 33312
rect 8202 33300 8208 33312
rect 7064 33272 8208 33300
rect 7064 33260 7070 33272
rect 8202 33260 8208 33272
rect 8260 33260 8266 33312
rect 9217 33303 9275 33309
rect 9217 33269 9229 33303
rect 9263 33300 9275 33303
rect 9582 33300 9588 33312
rect 9263 33272 9588 33300
rect 9263 33269 9275 33272
rect 9217 33263 9275 33269
rect 9582 33260 9588 33272
rect 9640 33272 9674 33312
rect 9640 33260 9646 33272
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 5859 33099 5917 33105
rect 5859 33065 5871 33099
rect 5905 33096 5917 33099
rect 6178 33096 6184 33108
rect 5905 33068 6184 33096
rect 5905 33065 5917 33068
rect 5859 33059 5917 33065
rect 6178 33056 6184 33068
rect 6236 33056 6242 33108
rect 7098 33096 7104 33108
rect 7059 33068 7104 33096
rect 7098 33056 7104 33068
rect 7156 33056 7162 33108
rect 7650 33096 7656 33108
rect 7611 33068 7656 33096
rect 7650 33056 7656 33068
rect 7708 33056 7714 33108
rect 7926 33096 7932 33108
rect 7887 33068 7932 33096
rect 7926 33056 7932 33068
rect 7984 33056 7990 33108
rect 9950 33056 9956 33108
rect 10008 33096 10014 33108
rect 10045 33099 10103 33105
rect 10045 33096 10057 33099
rect 10008 33068 10057 33096
rect 10008 33056 10014 33068
rect 10045 33065 10057 33068
rect 10091 33065 10103 33099
rect 10045 33059 10103 33065
rect 10410 33056 10416 33108
rect 10468 33096 10474 33108
rect 10597 33099 10655 33105
rect 10597 33096 10609 33099
rect 10468 33068 10609 33096
rect 10468 33056 10474 33068
rect 10597 33065 10609 33068
rect 10643 33065 10655 33099
rect 10597 33059 10655 33065
rect 11514 33056 11520 33108
rect 11572 33096 11578 33108
rect 12526 33096 12532 33108
rect 11572 33068 11836 33096
rect 12487 33068 12532 33096
rect 11572 33056 11578 33068
rect 7834 32988 7840 33040
rect 7892 33028 7898 33040
rect 8297 33031 8355 33037
rect 8297 33028 8309 33031
rect 7892 33000 8309 33028
rect 7892 32988 7898 33000
rect 8297 32997 8309 33000
rect 8343 33028 8355 33031
rect 8619 33031 8677 33037
rect 8619 33028 8631 33031
rect 8343 33000 8631 33028
rect 8343 32997 8355 33000
rect 8297 32991 8355 32997
rect 8619 32997 8631 33000
rect 8665 32997 8677 33031
rect 8619 32991 8677 32997
rect 10962 32988 10968 33040
rect 11020 33028 11026 33040
rect 11609 33031 11667 33037
rect 11609 33028 11621 33031
rect 11020 33000 11621 33028
rect 11020 32988 11026 33000
rect 11609 32997 11621 33000
rect 11655 33028 11667 33031
rect 11698 33028 11704 33040
rect 11655 33000 11704 33028
rect 11655 32997 11667 33000
rect 11609 32991 11667 32997
rect 11698 32988 11704 33000
rect 11756 32988 11762 33040
rect 11808 33028 11836 33068
rect 12526 33056 12532 33068
rect 12584 33056 12590 33108
rect 12161 33031 12219 33037
rect 12161 33028 12173 33031
rect 11808 33000 12173 33028
rect 12161 32997 12173 33000
rect 12207 33028 12219 33031
rect 12802 33028 12808 33040
rect 12207 33000 12808 33028
rect 12207 32997 12219 33000
rect 12161 32991 12219 32997
rect 12802 32988 12808 33000
rect 12860 32988 12866 33040
rect 4062 32920 4068 32972
rect 4120 32960 4126 32972
rect 5718 32960 5724 32972
rect 5776 32969 5782 32972
rect 5776 32963 5814 32969
rect 4120 32932 5724 32960
rect 4120 32920 4126 32932
rect 5718 32920 5724 32932
rect 5802 32929 5814 32963
rect 8516 32963 8574 32969
rect 8516 32960 8528 32963
rect 5776 32923 5814 32929
rect 8312 32932 8528 32960
rect 5776 32920 5782 32923
rect 8312 32904 8340 32932
rect 8516 32929 8528 32932
rect 8562 32960 8574 32963
rect 12986 32960 12992 32972
rect 8562 32932 11376 32960
rect 12947 32932 12992 32960
rect 8562 32929 8574 32932
rect 8516 32923 8574 32929
rect 6733 32895 6791 32901
rect 6733 32861 6745 32895
rect 6779 32892 6791 32895
rect 7374 32892 7380 32904
rect 6779 32864 7380 32892
rect 6779 32861 6791 32864
rect 6733 32855 6791 32861
rect 7374 32852 7380 32864
rect 7432 32852 7438 32904
rect 8294 32852 8300 32904
rect 8352 32852 8358 32904
rect 9677 32895 9735 32901
rect 9677 32861 9689 32895
rect 9723 32892 9735 32895
rect 10410 32892 10416 32904
rect 9723 32864 10416 32892
rect 9723 32861 9735 32864
rect 9677 32855 9735 32861
rect 10410 32852 10416 32864
rect 10468 32852 10474 32904
rect 5258 32784 5264 32836
rect 5316 32824 5322 32836
rect 10778 32824 10784 32836
rect 5316 32796 10784 32824
rect 5316 32784 5322 32796
rect 10778 32784 10784 32796
rect 10836 32784 10842 32836
rect 11348 32824 11376 32932
rect 12986 32920 12992 32932
rect 13044 32920 13050 32972
rect 11514 32892 11520 32904
rect 11475 32864 11520 32892
rect 11514 32852 11520 32864
rect 11572 32852 11578 32904
rect 12434 32824 12440 32836
rect 11348 32796 12440 32824
rect 12434 32784 12440 32796
rect 12492 32784 12498 32836
rect 8754 32716 8760 32768
rect 8812 32756 8818 32768
rect 8941 32759 8999 32765
rect 8941 32756 8953 32759
rect 8812 32728 8953 32756
rect 8812 32716 8818 32728
rect 8941 32725 8953 32728
rect 8987 32725 8999 32759
rect 9306 32756 9312 32768
rect 9267 32728 9312 32756
rect 8941 32719 8999 32725
rect 9306 32716 9312 32728
rect 9364 32716 9370 32768
rect 11330 32756 11336 32768
rect 11243 32728 11336 32756
rect 11330 32716 11336 32728
rect 11388 32756 11394 32768
rect 13127 32759 13185 32765
rect 13127 32756 13139 32759
rect 11388 32728 13139 32756
rect 11388 32716 11394 32728
rect 13127 32725 13139 32728
rect 13173 32725 13185 32759
rect 13127 32719 13185 32725
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 5718 32552 5724 32564
rect 5679 32524 5724 32552
rect 5718 32512 5724 32524
rect 5776 32552 5782 32564
rect 7466 32552 7472 32564
rect 5776 32524 7472 32552
rect 5776 32512 5782 32524
rect 7466 32512 7472 32524
rect 7524 32512 7530 32564
rect 7745 32555 7803 32561
rect 7745 32521 7757 32555
rect 7791 32552 7803 32555
rect 7926 32552 7932 32564
rect 7791 32524 7932 32552
rect 7791 32521 7803 32524
rect 7745 32515 7803 32521
rect 7926 32512 7932 32524
rect 7984 32512 7990 32564
rect 8294 32512 8300 32564
rect 8352 32552 8358 32564
rect 8389 32555 8447 32561
rect 8389 32552 8401 32555
rect 8352 32524 8401 32552
rect 8352 32512 8358 32524
rect 8389 32521 8401 32524
rect 8435 32521 8447 32555
rect 9490 32552 9496 32564
rect 9451 32524 9496 32552
rect 8389 32515 8447 32521
rect 9490 32512 9496 32524
rect 9548 32512 9554 32564
rect 11698 32552 11704 32564
rect 11659 32524 11704 32552
rect 11698 32512 11704 32524
rect 11756 32512 11762 32564
rect 12158 32512 12164 32564
rect 12216 32552 12222 32564
rect 12575 32555 12633 32561
rect 12575 32552 12587 32555
rect 12216 32524 12587 32552
rect 12216 32512 12222 32524
rect 12575 32521 12587 32524
rect 12621 32521 12633 32555
rect 12575 32515 12633 32521
rect 6822 32444 6828 32496
rect 6880 32484 6886 32496
rect 7834 32484 7840 32496
rect 6880 32456 7840 32484
rect 6880 32444 6886 32456
rect 7834 32444 7840 32456
rect 7892 32484 7898 32496
rect 12253 32487 12311 32493
rect 12253 32484 12265 32487
rect 7892 32456 12265 32484
rect 7892 32444 7898 32456
rect 12253 32453 12265 32456
rect 12299 32453 12311 32487
rect 12253 32447 12311 32453
rect 6273 32419 6331 32425
rect 6273 32385 6285 32419
rect 6319 32416 6331 32419
rect 6641 32419 6699 32425
rect 6641 32416 6653 32419
rect 6319 32388 6653 32416
rect 6319 32385 6331 32388
rect 6273 32379 6331 32385
rect 6641 32385 6653 32388
rect 6687 32416 6699 32419
rect 7098 32416 7104 32428
rect 6687 32388 7104 32416
rect 6687 32385 6699 32388
rect 6641 32379 6699 32385
rect 7098 32376 7104 32388
rect 7156 32416 7162 32428
rect 8573 32419 8631 32425
rect 7156 32388 7236 32416
rect 7156 32376 7162 32388
rect 6822 32348 6828 32360
rect 6783 32320 6828 32348
rect 6822 32308 6828 32320
rect 6880 32308 6886 32360
rect 7208 32221 7236 32388
rect 8573 32385 8585 32419
rect 8619 32416 8631 32419
rect 8754 32416 8760 32428
rect 8619 32388 8760 32416
rect 8619 32385 8631 32388
rect 8573 32379 8631 32385
rect 8754 32376 8760 32388
rect 8812 32376 8818 32428
rect 10318 32348 10324 32360
rect 10279 32320 10324 32348
rect 10318 32308 10324 32320
rect 10376 32308 10382 32360
rect 10781 32351 10839 32357
rect 10781 32348 10793 32351
rect 10520 32320 10793 32348
rect 8113 32283 8171 32289
rect 8113 32249 8125 32283
rect 8159 32280 8171 32283
rect 8935 32283 8993 32289
rect 8935 32280 8947 32283
rect 8159 32252 8947 32280
rect 8159 32249 8171 32252
rect 8113 32243 8171 32249
rect 8935 32249 8947 32252
rect 8981 32280 8993 32283
rect 10226 32280 10232 32292
rect 8981 32252 9628 32280
rect 10139 32252 10232 32280
rect 8981 32249 8993 32252
rect 8935 32243 8993 32249
rect 7193 32215 7251 32221
rect 7193 32181 7205 32215
rect 7239 32212 7251 32215
rect 7282 32212 7288 32224
rect 7239 32184 7288 32212
rect 7239 32181 7251 32184
rect 7193 32175 7251 32181
rect 7282 32172 7288 32184
rect 7340 32212 7346 32224
rect 8128 32212 8156 32243
rect 9600 32224 9628 32252
rect 10226 32240 10232 32252
rect 10284 32280 10290 32292
rect 10520 32280 10548 32320
rect 10781 32317 10793 32320
rect 10827 32317 10839 32351
rect 12268 32348 12296 32447
rect 12472 32351 12530 32357
rect 12472 32348 12484 32351
rect 12268 32320 12484 32348
rect 10781 32311 10839 32317
rect 12472 32317 12484 32320
rect 12518 32317 12530 32351
rect 12472 32311 12530 32317
rect 10284 32252 10548 32280
rect 10284 32240 10290 32252
rect 7340 32184 8156 32212
rect 7340 32172 7346 32184
rect 9582 32172 9588 32224
rect 9640 32212 9646 32224
rect 9769 32215 9827 32221
rect 9769 32212 9781 32215
rect 9640 32184 9781 32212
rect 9640 32172 9646 32184
rect 9769 32181 9781 32184
rect 9815 32181 9827 32215
rect 10410 32212 10416 32224
rect 10371 32184 10416 32212
rect 9769 32175 9827 32181
rect 10410 32172 10416 32184
rect 10468 32212 10474 32224
rect 11333 32215 11391 32221
rect 11333 32212 11345 32215
rect 10468 32184 11345 32212
rect 10468 32172 10474 32184
rect 11333 32181 11345 32184
rect 11379 32181 11391 32215
rect 11333 32175 11391 32181
rect 12342 32172 12348 32224
rect 12400 32212 12406 32224
rect 12986 32212 12992 32224
rect 12400 32184 12992 32212
rect 12400 32172 12406 32184
rect 12986 32172 12992 32184
rect 13044 32172 13050 32224
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 9766 32008 9772 32020
rect 9727 31980 9772 32008
rect 9766 31968 9772 31980
rect 9824 31968 9830 32020
rect 11379 32011 11437 32017
rect 11379 31977 11391 32011
rect 11425 32008 11437 32011
rect 11514 32008 11520 32020
rect 11425 31980 11520 32008
rect 11425 31977 11437 31980
rect 11379 31971 11437 31977
rect 11514 31968 11520 31980
rect 11572 32008 11578 32020
rect 11701 32011 11759 32017
rect 11701 32008 11713 32011
rect 11572 31980 11713 32008
rect 11572 31968 11578 31980
rect 11701 31977 11713 31980
rect 11747 31977 11759 32011
rect 11701 31971 11759 31977
rect 6822 31940 6828 31952
rect 6783 31912 6828 31940
rect 6822 31900 6828 31912
rect 6880 31940 6886 31952
rect 7469 31943 7527 31949
rect 7469 31940 7481 31943
rect 6880 31912 7481 31940
rect 6880 31900 6886 31912
rect 7469 31909 7481 31912
rect 7515 31909 7527 31943
rect 8389 31943 8447 31949
rect 7469 31903 7527 31909
rect 7852 31912 8248 31940
rect 5534 31832 5540 31884
rect 5592 31872 5598 31884
rect 6089 31875 6147 31881
rect 6089 31872 6101 31875
rect 5592 31844 6101 31872
rect 5592 31832 5598 31844
rect 6089 31841 6101 31844
rect 6135 31841 6147 31875
rect 6638 31872 6644 31884
rect 6599 31844 6644 31872
rect 6089 31835 6147 31841
rect 6104 31736 6132 31835
rect 6638 31832 6644 31844
rect 6696 31832 6702 31884
rect 7650 31832 7656 31884
rect 7708 31872 7714 31884
rect 7852 31881 7880 31912
rect 7837 31875 7895 31881
rect 7837 31872 7849 31875
rect 7708 31844 7849 31872
rect 7708 31832 7714 31844
rect 7837 31841 7849 31844
rect 7883 31841 7895 31875
rect 8110 31872 8116 31884
rect 8071 31844 8116 31872
rect 7837 31835 7895 31841
rect 8110 31832 8116 31844
rect 8168 31832 8174 31884
rect 8220 31872 8248 31912
rect 8389 31909 8401 31943
rect 8435 31940 8447 31943
rect 8754 31940 8760 31952
rect 8435 31912 8760 31940
rect 8435 31909 8447 31912
rect 8389 31903 8447 31909
rect 8754 31900 8760 31912
rect 8812 31900 8818 31952
rect 9950 31872 9956 31884
rect 8220 31844 9674 31872
rect 9911 31844 9956 31872
rect 9646 31804 9674 31844
rect 9950 31832 9956 31844
rect 10008 31832 10014 31884
rect 10226 31872 10232 31884
rect 10187 31844 10232 31872
rect 10226 31832 10232 31844
rect 10284 31832 10290 31884
rect 11238 31872 11244 31884
rect 11199 31844 11244 31872
rect 11238 31832 11244 31844
rect 11296 31832 11302 31884
rect 11514 31832 11520 31884
rect 11572 31872 11578 31884
rect 15470 31872 15476 31884
rect 11572 31844 15476 31872
rect 11572 31832 11578 31844
rect 15470 31832 15476 31844
rect 15528 31832 15534 31884
rect 9968 31804 9996 31832
rect 9646 31776 9996 31804
rect 10318 31736 10324 31748
rect 6104 31708 10324 31736
rect 10318 31696 10324 31708
rect 10376 31736 10382 31748
rect 10689 31739 10747 31745
rect 10689 31736 10701 31739
rect 10376 31708 10701 31736
rect 10376 31696 10382 31708
rect 10689 31705 10701 31708
rect 10735 31705 10747 31739
rect 10689 31699 10747 31705
rect 7193 31671 7251 31677
rect 7193 31637 7205 31671
rect 7239 31668 7251 31671
rect 7374 31668 7380 31680
rect 7239 31640 7380 31668
rect 7239 31637 7251 31640
rect 7193 31631 7251 31637
rect 7374 31628 7380 31640
rect 7432 31628 7438 31680
rect 8662 31668 8668 31680
rect 8623 31640 8668 31668
rect 8662 31628 8668 31640
rect 8720 31628 8726 31680
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 9769 31467 9827 31473
rect 9769 31433 9781 31467
rect 9815 31464 9827 31467
rect 10226 31464 10232 31476
rect 9815 31436 10232 31464
rect 9815 31433 9827 31436
rect 9769 31427 9827 31433
rect 6932 31368 7512 31396
rect 6932 31272 6960 31368
rect 7374 31328 7380 31340
rect 7335 31300 7380 31328
rect 7374 31288 7380 31300
rect 7432 31288 7438 31340
rect 6914 31260 6920 31272
rect 6875 31232 6920 31260
rect 6914 31220 6920 31232
rect 6972 31220 6978 31272
rect 7285 31263 7343 31269
rect 7285 31229 7297 31263
rect 7331 31229 7343 31263
rect 7484 31260 7512 31368
rect 9306 31328 9312 31340
rect 9267 31300 9312 31328
rect 9306 31288 9312 31300
rect 9364 31288 9370 31340
rect 8662 31260 8668 31272
rect 7484 31232 8668 31260
rect 7285 31223 7343 31229
rect 5534 31084 5540 31136
rect 5592 31124 5598 31136
rect 5721 31127 5779 31133
rect 5721 31124 5733 31127
rect 5592 31096 5733 31124
rect 5592 31084 5598 31096
rect 5721 31093 5733 31096
rect 5767 31093 5779 31127
rect 5721 31087 5779 31093
rect 6181 31127 6239 31133
rect 6181 31093 6193 31127
rect 6227 31124 6239 31127
rect 6638 31124 6644 31136
rect 6227 31096 6644 31124
rect 6227 31093 6239 31096
rect 6181 31087 6239 31093
rect 6638 31084 6644 31096
rect 6696 31124 6702 31136
rect 7300 31124 7328 31223
rect 8662 31220 8668 31232
rect 8720 31220 8726 31272
rect 9217 31263 9275 31269
rect 9217 31229 9229 31263
rect 9263 31260 9275 31263
rect 9784 31260 9812 31427
rect 10226 31424 10232 31436
rect 10284 31424 10290 31476
rect 9950 31356 9956 31408
rect 10008 31396 10014 31408
rect 10137 31399 10195 31405
rect 10137 31396 10149 31399
rect 10008 31368 10149 31396
rect 10008 31356 10014 31368
rect 10137 31365 10149 31368
rect 10183 31396 10195 31399
rect 12066 31396 12072 31408
rect 10183 31368 12072 31396
rect 10183 31365 10195 31368
rect 10137 31359 10195 31365
rect 12066 31356 12072 31368
rect 12124 31356 12130 31408
rect 10689 31331 10747 31337
rect 10689 31297 10701 31331
rect 10735 31328 10747 31331
rect 11054 31328 11060 31340
rect 10735 31300 11060 31328
rect 10735 31297 10747 31300
rect 10689 31291 10747 31297
rect 11054 31288 11060 31300
rect 11112 31288 11118 31340
rect 9263 31232 9812 31260
rect 9263 31229 9275 31232
rect 9217 31223 9275 31229
rect 8573 31195 8631 31201
rect 8573 31161 8585 31195
rect 8619 31192 8631 31195
rect 9232 31192 9260 31223
rect 8619 31164 9260 31192
rect 10781 31195 10839 31201
rect 8619 31161 8631 31164
rect 8573 31155 8631 31161
rect 8680 31136 8708 31164
rect 10781 31161 10793 31195
rect 10827 31192 10839 31195
rect 10962 31192 10968 31204
rect 10827 31164 10968 31192
rect 10827 31161 10839 31164
rect 10781 31155 10839 31161
rect 7837 31127 7895 31133
rect 7837 31124 7849 31127
rect 6696 31096 7849 31124
rect 6696 31084 6702 31096
rect 7837 31093 7849 31096
rect 7883 31124 7895 31127
rect 8110 31124 8116 31136
rect 7883 31096 8116 31124
rect 7883 31093 7895 31096
rect 7837 31087 7895 31093
rect 8110 31084 8116 31096
rect 8168 31084 8174 31136
rect 8662 31084 8668 31136
rect 8720 31084 8726 31136
rect 10505 31127 10563 31133
rect 10505 31093 10517 31127
rect 10551 31124 10563 31127
rect 10796 31124 10824 31155
rect 10962 31152 10968 31164
rect 11020 31152 11026 31204
rect 11333 31195 11391 31201
rect 11333 31161 11345 31195
rect 11379 31192 11391 31195
rect 12158 31192 12164 31204
rect 11379 31164 12164 31192
rect 11379 31161 11391 31164
rect 11333 31155 11391 31161
rect 12158 31152 12164 31164
rect 12216 31152 12222 31204
rect 10551 31096 10824 31124
rect 10551 31093 10563 31096
rect 10505 31087 10563 31093
rect 11238 31084 11244 31136
rect 11296 31124 11302 31136
rect 11701 31127 11759 31133
rect 11701 31124 11713 31127
rect 11296 31096 11713 31124
rect 11296 31084 11302 31096
rect 11701 31093 11713 31096
rect 11747 31124 11759 31127
rect 12434 31124 12440 31136
rect 11747 31096 12440 31124
rect 11747 31093 11759 31096
rect 11701 31087 11759 31093
rect 12434 31084 12440 31096
rect 12492 31084 12498 31136
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 7650 30920 7656 30932
rect 7611 30892 7656 30920
rect 7650 30880 7656 30892
rect 7708 30880 7714 30932
rect 8018 30880 8024 30932
rect 8076 30920 8082 30932
rect 8076 30892 8156 30920
rect 8076 30880 8082 30892
rect 8128 30861 8156 30892
rect 8570 30880 8576 30932
rect 8628 30920 8634 30932
rect 9401 30923 9459 30929
rect 9401 30920 9413 30923
rect 8628 30892 9413 30920
rect 8628 30880 8634 30892
rect 8113 30855 8171 30861
rect 8113 30821 8125 30855
rect 8159 30821 8171 30855
rect 8113 30815 8171 30821
rect 8205 30855 8263 30861
rect 8205 30821 8217 30855
rect 8251 30852 8263 30855
rect 8294 30852 8300 30864
rect 8251 30824 8300 30852
rect 8251 30821 8263 30824
rect 8205 30815 8263 30821
rect 8294 30812 8300 30824
rect 8352 30812 8358 30864
rect 6730 30744 6736 30796
rect 6788 30784 6794 30796
rect 6788 30756 7144 30784
rect 6788 30744 6794 30756
rect 7116 30728 7144 30756
rect 5258 30676 5264 30728
rect 5316 30716 5322 30728
rect 7009 30719 7067 30725
rect 7009 30716 7021 30719
rect 5316 30688 7021 30716
rect 5316 30676 5322 30688
rect 7009 30685 7021 30688
rect 7055 30685 7067 30719
rect 7009 30679 7067 30685
rect 7098 30676 7104 30728
rect 7156 30716 7162 30728
rect 8389 30719 8447 30725
rect 8389 30716 8401 30719
rect 7156 30688 8401 30716
rect 7156 30676 7162 30688
rect 8389 30685 8401 30688
rect 8435 30685 8447 30719
rect 9232 30716 9260 30892
rect 9401 30889 9413 30892
rect 9447 30889 9459 30923
rect 9401 30883 9459 30889
rect 10781 30923 10839 30929
rect 10781 30889 10793 30923
rect 10827 30920 10839 30923
rect 11054 30920 11060 30932
rect 10827 30892 11060 30920
rect 10827 30889 10839 30892
rect 10781 30883 10839 30889
rect 11054 30880 11060 30892
rect 11112 30880 11118 30932
rect 9306 30812 9312 30864
rect 9364 30852 9370 30864
rect 9861 30855 9919 30861
rect 9861 30852 9873 30855
rect 9364 30824 9873 30852
rect 9364 30812 9370 30824
rect 9861 30821 9873 30824
rect 9907 30821 9919 30855
rect 11422 30852 11428 30864
rect 11383 30824 11428 30852
rect 9861 30815 9919 30821
rect 11422 30812 11428 30824
rect 11480 30812 11486 30864
rect 9769 30719 9827 30725
rect 9769 30716 9781 30719
rect 9232 30688 9781 30716
rect 8389 30679 8447 30685
rect 9769 30685 9781 30688
rect 9815 30685 9827 30719
rect 9769 30679 9827 30685
rect 10045 30719 10103 30725
rect 10045 30685 10057 30719
rect 10091 30685 10103 30719
rect 11330 30716 11336 30728
rect 11291 30688 11336 30716
rect 10045 30679 10103 30685
rect 8404 30648 8432 30679
rect 10060 30648 10088 30679
rect 11330 30676 11336 30688
rect 11388 30676 11394 30728
rect 11977 30719 12035 30725
rect 11977 30685 11989 30719
rect 12023 30716 12035 30719
rect 12158 30716 12164 30728
rect 12023 30688 12164 30716
rect 12023 30685 12035 30688
rect 11977 30679 12035 30685
rect 12158 30676 12164 30688
rect 12216 30676 12222 30728
rect 8404 30620 10088 30648
rect 6914 30580 6920 30592
rect 6875 30552 6920 30580
rect 6914 30540 6920 30552
rect 6972 30540 6978 30592
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 8478 30336 8484 30388
rect 8536 30376 8542 30388
rect 8987 30379 9045 30385
rect 8987 30376 8999 30379
rect 8536 30348 8999 30376
rect 8536 30336 8542 30348
rect 8987 30345 8999 30348
rect 9033 30345 9045 30379
rect 8987 30339 9045 30345
rect 10781 30379 10839 30385
rect 10781 30345 10793 30379
rect 10827 30376 10839 30379
rect 11333 30379 11391 30385
rect 11333 30376 11345 30379
rect 10827 30348 11345 30376
rect 10827 30345 10839 30348
rect 10781 30339 10839 30345
rect 11333 30345 11345 30348
rect 11379 30376 11391 30379
rect 11422 30376 11428 30388
rect 11379 30348 11428 30376
rect 11379 30345 11391 30348
rect 11333 30339 11391 30345
rect 11422 30336 11428 30348
rect 11480 30336 11486 30388
rect 8757 30311 8815 30317
rect 8757 30277 8769 30311
rect 8803 30308 8815 30311
rect 12158 30308 12164 30320
rect 8803 30280 12164 30308
rect 8803 30277 8815 30280
rect 8757 30271 8815 30277
rect 7466 30172 7472 30184
rect 7427 30144 7472 30172
rect 7466 30132 7472 30144
rect 7524 30132 7530 30184
rect 8931 30181 8959 30280
rect 12158 30268 12164 30280
rect 12216 30268 12222 30320
rect 11330 30200 11336 30252
rect 11388 30240 11394 30252
rect 11609 30243 11667 30249
rect 11609 30240 11621 30243
rect 11388 30212 11621 30240
rect 11388 30200 11394 30212
rect 11609 30209 11621 30212
rect 11655 30209 11667 30243
rect 11609 30203 11667 30209
rect 7745 30175 7803 30181
rect 7745 30141 7757 30175
rect 7791 30141 7803 30175
rect 7745 30135 7803 30141
rect 8916 30175 8974 30181
rect 8916 30141 8928 30175
rect 8962 30141 8974 30175
rect 8916 30135 8974 30141
rect 9861 30175 9919 30181
rect 9861 30141 9873 30175
rect 9907 30172 9919 30175
rect 9950 30172 9956 30184
rect 9907 30144 9956 30172
rect 9907 30141 9919 30144
rect 9861 30135 9919 30141
rect 7760 30104 7788 30135
rect 9950 30132 9956 30144
rect 10008 30132 10014 30184
rect 7116 30076 7788 30104
rect 6638 29996 6644 30048
rect 6696 30036 6702 30048
rect 7116 30045 7144 30076
rect 7101 30039 7159 30045
rect 7101 30036 7113 30039
rect 6696 30008 7113 30036
rect 6696 29996 6702 30008
rect 7101 30005 7113 30008
rect 7147 30005 7159 30039
rect 7558 30036 7564 30048
rect 7519 30008 7564 30036
rect 7101 29999 7159 30005
rect 7558 29996 7564 30008
rect 7616 29996 7622 30048
rect 8294 30036 8300 30048
rect 8255 30008 8300 30036
rect 8294 29996 8300 30008
rect 8352 29996 8358 30048
rect 9306 30036 9312 30048
rect 9267 30008 9312 30036
rect 9306 29996 9312 30008
rect 9364 29996 9370 30048
rect 9769 30039 9827 30045
rect 9769 30005 9781 30039
rect 9815 30036 9827 30039
rect 10226 30036 10232 30048
rect 9815 30008 10232 30036
rect 9815 30005 9827 30008
rect 9769 29999 9827 30005
rect 10226 29996 10232 30008
rect 10284 29996 10290 30048
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 7466 29832 7472 29844
rect 7427 29804 7472 29832
rect 7466 29792 7472 29804
rect 7524 29792 7530 29844
rect 7929 29835 7987 29841
rect 7929 29801 7941 29835
rect 7975 29832 7987 29835
rect 8018 29832 8024 29844
rect 7975 29804 8024 29832
rect 7975 29801 7987 29804
rect 7929 29795 7987 29801
rect 8018 29792 8024 29804
rect 8076 29792 8082 29844
rect 10962 29832 10968 29844
rect 10923 29804 10968 29832
rect 10962 29792 10968 29804
rect 11020 29792 11026 29844
rect 10226 29724 10232 29776
rect 10284 29764 10290 29776
rect 10366 29767 10424 29773
rect 10366 29764 10378 29767
rect 10284 29736 10378 29764
rect 10284 29724 10290 29736
rect 10366 29733 10378 29736
rect 10412 29733 10424 29767
rect 11974 29764 11980 29776
rect 11935 29736 11980 29764
rect 10366 29727 10424 29733
rect 11974 29724 11980 29736
rect 12032 29724 12038 29776
rect 6549 29699 6607 29705
rect 6549 29665 6561 29699
rect 6595 29665 6607 29699
rect 6549 29659 6607 29665
rect 6564 29628 6592 29659
rect 6638 29656 6644 29708
rect 6696 29696 6702 29708
rect 6917 29699 6975 29705
rect 6917 29696 6929 29699
rect 6696 29668 6929 29696
rect 6696 29656 6702 29668
rect 6917 29665 6929 29668
rect 6963 29665 6975 29699
rect 8018 29696 8024 29708
rect 7979 29668 8024 29696
rect 6917 29659 6975 29665
rect 8018 29656 8024 29668
rect 8076 29656 8082 29708
rect 8573 29699 8631 29705
rect 8573 29665 8585 29699
rect 8619 29696 8631 29699
rect 8662 29696 8668 29708
rect 8619 29668 8668 29696
rect 8619 29665 8631 29668
rect 8573 29659 8631 29665
rect 8662 29656 8668 29668
rect 8720 29656 8726 29708
rect 6730 29628 6736 29640
rect 6564 29600 6736 29628
rect 6730 29588 6736 29600
rect 6788 29588 6794 29640
rect 7190 29628 7196 29640
rect 7151 29600 7196 29628
rect 7190 29588 7196 29600
rect 7248 29588 7254 29640
rect 8757 29631 8815 29637
rect 8757 29597 8769 29631
rect 8803 29628 8815 29631
rect 8846 29628 8852 29640
rect 8803 29600 8852 29628
rect 8803 29597 8815 29600
rect 8757 29591 8815 29597
rect 8846 29588 8852 29600
rect 8904 29628 8910 29640
rect 9125 29631 9183 29637
rect 9125 29628 9137 29631
rect 8904 29600 9137 29628
rect 8904 29588 8910 29600
rect 9125 29597 9137 29600
rect 9171 29597 9183 29631
rect 9125 29591 9183 29597
rect 10045 29631 10103 29637
rect 10045 29597 10057 29631
rect 10091 29628 10103 29631
rect 10594 29628 10600 29640
rect 10091 29600 10600 29628
rect 10091 29597 10103 29600
rect 10045 29591 10103 29597
rect 10594 29588 10600 29600
rect 10652 29588 10658 29640
rect 11882 29628 11888 29640
rect 11843 29600 11888 29628
rect 11882 29588 11888 29600
rect 11940 29588 11946 29640
rect 12158 29628 12164 29640
rect 12119 29600 12164 29628
rect 12158 29588 12164 29600
rect 12216 29588 12222 29640
rect 5261 29495 5319 29501
rect 5261 29461 5273 29495
rect 5307 29492 5319 29495
rect 5626 29492 5632 29504
rect 5307 29464 5632 29492
rect 5307 29461 5319 29464
rect 5261 29455 5319 29461
rect 5626 29452 5632 29464
rect 5684 29452 5690 29504
rect 9950 29492 9956 29504
rect 9911 29464 9956 29492
rect 9950 29452 9956 29464
rect 10008 29452 10014 29504
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 5074 29248 5080 29300
rect 5132 29288 5138 29300
rect 5902 29288 5908 29300
rect 5132 29260 5908 29288
rect 5132 29248 5138 29260
rect 5902 29248 5908 29260
rect 5960 29288 5966 29300
rect 8110 29288 8116 29300
rect 5960 29260 8116 29288
rect 5960 29248 5966 29260
rect 8110 29248 8116 29260
rect 8168 29248 8174 29300
rect 8294 29288 8300 29300
rect 8255 29260 8300 29288
rect 8294 29248 8300 29260
rect 8352 29248 8358 29300
rect 8662 29288 8668 29300
rect 8623 29260 8668 29288
rect 8662 29248 8668 29260
rect 8720 29248 8726 29300
rect 10226 29288 10232 29300
rect 9646 29260 10232 29288
rect 4522 29180 4528 29232
rect 4580 29220 4586 29232
rect 7006 29220 7012 29232
rect 4580 29192 7012 29220
rect 4580 29180 4586 29192
rect 7006 29180 7012 29192
rect 7064 29220 7070 29232
rect 8386 29220 8392 29232
rect 7064 29192 8392 29220
rect 7064 29180 7070 29192
rect 8386 29180 8392 29192
rect 8444 29180 8450 29232
rect 5077 29155 5135 29161
rect 5077 29121 5089 29155
rect 5123 29152 5135 29155
rect 5258 29152 5264 29164
rect 5123 29124 5264 29152
rect 5123 29121 5135 29124
rect 5077 29115 5135 29121
rect 5258 29112 5264 29124
rect 5316 29112 5322 29164
rect 5905 29155 5963 29161
rect 5905 29121 5917 29155
rect 5951 29152 5963 29155
rect 7098 29152 7104 29164
rect 5951 29124 7104 29152
rect 5951 29121 5963 29124
rect 5905 29115 5963 29121
rect 7098 29112 7104 29124
rect 7156 29112 7162 29164
rect 7190 29112 7196 29164
rect 7248 29152 7254 29164
rect 7377 29155 7435 29161
rect 7377 29152 7389 29155
rect 7248 29124 7389 29152
rect 7248 29112 7254 29124
rect 7377 29121 7389 29124
rect 7423 29121 7435 29155
rect 7377 29115 7435 29121
rect 8846 29112 8852 29164
rect 8904 29152 8910 29164
rect 9125 29155 9183 29161
rect 9125 29152 9137 29155
rect 8904 29124 9137 29152
rect 8904 29112 8910 29124
rect 9125 29121 9137 29124
rect 9171 29121 9183 29155
rect 9125 29115 9183 29121
rect 7282 29084 7288 29096
rect 7243 29056 7288 29084
rect 7282 29044 7288 29056
rect 7340 29084 7346 29096
rect 7926 29084 7932 29096
rect 7340 29056 7932 29084
rect 7340 29044 7346 29056
rect 5353 29019 5411 29025
rect 5353 28985 5365 29019
rect 5399 29016 5411 29019
rect 5626 29016 5632 29028
rect 5399 28988 5632 29016
rect 5399 28985 5411 28988
rect 5353 28979 5411 28985
rect 5626 28976 5632 28988
rect 5684 28976 5690 29028
rect 7754 29025 7782 29056
rect 7926 29044 7932 29056
rect 7984 29084 7990 29096
rect 8294 29084 8300 29096
rect 7984 29056 8300 29084
rect 7984 29044 7990 29056
rect 8294 29044 8300 29056
rect 8352 29084 8358 29096
rect 8941 29087 8999 29093
rect 8941 29084 8953 29087
rect 8352 29056 8953 29084
rect 8352 29044 8358 29056
rect 8941 29053 8953 29056
rect 8987 29084 8999 29087
rect 9646 29084 9674 29260
rect 10226 29248 10232 29260
rect 10284 29288 10290 29300
rect 10321 29291 10379 29297
rect 10321 29288 10333 29291
rect 10284 29260 10333 29288
rect 10284 29248 10290 29260
rect 10321 29257 10333 29260
rect 10367 29257 10379 29291
rect 11882 29288 11888 29300
rect 11843 29260 11888 29288
rect 10321 29251 10379 29257
rect 11882 29248 11888 29260
rect 11940 29248 11946 29300
rect 10873 29155 10931 29161
rect 10873 29121 10885 29155
rect 10919 29152 10931 29155
rect 11900 29152 11928 29248
rect 10919 29124 11928 29152
rect 10919 29121 10931 29124
rect 10873 29115 10931 29121
rect 8987 29056 9674 29084
rect 10045 29087 10103 29093
rect 8987 29053 8999 29056
rect 8941 29047 8999 29053
rect 9502 29025 9530 29056
rect 10045 29053 10057 29087
rect 10091 29084 10103 29087
rect 11974 29084 11980 29096
rect 10091 29056 11980 29084
rect 10091 29053 10103 29056
rect 10045 29047 10103 29053
rect 11974 29044 11980 29056
rect 12032 29084 12038 29096
rect 12161 29087 12219 29093
rect 12161 29084 12173 29087
rect 12032 29056 12173 29084
rect 12032 29044 12038 29056
rect 12161 29053 12173 29056
rect 12207 29053 12219 29087
rect 12161 29047 12219 29053
rect 7739 29019 7797 29025
rect 7739 29016 7751 29019
rect 7717 28988 7751 29016
rect 7739 28985 7751 28988
rect 7785 28985 7797 29019
rect 9487 29019 9545 29025
rect 9487 29016 9499 29019
rect 9465 28988 9499 29016
rect 7739 28979 7797 28985
rect 9487 28985 9499 28988
rect 9533 28985 9545 29019
rect 9487 28979 9545 28985
rect 6549 28951 6607 28957
rect 6549 28917 6561 28951
rect 6595 28948 6607 28951
rect 6638 28948 6644 28960
rect 6595 28920 6644 28948
rect 6595 28917 6607 28920
rect 6549 28911 6607 28917
rect 6638 28908 6644 28920
rect 6696 28908 6702 28960
rect 10594 28908 10600 28960
rect 10652 28948 10658 28960
rect 10689 28951 10747 28957
rect 10689 28948 10701 28951
rect 10652 28920 10701 28948
rect 10652 28908 10658 28920
rect 10689 28917 10701 28920
rect 10735 28917 10747 28951
rect 10689 28911 10747 28917
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 7190 28704 7196 28756
rect 7248 28744 7254 28756
rect 7469 28747 7527 28753
rect 7469 28744 7481 28747
rect 7248 28716 7481 28744
rect 7248 28704 7254 28716
rect 7469 28713 7481 28716
rect 7515 28713 7527 28747
rect 7469 28707 7527 28713
rect 7926 28704 7932 28756
rect 7984 28744 7990 28756
rect 8021 28747 8079 28753
rect 8021 28744 8033 28747
rect 7984 28716 8033 28744
rect 7984 28704 7990 28716
rect 8021 28713 8033 28716
rect 8067 28713 8079 28747
rect 8021 28707 8079 28713
rect 8573 28747 8631 28753
rect 8573 28713 8585 28747
rect 8619 28744 8631 28747
rect 9306 28744 9312 28756
rect 8619 28716 9312 28744
rect 8619 28713 8631 28716
rect 8573 28707 8631 28713
rect 9306 28704 9312 28716
rect 9364 28704 9370 28756
rect 9950 28744 9956 28756
rect 9911 28716 9956 28744
rect 9950 28704 9956 28716
rect 10008 28704 10014 28756
rect 11425 28747 11483 28753
rect 11425 28744 11437 28747
rect 10152 28716 11437 28744
rect 8662 28636 8668 28688
rect 8720 28676 8726 28688
rect 10152 28676 10180 28716
rect 11425 28713 11437 28716
rect 11471 28713 11483 28747
rect 11425 28707 11483 28713
rect 8720 28648 10180 28676
rect 8720 28636 8726 28648
rect 4801 28611 4859 28617
rect 4801 28577 4813 28611
rect 4847 28608 4859 28611
rect 4890 28608 4896 28620
rect 4847 28580 4896 28608
rect 4847 28577 4859 28580
rect 4801 28571 4859 28577
rect 4890 28568 4896 28580
rect 4948 28568 4954 28620
rect 6178 28608 6184 28620
rect 6139 28580 6184 28608
rect 6178 28568 6184 28580
rect 6236 28568 6242 28620
rect 6638 28608 6644 28620
rect 6551 28580 6644 28608
rect 6638 28568 6644 28580
rect 6696 28608 6702 28620
rect 6696 28580 7230 28608
rect 6696 28568 6702 28580
rect 6822 28540 6828 28552
rect 6783 28512 6828 28540
rect 6822 28500 6828 28512
rect 6880 28500 6886 28552
rect 7202 28540 7230 28580
rect 7558 28568 7564 28620
rect 7616 28608 7622 28620
rect 7653 28611 7711 28617
rect 7653 28608 7665 28611
rect 7616 28580 7665 28608
rect 7616 28568 7622 28580
rect 7653 28577 7665 28580
rect 7699 28577 7711 28611
rect 9674 28608 9680 28620
rect 9635 28580 9680 28608
rect 7653 28571 7711 28577
rect 9674 28568 9680 28580
rect 9732 28568 9738 28620
rect 10152 28617 10180 28648
rect 10137 28611 10195 28617
rect 10137 28577 10149 28611
rect 10183 28577 10195 28611
rect 10137 28571 10195 28577
rect 10962 28568 10968 28620
rect 11020 28608 11026 28620
rect 11241 28611 11299 28617
rect 11241 28608 11253 28611
rect 11020 28580 11253 28608
rect 11020 28568 11026 28580
rect 11241 28577 11253 28580
rect 11287 28577 11299 28611
rect 11241 28571 11299 28577
rect 11054 28540 11060 28552
rect 7202 28512 11060 28540
rect 11054 28500 11060 28512
rect 11112 28500 11118 28552
rect 8018 28432 8024 28484
rect 8076 28472 8082 28484
rect 8386 28472 8392 28484
rect 8076 28444 8392 28472
rect 8076 28432 8082 28444
rect 8386 28432 8392 28444
rect 8444 28472 8450 28484
rect 8849 28475 8907 28481
rect 8849 28472 8861 28475
rect 8444 28444 8861 28472
rect 8444 28432 8450 28444
rect 8849 28441 8861 28444
rect 8895 28441 8907 28475
rect 8849 28435 8907 28441
rect 4798 28364 4804 28416
rect 4856 28404 4862 28416
rect 4939 28407 4997 28413
rect 4939 28404 4951 28407
rect 4856 28376 4951 28404
rect 4856 28364 4862 28376
rect 4939 28373 4951 28376
rect 4985 28373 4997 28407
rect 5258 28404 5264 28416
rect 5219 28376 5264 28404
rect 4939 28367 4997 28373
rect 5258 28364 5264 28376
rect 5316 28364 5322 28416
rect 5350 28364 5356 28416
rect 5408 28404 5414 28416
rect 5629 28407 5687 28413
rect 5629 28404 5641 28407
rect 5408 28376 5641 28404
rect 5408 28364 5414 28376
rect 5629 28373 5641 28376
rect 5675 28373 5687 28407
rect 5629 28367 5687 28373
rect 6730 28364 6736 28416
rect 6788 28404 6794 28416
rect 7193 28407 7251 28413
rect 7193 28404 7205 28407
rect 6788 28376 7205 28404
rect 6788 28364 6794 28376
rect 7193 28373 7205 28376
rect 7239 28404 7251 28407
rect 9582 28404 9588 28416
rect 7239 28376 9588 28404
rect 7239 28373 7251 28376
rect 7193 28367 7251 28373
rect 9582 28364 9588 28376
rect 9640 28364 9646 28416
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 4430 28200 4436 28212
rect 4391 28172 4436 28200
rect 4430 28160 4436 28172
rect 4488 28160 4494 28212
rect 4890 28200 4896 28212
rect 4851 28172 4896 28200
rect 4890 28160 4896 28172
rect 4948 28160 4954 28212
rect 6181 28203 6239 28209
rect 6181 28169 6193 28203
rect 6227 28200 6239 28203
rect 6638 28200 6644 28212
rect 6227 28172 6644 28200
rect 6227 28169 6239 28172
rect 6181 28163 6239 28169
rect 6638 28160 6644 28172
rect 6696 28160 6702 28212
rect 7558 28160 7564 28212
rect 7616 28200 7622 28212
rect 8389 28203 8447 28209
rect 8389 28200 8401 28203
rect 7616 28172 8401 28200
rect 7616 28160 7622 28172
rect 8389 28169 8401 28172
rect 8435 28169 8447 28203
rect 8389 28163 8447 28169
rect 8662 28160 8668 28212
rect 8720 28200 8726 28212
rect 9125 28203 9183 28209
rect 9125 28200 9137 28203
rect 8720 28172 9137 28200
rect 8720 28160 8726 28172
rect 9125 28169 9137 28172
rect 9171 28200 9183 28203
rect 10321 28203 10379 28209
rect 10321 28200 10333 28203
rect 9171 28172 10333 28200
rect 9171 28169 9183 28172
rect 9125 28163 9183 28169
rect 5626 28092 5632 28144
rect 5684 28132 5690 28144
rect 7745 28135 7803 28141
rect 7745 28132 7757 28135
rect 5684 28104 7757 28132
rect 5684 28092 5690 28104
rect 7745 28101 7757 28104
rect 7791 28101 7803 28135
rect 7745 28095 7803 28101
rect 7837 28135 7895 28141
rect 7837 28101 7849 28135
rect 7883 28132 7895 28135
rect 8113 28135 8171 28141
rect 8113 28132 8125 28135
rect 7883 28104 8125 28132
rect 7883 28101 7895 28104
rect 7837 28095 7895 28101
rect 8113 28101 8125 28104
rect 8159 28132 8171 28135
rect 8294 28132 8300 28144
rect 8159 28104 8300 28132
rect 8159 28101 8171 28104
rect 8113 28095 8171 28101
rect 8294 28092 8300 28104
rect 8352 28092 8358 28144
rect 5077 28067 5135 28073
rect 5077 28033 5089 28067
rect 5123 28064 5135 28067
rect 5350 28064 5356 28076
rect 5123 28036 5356 28064
rect 5123 28033 5135 28036
rect 5077 28027 5135 28033
rect 5350 28024 5356 28036
rect 5408 28024 5414 28076
rect 6822 28064 6828 28076
rect 6783 28036 6828 28064
rect 6822 28024 6828 28036
rect 6880 28024 6886 28076
rect 7466 28024 7472 28076
rect 7524 28064 7530 28076
rect 8757 28067 8815 28073
rect 8757 28064 8769 28067
rect 7524 28036 8769 28064
rect 7524 28024 7530 28036
rect 8757 28033 8769 28036
rect 8803 28064 8815 28067
rect 9674 28064 9680 28076
rect 8803 28036 9680 28064
rect 8803 28033 8815 28036
rect 8757 28027 8815 28033
rect 9674 28024 9680 28036
rect 9732 28024 9738 28076
rect 3510 27956 3516 28008
rect 3568 27996 3574 28008
rect 4008 27999 4066 28005
rect 4008 27996 4020 27999
rect 3568 27968 4020 27996
rect 3568 27956 3574 27968
rect 4008 27965 4020 27968
rect 4054 27996 4066 27999
rect 4430 27996 4436 28008
rect 4054 27968 4436 27996
rect 4054 27965 4066 27968
rect 4008 27959 4066 27965
rect 4430 27956 4436 27968
rect 4488 27956 4494 28008
rect 9582 27996 9588 28008
rect 9543 27968 9588 27996
rect 9582 27956 9588 27968
rect 9640 27956 9646 28008
rect 9784 28005 9812 28172
rect 10321 28169 10333 28172
rect 10367 28169 10379 28203
rect 11054 28200 11060 28212
rect 11015 28172 11060 28200
rect 10321 28163 10379 28169
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 10045 28067 10103 28073
rect 10045 28033 10057 28067
rect 10091 28064 10103 28067
rect 10594 28064 10600 28076
rect 10091 28036 10600 28064
rect 10091 28033 10103 28036
rect 10045 28027 10103 28033
rect 10594 28024 10600 28036
rect 10652 28024 10658 28076
rect 9769 27999 9827 28005
rect 9769 27965 9781 27999
rect 9815 27965 9827 27999
rect 9769 27959 9827 27965
rect 10873 27999 10931 28005
rect 10873 27965 10885 27999
rect 10919 27996 10931 27999
rect 11701 27999 11759 28005
rect 11701 27996 11713 27999
rect 10919 27968 11713 27996
rect 10919 27965 10931 27968
rect 10873 27959 10931 27965
rect 11701 27965 11713 27968
rect 11747 27965 11759 27999
rect 11701 27959 11759 27965
rect 3050 27888 3056 27940
rect 3108 27928 3114 27940
rect 4890 27928 4896 27940
rect 3108 27900 4896 27928
rect 3108 27888 3114 27900
rect 4890 27888 4896 27900
rect 4948 27888 4954 27940
rect 5169 27931 5227 27937
rect 5169 27897 5181 27931
rect 5215 27928 5227 27931
rect 5258 27928 5264 27940
rect 5215 27900 5264 27928
rect 5215 27897 5227 27900
rect 5169 27891 5227 27897
rect 5258 27888 5264 27900
rect 5316 27888 5322 27940
rect 5721 27931 5779 27937
rect 5721 27897 5733 27931
rect 5767 27928 5779 27931
rect 5902 27928 5908 27940
rect 5767 27900 5908 27928
rect 5767 27897 5779 27900
rect 5721 27891 5779 27897
rect 5902 27888 5908 27900
rect 5960 27888 5966 27940
rect 6641 27931 6699 27937
rect 6641 27897 6653 27931
rect 6687 27928 6699 27931
rect 7187 27931 7245 27937
rect 7187 27928 7199 27931
rect 6687 27900 7199 27928
rect 6687 27897 6699 27900
rect 6641 27891 6699 27897
rect 7187 27897 7199 27900
rect 7233 27928 7245 27931
rect 7837 27931 7895 27937
rect 7837 27928 7849 27931
rect 7233 27900 7849 27928
rect 7233 27897 7245 27900
rect 7187 27891 7245 27897
rect 7837 27897 7849 27900
rect 7883 27897 7895 27931
rect 7837 27891 7895 27897
rect 8570 27888 8576 27940
rect 8628 27928 8634 27940
rect 10888 27928 10916 27959
rect 8628 27900 10916 27928
rect 8628 27888 8634 27900
rect 10962 27888 10968 27940
rect 11020 27928 11026 27940
rect 11333 27931 11391 27937
rect 11333 27928 11345 27931
rect 11020 27900 11345 27928
rect 11020 27888 11026 27900
rect 11333 27897 11345 27900
rect 11379 27897 11391 27931
rect 11333 27891 11391 27897
rect 4111 27863 4169 27869
rect 4111 27829 4123 27863
rect 4157 27860 4169 27863
rect 5994 27860 6000 27872
rect 4157 27832 6000 27860
rect 4157 27829 4169 27832
rect 4111 27823 4169 27829
rect 5994 27820 6000 27832
rect 6052 27820 6058 27872
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 4798 27656 4804 27668
rect 4759 27628 4804 27656
rect 4798 27616 4804 27628
rect 4856 27616 4862 27668
rect 5169 27659 5227 27665
rect 5169 27625 5181 27659
rect 5215 27656 5227 27659
rect 5258 27656 5264 27668
rect 5215 27628 5264 27656
rect 5215 27625 5227 27628
rect 5169 27619 5227 27625
rect 5258 27616 5264 27628
rect 5316 27616 5322 27668
rect 6733 27659 6791 27665
rect 6733 27625 6745 27659
rect 6779 27656 6791 27659
rect 6822 27656 6828 27668
rect 6779 27628 6828 27656
rect 6779 27625 6791 27628
rect 6733 27619 6791 27625
rect 6822 27616 6828 27628
rect 6880 27616 6886 27668
rect 4387 27591 4445 27597
rect 4387 27557 4399 27591
rect 4433 27588 4445 27591
rect 5350 27588 5356 27600
rect 4433 27560 5356 27588
rect 4433 27557 4445 27560
rect 4387 27551 4445 27557
rect 5350 27548 5356 27560
rect 5408 27548 5414 27600
rect 5445 27591 5503 27597
rect 5445 27557 5457 27591
rect 5491 27588 5503 27591
rect 5626 27588 5632 27600
rect 5491 27560 5632 27588
rect 5491 27557 5503 27560
rect 5445 27551 5503 27557
rect 5626 27548 5632 27560
rect 5684 27588 5690 27600
rect 6270 27588 6276 27600
rect 5684 27560 6276 27588
rect 5684 27548 5690 27560
rect 6270 27548 6276 27560
rect 6328 27588 6334 27600
rect 7009 27591 7067 27597
rect 7009 27588 7021 27591
rect 6328 27560 7021 27588
rect 6328 27548 6334 27560
rect 7009 27557 7021 27560
rect 7055 27557 7067 27591
rect 9858 27588 9864 27600
rect 9819 27560 9864 27588
rect 7009 27551 7067 27557
rect 9858 27548 9864 27560
rect 9916 27548 9922 27600
rect 11425 27591 11483 27597
rect 11425 27557 11437 27591
rect 11471 27588 11483 27591
rect 11974 27588 11980 27600
rect 11471 27560 11980 27588
rect 11471 27557 11483 27560
rect 11425 27551 11483 27557
rect 11974 27548 11980 27560
rect 12032 27548 12038 27600
rect 4300 27523 4358 27529
rect 4300 27489 4312 27523
rect 4346 27520 4358 27523
rect 4522 27520 4528 27532
rect 4346 27492 4528 27520
rect 4346 27489 4358 27492
rect 4300 27483 4358 27489
rect 4522 27480 4528 27492
rect 4580 27480 4586 27532
rect 8202 27480 8208 27532
rect 8260 27520 8266 27532
rect 8456 27523 8514 27529
rect 8456 27520 8468 27523
rect 8260 27492 8468 27520
rect 8260 27480 8266 27492
rect 8456 27489 8468 27492
rect 8502 27520 8514 27523
rect 8754 27520 8760 27532
rect 8502 27492 8760 27520
rect 8502 27489 8514 27492
rect 8456 27483 8514 27489
rect 8754 27480 8760 27492
rect 8812 27480 8818 27532
rect 12434 27480 12440 27532
rect 12492 27520 12498 27532
rect 12872 27523 12930 27529
rect 12872 27520 12884 27523
rect 12492 27492 12884 27520
rect 12492 27480 12498 27492
rect 12872 27489 12884 27492
rect 12918 27520 12930 27523
rect 13262 27520 13268 27532
rect 12918 27492 13268 27520
rect 12918 27489 12930 27492
rect 12872 27483 12930 27489
rect 13262 27480 13268 27492
rect 13320 27480 13326 27532
rect 5353 27455 5411 27461
rect 5353 27421 5365 27455
rect 5399 27452 5411 27455
rect 5718 27452 5724 27464
rect 5399 27424 5724 27452
rect 5399 27421 5411 27424
rect 5353 27415 5411 27421
rect 5718 27412 5724 27424
rect 5776 27412 5782 27464
rect 6917 27455 6975 27461
rect 6917 27421 6929 27455
rect 6963 27452 6975 27455
rect 7834 27452 7840 27464
rect 6963 27424 7840 27452
rect 6963 27421 6975 27424
rect 6917 27415 6975 27421
rect 7834 27412 7840 27424
rect 7892 27412 7898 27464
rect 9398 27412 9404 27464
rect 9456 27452 9462 27464
rect 9769 27455 9827 27461
rect 9769 27452 9781 27455
rect 9456 27424 9781 27452
rect 9456 27412 9462 27424
rect 9769 27421 9781 27424
rect 9815 27421 9827 27455
rect 9769 27415 9827 27421
rect 10413 27455 10471 27461
rect 10413 27421 10425 27455
rect 10459 27452 10471 27455
rect 11146 27452 11152 27464
rect 10459 27424 11152 27452
rect 10459 27421 10471 27424
rect 10413 27415 10471 27421
rect 11146 27412 11152 27424
rect 11204 27452 11210 27464
rect 11333 27455 11391 27461
rect 11333 27452 11345 27455
rect 11204 27424 11345 27452
rect 11204 27412 11210 27424
rect 11333 27421 11345 27424
rect 11379 27421 11391 27455
rect 11333 27415 11391 27421
rect 11514 27412 11520 27464
rect 11572 27452 11578 27464
rect 11609 27455 11667 27461
rect 11609 27452 11621 27455
rect 11572 27424 11621 27452
rect 11572 27412 11578 27424
rect 11609 27421 11621 27424
rect 11655 27421 11667 27455
rect 11609 27415 11667 27421
rect 5902 27384 5908 27396
rect 5863 27356 5908 27384
rect 5902 27344 5908 27356
rect 5960 27344 5966 27396
rect 7466 27384 7472 27396
rect 7427 27356 7472 27384
rect 7466 27344 7472 27356
rect 7524 27344 7530 27396
rect 6178 27276 6184 27328
rect 6236 27316 6242 27328
rect 6365 27319 6423 27325
rect 6365 27316 6377 27319
rect 6236 27288 6377 27316
rect 6236 27276 6242 27288
rect 6365 27285 6377 27288
rect 6411 27316 6423 27319
rect 6638 27316 6644 27328
rect 6411 27288 6644 27316
rect 6411 27285 6423 27288
rect 6365 27279 6423 27285
rect 6638 27276 6644 27288
rect 6696 27316 6702 27328
rect 8386 27316 8392 27328
rect 6696 27288 8392 27316
rect 6696 27276 6702 27288
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 8527 27319 8585 27325
rect 8527 27285 8539 27319
rect 8573 27316 8585 27319
rect 8846 27316 8852 27328
rect 8573 27288 8852 27316
rect 8573 27285 8585 27288
rect 8527 27279 8585 27285
rect 8846 27276 8852 27288
rect 8904 27276 8910 27328
rect 9401 27319 9459 27325
rect 9401 27285 9413 27319
rect 9447 27316 9459 27319
rect 9582 27316 9588 27328
rect 9447 27288 9588 27316
rect 9447 27285 9459 27288
rect 9401 27279 9459 27285
rect 9582 27276 9588 27288
rect 9640 27276 9646 27328
rect 12526 27276 12532 27328
rect 12584 27316 12590 27328
rect 12943 27319 13001 27325
rect 12943 27316 12955 27319
rect 12584 27288 12955 27316
rect 12584 27276 12590 27288
rect 12943 27285 12955 27288
rect 12989 27285 13001 27319
rect 12943 27279 13001 27285
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 3191 27115 3249 27121
rect 3191 27081 3203 27115
rect 3237 27112 3249 27115
rect 5718 27112 5724 27124
rect 3237 27084 5724 27112
rect 3237 27081 3249 27084
rect 3191 27075 3249 27081
rect 5718 27072 5724 27084
rect 5776 27072 5782 27124
rect 6270 27112 6276 27124
rect 6231 27084 6276 27112
rect 6270 27072 6276 27084
rect 6328 27072 6334 27124
rect 7834 27112 7840 27124
rect 7795 27084 7840 27112
rect 7834 27072 7840 27084
rect 7892 27112 7898 27124
rect 8527 27115 8585 27121
rect 8527 27112 8539 27115
rect 7892 27084 8539 27112
rect 7892 27072 7898 27084
rect 8527 27081 8539 27084
rect 8573 27081 8585 27115
rect 8527 27075 8585 27081
rect 13630 27072 13636 27124
rect 13688 27112 13694 27124
rect 13725 27115 13783 27121
rect 13725 27112 13737 27115
rect 13688 27084 13737 27112
rect 13688 27072 13694 27084
rect 13725 27081 13737 27084
rect 13771 27081 13783 27115
rect 13725 27075 13783 27081
rect 4154 27044 4160 27056
rect 3135 27016 4160 27044
rect 3135 26917 3163 27016
rect 4154 27004 4160 27016
rect 4212 27004 4218 27056
rect 4522 27044 4528 27056
rect 4483 27016 4528 27044
rect 4522 27004 4528 27016
rect 4580 27004 4586 27056
rect 7466 27044 7472 27056
rect 5828 27016 7472 27044
rect 4798 26936 4804 26988
rect 4856 26976 4862 26988
rect 5828 26985 5856 27016
rect 7466 27004 7472 27016
rect 7524 27004 7530 27056
rect 10229 27047 10287 27053
rect 10229 27013 10241 27047
rect 10275 27044 10287 27047
rect 11146 27044 11152 27056
rect 10275 27016 11152 27044
rect 10275 27013 10287 27016
rect 10229 27007 10287 27013
rect 11146 27004 11152 27016
rect 11204 27004 11210 27056
rect 5169 26979 5227 26985
rect 5169 26976 5181 26979
rect 4856 26948 5181 26976
rect 4856 26936 4862 26948
rect 5169 26945 5181 26948
rect 5215 26945 5227 26979
rect 5169 26939 5227 26945
rect 5813 26979 5871 26985
rect 5813 26945 5825 26979
rect 5859 26945 5871 26979
rect 5813 26939 5871 26945
rect 5994 26936 6000 26988
rect 6052 26976 6058 26988
rect 6917 26979 6975 26985
rect 6917 26976 6929 26979
rect 6052 26948 6929 26976
rect 6052 26936 6058 26948
rect 6917 26945 6929 26948
rect 6963 26976 6975 26979
rect 7098 26976 7104 26988
rect 6963 26948 7104 26976
rect 6963 26945 6975 26948
rect 6917 26939 6975 26945
rect 7098 26936 7104 26948
rect 7156 26936 7162 26988
rect 9858 26936 9864 26988
rect 9916 26976 9922 26988
rect 10965 26979 11023 26985
rect 10965 26976 10977 26979
rect 9916 26948 10977 26976
rect 9916 26936 9922 26948
rect 10965 26945 10977 26948
rect 11011 26945 11023 26979
rect 10965 26939 11023 26945
rect 3120 26911 3178 26917
rect 3120 26877 3132 26911
rect 3166 26877 3178 26911
rect 3120 26871 3178 26877
rect 3135 26840 3163 26871
rect 3234 26868 3240 26920
rect 3292 26908 3298 26920
rect 4116 26911 4174 26917
rect 4116 26908 4128 26911
rect 3292 26880 4128 26908
rect 3292 26868 3298 26880
rect 4116 26877 4128 26880
rect 4162 26908 4174 26911
rect 4614 26908 4620 26920
rect 4162 26880 4620 26908
rect 4162 26877 4174 26880
rect 4116 26871 4174 26877
rect 4614 26868 4620 26880
rect 4672 26868 4678 26920
rect 6178 26868 6184 26920
rect 6236 26908 6242 26920
rect 6549 26911 6607 26917
rect 6549 26908 6561 26911
rect 6236 26880 6561 26908
rect 6236 26868 6242 26880
rect 6549 26877 6561 26880
rect 6595 26877 6607 26911
rect 6549 26871 6607 26877
rect 4203 26843 4261 26849
rect 3135 26812 3280 26840
rect 3252 26784 3280 26812
rect 4203 26809 4215 26843
rect 4249 26840 4261 26843
rect 4982 26840 4988 26852
rect 4249 26812 4988 26840
rect 4249 26809 4261 26812
rect 4203 26803 4261 26809
rect 4982 26800 4988 26812
rect 5040 26800 5046 26852
rect 5258 26840 5264 26852
rect 5219 26812 5264 26840
rect 5258 26800 5264 26812
rect 5316 26800 5322 26852
rect 3234 26732 3240 26784
rect 3292 26772 3298 26784
rect 3513 26775 3571 26781
rect 3513 26772 3525 26775
rect 3292 26744 3525 26772
rect 3292 26732 3298 26744
rect 3513 26741 3525 26744
rect 3559 26741 3571 26775
rect 3513 26735 3571 26741
rect 4614 26732 4620 26784
rect 4672 26772 4678 26784
rect 4893 26775 4951 26781
rect 4893 26772 4905 26775
rect 4672 26744 4905 26772
rect 4672 26732 4678 26744
rect 4893 26741 4905 26744
rect 4939 26741 4951 26775
rect 6564 26772 6592 26871
rect 8110 26868 8116 26920
rect 8168 26908 8174 26920
rect 8424 26911 8482 26917
rect 8424 26908 8436 26911
rect 8168 26880 8436 26908
rect 8168 26868 8174 26880
rect 8424 26877 8436 26880
rect 8470 26908 8482 26911
rect 9217 26911 9275 26917
rect 9217 26908 9229 26911
rect 8470 26880 9229 26908
rect 8470 26877 8482 26880
rect 8424 26871 8482 26877
rect 9217 26877 9229 26880
rect 9263 26877 9275 26911
rect 9217 26871 9275 26877
rect 11054 26868 11060 26920
rect 11112 26908 11118 26920
rect 11184 26911 11242 26917
rect 11184 26908 11196 26911
rect 11112 26880 11196 26908
rect 11112 26868 11118 26880
rect 11184 26877 11196 26880
rect 11230 26908 11242 26911
rect 11609 26911 11667 26917
rect 11609 26908 11621 26911
rect 11230 26880 11621 26908
rect 11230 26877 11242 26880
rect 11184 26871 11242 26877
rect 11609 26877 11621 26880
rect 11655 26877 11667 26911
rect 11609 26871 11667 26877
rect 12250 26868 12256 26920
rect 12308 26908 12314 26920
rect 12472 26911 12530 26917
rect 12472 26908 12484 26911
rect 12308 26880 12484 26908
rect 12308 26868 12314 26880
rect 12472 26877 12484 26880
rect 12518 26908 12530 26911
rect 12710 26908 12716 26920
rect 12518 26880 12716 26908
rect 12518 26877 12530 26880
rect 12472 26871 12530 26877
rect 12710 26868 12716 26880
rect 12768 26908 12774 26920
rect 12897 26911 12955 26917
rect 12897 26908 12909 26911
rect 12768 26880 12909 26908
rect 12768 26868 12774 26880
rect 12897 26877 12909 26880
rect 12943 26877 12955 26911
rect 12897 26871 12955 26877
rect 13484 26911 13542 26917
rect 13484 26877 13496 26911
rect 13530 26877 13542 26911
rect 13484 26871 13542 26877
rect 7009 26843 7067 26849
rect 7009 26809 7021 26843
rect 7055 26809 7067 26843
rect 7009 26803 7067 26809
rect 7024 26772 7052 26803
rect 9490 26800 9496 26852
rect 9548 26840 9554 26852
rect 9677 26843 9735 26849
rect 9677 26840 9689 26843
rect 9548 26812 9689 26840
rect 9548 26800 9554 26812
rect 9677 26809 9689 26812
rect 9723 26809 9735 26843
rect 9677 26803 9735 26809
rect 9766 26800 9772 26852
rect 9824 26840 9830 26852
rect 10597 26843 10655 26849
rect 10597 26840 10609 26843
rect 9824 26812 10609 26840
rect 9824 26800 9830 26812
rect 10597 26809 10609 26812
rect 10643 26809 10655 26843
rect 10597 26803 10655 26809
rect 11514 26800 11520 26852
rect 11572 26840 11578 26852
rect 13499 26840 13527 26871
rect 13909 26843 13967 26849
rect 13909 26840 13921 26843
rect 11572 26812 13921 26840
rect 11572 26800 11578 26812
rect 13909 26809 13921 26812
rect 13955 26809 13967 26843
rect 13909 26803 13967 26809
rect 6564 26744 7052 26772
rect 4893 26735 4951 26741
rect 8754 26732 8760 26784
rect 8812 26772 8818 26784
rect 8849 26775 8907 26781
rect 8849 26772 8861 26775
rect 8812 26744 8861 26772
rect 8812 26732 8818 26744
rect 8849 26741 8861 26744
rect 8895 26741 8907 26775
rect 8849 26735 8907 26741
rect 11054 26732 11060 26784
rect 11112 26772 11118 26784
rect 11287 26775 11345 26781
rect 11287 26772 11299 26775
rect 11112 26744 11299 26772
rect 11112 26732 11118 26744
rect 11287 26741 11299 26744
rect 11333 26741 11345 26775
rect 11974 26772 11980 26784
rect 11935 26744 11980 26772
rect 11287 26735 11345 26741
rect 11974 26732 11980 26744
rect 12032 26732 12038 26784
rect 12066 26732 12072 26784
rect 12124 26772 12130 26784
rect 12575 26775 12633 26781
rect 12575 26772 12587 26775
rect 12124 26744 12587 26772
rect 12124 26732 12130 26744
rect 12575 26741 12587 26744
rect 12621 26741 12633 26775
rect 13262 26772 13268 26784
rect 13223 26744 13268 26772
rect 12575 26735 12633 26741
rect 13262 26732 13268 26744
rect 13320 26732 13326 26784
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 5261 26571 5319 26577
rect 5261 26537 5273 26571
rect 5307 26568 5319 26571
rect 5626 26568 5632 26580
rect 5307 26540 5632 26568
rect 5307 26537 5319 26540
rect 5261 26531 5319 26537
rect 5626 26528 5632 26540
rect 5684 26528 5690 26580
rect 5718 26528 5724 26580
rect 5776 26568 5782 26580
rect 5905 26571 5963 26577
rect 5905 26568 5917 26571
rect 5776 26540 5917 26568
rect 5776 26528 5782 26540
rect 5905 26537 5917 26540
rect 5951 26537 5963 26571
rect 7098 26568 7104 26580
rect 7059 26540 7104 26568
rect 5905 26531 5963 26537
rect 7098 26528 7104 26540
rect 7156 26528 7162 26580
rect 10042 26528 10048 26580
rect 10100 26568 10106 26580
rect 12897 26571 12955 26577
rect 12897 26568 12909 26571
rect 10100 26540 12909 26568
rect 10100 26528 10106 26540
rect 12897 26537 12909 26540
rect 12943 26537 12955 26571
rect 12897 26531 12955 26537
rect 4154 26460 4160 26512
rect 4212 26500 4218 26512
rect 4662 26503 4720 26509
rect 4662 26500 4674 26503
rect 4212 26472 4674 26500
rect 4212 26460 4218 26472
rect 4662 26469 4674 26472
rect 4708 26469 4720 26503
rect 4662 26463 4720 26469
rect 6178 26460 6184 26512
rect 6236 26500 6242 26512
rect 6273 26503 6331 26509
rect 6273 26500 6285 26503
rect 6236 26472 6285 26500
rect 6236 26460 6242 26472
rect 6273 26469 6285 26472
rect 6319 26469 6331 26503
rect 9858 26500 9864 26512
rect 9819 26472 9864 26500
rect 6273 26463 6331 26469
rect 9858 26460 9864 26472
rect 9916 26460 9922 26512
rect 11425 26503 11483 26509
rect 11425 26469 11437 26503
rect 11471 26500 11483 26503
rect 12618 26500 12624 26512
rect 11471 26472 12624 26500
rect 11471 26469 11483 26472
rect 11425 26463 11483 26469
rect 12618 26460 12624 26472
rect 12676 26460 12682 26512
rect 7834 26432 7840 26444
rect 7795 26404 7840 26432
rect 7834 26392 7840 26404
rect 7892 26392 7898 26444
rect 8294 26432 8300 26444
rect 8255 26404 8300 26432
rect 8294 26392 8300 26404
rect 8352 26392 8358 26444
rect 13078 26432 13084 26444
rect 13039 26404 13084 26432
rect 13078 26392 13084 26404
rect 13136 26392 13142 26444
rect 13265 26435 13323 26441
rect 13265 26401 13277 26435
rect 13311 26401 13323 26435
rect 13265 26395 13323 26401
rect 4341 26367 4399 26373
rect 4341 26333 4353 26367
rect 4387 26364 4399 26367
rect 4798 26364 4804 26376
rect 4387 26336 4804 26364
rect 4387 26333 4399 26336
rect 4341 26327 4399 26333
rect 4798 26324 4804 26336
rect 4856 26324 4862 26376
rect 4982 26324 4988 26376
rect 5040 26364 5046 26376
rect 6181 26367 6239 26373
rect 6181 26364 6193 26367
rect 5040 26336 6193 26364
rect 5040 26324 5046 26336
rect 6181 26333 6193 26336
rect 6227 26364 6239 26367
rect 6454 26364 6460 26376
rect 6227 26336 6460 26364
rect 6227 26333 6239 26336
rect 6181 26327 6239 26333
rect 6454 26324 6460 26336
rect 6512 26324 6518 26376
rect 8386 26364 8392 26376
rect 8347 26336 8392 26364
rect 8386 26324 8392 26336
rect 8444 26324 8450 26376
rect 9769 26367 9827 26373
rect 9769 26333 9781 26367
rect 9815 26364 9827 26367
rect 9950 26364 9956 26376
rect 9815 26336 9956 26364
rect 9815 26333 9827 26336
rect 9769 26327 9827 26333
rect 9950 26324 9956 26336
rect 10008 26364 10014 26376
rect 11054 26364 11060 26376
rect 10008 26336 11060 26364
rect 10008 26324 10014 26336
rect 11054 26324 11060 26336
rect 11112 26324 11118 26376
rect 11333 26367 11391 26373
rect 11333 26333 11345 26367
rect 11379 26364 11391 26367
rect 11698 26364 11704 26376
rect 11379 26336 11704 26364
rect 11379 26333 11391 26336
rect 11333 26327 11391 26333
rect 11698 26324 11704 26336
rect 11756 26364 11762 26376
rect 12066 26364 12072 26376
rect 11756 26336 12072 26364
rect 11756 26324 11762 26336
rect 12066 26324 12072 26336
rect 12124 26324 12130 26376
rect 12250 26324 12256 26376
rect 12308 26364 12314 26376
rect 13280 26364 13308 26395
rect 12308 26336 13308 26364
rect 12308 26324 12314 26336
rect 5350 26256 5356 26308
rect 5408 26296 5414 26308
rect 5902 26296 5908 26308
rect 5408 26268 5908 26296
rect 5408 26256 5414 26268
rect 5902 26256 5908 26268
rect 5960 26296 5966 26308
rect 6733 26299 6791 26305
rect 6733 26296 6745 26299
rect 5960 26268 6745 26296
rect 5960 26256 5966 26268
rect 6733 26265 6745 26268
rect 6779 26265 6791 26299
rect 6733 26259 6791 26265
rect 9125 26299 9183 26305
rect 9125 26265 9137 26299
rect 9171 26296 9183 26299
rect 9398 26296 9404 26308
rect 9171 26268 9404 26296
rect 9171 26265 9183 26268
rect 9125 26259 9183 26265
rect 9398 26256 9404 26268
rect 9456 26256 9462 26308
rect 10321 26299 10379 26305
rect 10321 26265 10333 26299
rect 10367 26296 10379 26299
rect 11238 26296 11244 26308
rect 10367 26268 11244 26296
rect 10367 26265 10379 26268
rect 10321 26259 10379 26265
rect 11238 26256 11244 26268
rect 11296 26296 11302 26308
rect 11885 26299 11943 26305
rect 11885 26296 11897 26299
rect 11296 26268 11897 26296
rect 11296 26256 11302 26268
rect 11885 26265 11897 26268
rect 11931 26265 11943 26299
rect 11885 26259 11943 26265
rect 2866 26188 2872 26240
rect 2924 26228 2930 26240
rect 5534 26228 5540 26240
rect 2924 26200 5540 26228
rect 2924 26188 2930 26200
rect 5534 26188 5540 26200
rect 5592 26228 5598 26240
rect 7190 26228 7196 26240
rect 5592 26200 7196 26228
rect 5592 26188 5598 26200
rect 7190 26188 7196 26200
rect 7248 26188 7254 26240
rect 7561 26231 7619 26237
rect 7561 26197 7573 26231
rect 7607 26228 7619 26231
rect 7650 26228 7656 26240
rect 7607 26200 7656 26228
rect 7607 26197 7619 26200
rect 7561 26191 7619 26197
rect 7650 26188 7656 26200
rect 7708 26188 7714 26240
rect 9490 26228 9496 26240
rect 9451 26200 9496 26228
rect 9490 26188 9496 26200
rect 9548 26188 9554 26240
rect 10686 26228 10692 26240
rect 10647 26200 10692 26228
rect 10686 26188 10692 26200
rect 10744 26188 10750 26240
rect 11146 26228 11152 26240
rect 11107 26200 11152 26228
rect 11146 26188 11152 26200
rect 11204 26188 11210 26240
rect 12529 26231 12587 26237
rect 12529 26197 12541 26231
rect 12575 26228 12587 26231
rect 12618 26228 12624 26240
rect 12575 26200 12624 26228
rect 12575 26197 12587 26200
rect 12529 26191 12587 26197
rect 12618 26188 12624 26200
rect 12676 26188 12682 26240
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 5169 26027 5227 26033
rect 5169 25993 5181 26027
rect 5215 26024 5227 26027
rect 5258 26024 5264 26036
rect 5215 25996 5264 26024
rect 5215 25993 5227 25996
rect 5169 25987 5227 25993
rect 5258 25984 5264 25996
rect 5316 25984 5322 26036
rect 6454 26024 6460 26036
rect 6415 25996 6460 26024
rect 6454 25984 6460 25996
rect 6512 25984 6518 26036
rect 6914 26024 6920 26036
rect 6564 25996 6920 26024
rect 2958 25916 2964 25968
rect 3016 25956 3022 25968
rect 6564 25956 6592 25996
rect 6914 25984 6920 25996
rect 6972 26024 6978 26036
rect 7469 26027 7527 26033
rect 7469 26024 7481 26027
rect 6972 25996 7481 26024
rect 6972 25984 6978 25996
rect 7469 25993 7481 25996
rect 7515 26024 7527 26027
rect 8294 26024 8300 26036
rect 7515 25996 8300 26024
rect 7515 25993 7527 25996
rect 7469 25987 7527 25993
rect 8294 25984 8300 25996
rect 8352 25984 8358 26036
rect 9585 26027 9643 26033
rect 9585 25993 9597 26027
rect 9631 26024 9643 26027
rect 9858 26024 9864 26036
rect 9631 25996 9864 26024
rect 9631 25993 9643 25996
rect 9585 25987 9643 25993
rect 9858 25984 9864 25996
rect 9916 26024 9922 26036
rect 10965 26027 11023 26033
rect 10965 26024 10977 26027
rect 9916 25996 10977 26024
rect 9916 25984 9922 25996
rect 10965 25993 10977 25996
rect 11011 25993 11023 26027
rect 11698 26024 11704 26036
rect 11659 25996 11704 26024
rect 10965 25987 11023 25993
rect 11698 25984 11704 25996
rect 11756 25984 11762 26036
rect 13078 25984 13084 26036
rect 13136 26024 13142 26036
rect 13449 26027 13507 26033
rect 13449 26024 13461 26027
rect 13136 25996 13461 26024
rect 13136 25984 13142 25996
rect 13449 25993 13461 25996
rect 13495 25993 13507 26027
rect 13449 25987 13507 25993
rect 7745 25959 7803 25965
rect 7745 25956 7757 25959
rect 3016 25928 6592 25956
rect 6656 25928 7757 25956
rect 3016 25916 3022 25928
rect 2682 25848 2688 25900
rect 2740 25888 2746 25900
rect 6656 25888 6684 25928
rect 7745 25925 7757 25928
rect 7791 25956 7803 25959
rect 7834 25956 7840 25968
rect 7791 25928 7840 25956
rect 7791 25925 7803 25928
rect 7745 25919 7803 25925
rect 7834 25916 7840 25928
rect 7892 25916 7898 25968
rect 8202 25956 8208 25968
rect 8163 25928 8208 25956
rect 8202 25916 8208 25928
rect 8260 25916 8266 25968
rect 9217 25959 9275 25965
rect 9217 25925 9229 25959
rect 9263 25956 9275 25959
rect 9306 25956 9312 25968
rect 9263 25928 9312 25956
rect 9263 25925 9275 25928
rect 9217 25919 9275 25925
rect 9306 25916 9312 25928
rect 9364 25956 9370 25968
rect 9766 25956 9772 25968
rect 9364 25928 9772 25956
rect 9364 25916 9370 25928
rect 9766 25916 9772 25928
rect 9824 25916 9830 25968
rect 11146 25916 11152 25968
rect 11204 25956 11210 25968
rect 11204 25928 12664 25956
rect 11204 25916 11210 25928
rect 2740 25860 6684 25888
rect 2740 25848 2746 25860
rect 6730 25848 6736 25900
rect 6788 25888 6794 25900
rect 6963 25891 7021 25897
rect 6963 25888 6975 25891
rect 6788 25860 6975 25888
rect 6788 25848 6794 25860
rect 6963 25857 6975 25860
rect 7009 25857 7021 25891
rect 6963 25851 7021 25857
rect 8297 25891 8355 25897
rect 8297 25857 8309 25891
rect 8343 25888 8355 25891
rect 8386 25888 8392 25900
rect 8343 25860 8392 25888
rect 8343 25857 8355 25860
rect 8297 25851 8355 25857
rect 8386 25848 8392 25860
rect 8444 25848 8450 25900
rect 9953 25891 10011 25897
rect 9953 25888 9965 25891
rect 9646 25860 9965 25888
rect 3789 25823 3847 25829
rect 3789 25789 3801 25823
rect 3835 25820 3847 25823
rect 3970 25820 3976 25832
rect 3835 25792 3976 25820
rect 3835 25789 3847 25792
rect 3789 25783 3847 25789
rect 3970 25780 3976 25792
rect 4028 25820 4034 25832
rect 4249 25823 4307 25829
rect 4249 25820 4261 25823
rect 4028 25792 4261 25820
rect 4028 25780 4034 25792
rect 4249 25789 4261 25792
rect 4295 25789 4307 25823
rect 4249 25783 4307 25789
rect 6876 25823 6934 25829
rect 6876 25789 6888 25823
rect 6922 25820 6934 25823
rect 7650 25820 7656 25832
rect 6922 25792 7656 25820
rect 6922 25789 6934 25792
rect 6876 25783 6934 25789
rect 7650 25780 7656 25792
rect 7708 25780 7714 25832
rect 4154 25752 4160 25764
rect 4115 25724 4160 25752
rect 4154 25712 4160 25724
rect 4212 25752 4218 25764
rect 4570 25755 4628 25761
rect 4570 25752 4582 25755
rect 4212 25724 4582 25752
rect 4212 25712 4218 25724
rect 4570 25721 4582 25724
rect 4616 25721 4628 25755
rect 4570 25715 4628 25721
rect 8202 25712 8208 25764
rect 8260 25752 8266 25764
rect 8618 25755 8676 25761
rect 8618 25752 8630 25755
rect 8260 25724 8630 25752
rect 8260 25712 8266 25724
rect 8618 25721 8630 25724
rect 8664 25752 8676 25755
rect 9646 25752 9674 25860
rect 8664 25724 9674 25752
rect 9784 25752 9812 25860
rect 9953 25857 9965 25860
rect 9999 25857 10011 25891
rect 12526 25888 12532 25900
rect 12487 25860 12532 25888
rect 9953 25851 10011 25857
rect 12526 25848 12532 25860
rect 12584 25848 12590 25900
rect 12636 25888 12664 25928
rect 12805 25891 12863 25897
rect 12805 25888 12817 25891
rect 12636 25860 12817 25888
rect 12805 25857 12817 25860
rect 12851 25857 12863 25891
rect 12805 25851 12863 25857
rect 9858 25780 9864 25832
rect 9916 25820 9922 25832
rect 10045 25823 10103 25829
rect 10045 25820 10057 25823
rect 9916 25792 10057 25820
rect 9916 25780 9922 25792
rect 10045 25789 10057 25792
rect 10091 25820 10103 25823
rect 10686 25820 10692 25832
rect 10091 25792 10692 25820
rect 10091 25789 10103 25792
rect 10045 25783 10103 25789
rect 10686 25780 10692 25792
rect 10744 25780 10750 25832
rect 10410 25761 10416 25764
rect 10366 25755 10416 25761
rect 10366 25752 10378 25755
rect 9784 25724 10378 25752
rect 8664 25721 8676 25724
rect 8618 25715 8676 25721
rect 10366 25721 10378 25724
rect 10412 25721 10416 25755
rect 10366 25715 10416 25721
rect 10410 25712 10416 25715
rect 10468 25712 10474 25764
rect 11330 25752 11336 25764
rect 11243 25724 11336 25752
rect 11330 25712 11336 25724
rect 11388 25752 11394 25764
rect 12618 25752 12624 25764
rect 11388 25724 12624 25752
rect 11388 25712 11394 25724
rect 12618 25712 12624 25724
rect 12676 25712 12682 25764
rect 4798 25644 4804 25696
rect 4856 25684 4862 25696
rect 5445 25687 5503 25693
rect 5445 25684 5457 25687
rect 4856 25656 5457 25684
rect 4856 25644 4862 25656
rect 5445 25653 5457 25656
rect 5491 25653 5503 25687
rect 6086 25684 6092 25696
rect 6047 25656 6092 25684
rect 5445 25647 5503 25653
rect 6086 25644 6092 25656
rect 6144 25644 6150 25696
rect 12250 25684 12256 25696
rect 12211 25656 12256 25684
rect 12250 25644 12256 25656
rect 12308 25644 12314 25696
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 4154 25440 4160 25492
rect 4212 25480 4218 25492
rect 4341 25483 4399 25489
rect 4341 25480 4353 25483
rect 4212 25452 4353 25480
rect 4212 25440 4218 25452
rect 4341 25449 4353 25452
rect 4387 25480 4399 25483
rect 5258 25480 5264 25492
rect 4387 25452 5264 25480
rect 4387 25449 4399 25452
rect 4341 25443 4399 25449
rect 5258 25440 5264 25452
rect 5316 25440 5322 25492
rect 5813 25483 5871 25489
rect 5813 25449 5825 25483
rect 5859 25480 5871 25483
rect 6086 25480 6092 25492
rect 5859 25452 6092 25480
rect 5859 25449 5871 25452
rect 5813 25443 5871 25449
rect 6086 25440 6092 25452
rect 6144 25440 6150 25492
rect 8386 25480 8392 25492
rect 8347 25452 8392 25480
rect 8386 25440 8392 25452
rect 8444 25440 8450 25492
rect 8846 25440 8852 25492
rect 8904 25480 8910 25492
rect 8941 25483 8999 25489
rect 8941 25480 8953 25483
rect 8904 25452 8953 25480
rect 8904 25440 8910 25452
rect 8941 25449 8953 25452
rect 8987 25449 8999 25483
rect 9950 25480 9956 25492
rect 9911 25452 9956 25480
rect 8941 25443 8999 25449
rect 9950 25440 9956 25452
rect 10008 25440 10014 25492
rect 10410 25480 10416 25492
rect 10371 25452 10416 25480
rect 10410 25440 10416 25452
rect 10468 25440 10474 25492
rect 10965 25483 11023 25489
rect 10965 25449 10977 25483
rect 11011 25480 11023 25483
rect 11330 25480 11336 25492
rect 11011 25452 11336 25480
rect 11011 25449 11023 25452
rect 10965 25443 11023 25449
rect 11330 25440 11336 25452
rect 11388 25440 11394 25492
rect 12526 25440 12532 25492
rect 12584 25480 12590 25492
rect 12989 25483 13047 25489
rect 12989 25480 13001 25483
rect 12584 25452 13001 25480
rect 12584 25440 12590 25452
rect 12989 25449 13001 25452
rect 13035 25449 13047 25483
rect 12989 25443 13047 25449
rect 6730 25372 6736 25424
rect 6788 25412 6794 25424
rect 7095 25415 7153 25421
rect 7095 25412 7107 25415
rect 6788 25384 7107 25412
rect 6788 25372 6794 25384
rect 7095 25381 7107 25384
rect 7141 25412 7153 25415
rect 8202 25412 8208 25424
rect 7141 25384 8208 25412
rect 7141 25381 7153 25384
rect 7095 25375 7153 25381
rect 8202 25372 8208 25384
rect 8260 25372 8266 25424
rect 10428 25412 10456 25440
rect 11790 25412 11796 25424
rect 10428 25384 11796 25412
rect 11790 25372 11796 25384
rect 11848 25412 11854 25424
rect 12114 25415 12172 25421
rect 12114 25412 12126 25415
rect 11848 25384 12126 25412
rect 11848 25372 11854 25384
rect 12114 25381 12126 25384
rect 12160 25381 12172 25415
rect 12114 25375 12172 25381
rect 2682 25344 2688 25356
rect 2643 25316 2688 25344
rect 2682 25304 2688 25316
rect 2740 25304 2746 25356
rect 2866 25344 2872 25356
rect 2827 25316 2872 25344
rect 2866 25304 2872 25316
rect 2924 25304 2930 25356
rect 3145 25347 3203 25353
rect 3145 25313 3157 25347
rect 3191 25344 3203 25347
rect 9858 25344 9864 25356
rect 3191 25316 9864 25344
rect 3191 25313 3203 25316
rect 3145 25307 3203 25313
rect 9858 25304 9864 25316
rect 9916 25304 9922 25356
rect 10042 25344 10048 25356
rect 10003 25316 10048 25344
rect 10042 25304 10048 25316
rect 10100 25304 10106 25356
rect 11974 25304 11980 25356
rect 12032 25344 12038 25356
rect 12713 25347 12771 25353
rect 12713 25344 12725 25347
rect 12032 25316 12725 25344
rect 12032 25304 12038 25316
rect 12713 25313 12725 25316
rect 12759 25313 12771 25347
rect 13538 25344 13544 25356
rect 13499 25316 13544 25344
rect 12713 25307 12771 25313
rect 13538 25304 13544 25316
rect 13596 25304 13602 25356
rect 4893 25279 4951 25285
rect 4893 25276 4905 25279
rect 4724 25248 4905 25276
rect 4338 25100 4344 25152
rect 4396 25140 4402 25152
rect 4724 25149 4752 25248
rect 4893 25245 4905 25248
rect 4939 25245 4951 25279
rect 4893 25239 4951 25245
rect 6733 25279 6791 25285
rect 6733 25245 6745 25279
rect 6779 25245 6791 25279
rect 8478 25276 8484 25288
rect 8439 25248 8484 25276
rect 6733 25239 6791 25245
rect 4709 25143 4767 25149
rect 4709 25140 4721 25143
rect 4396 25112 4721 25140
rect 4396 25100 4402 25112
rect 4709 25109 4721 25112
rect 4755 25109 4767 25143
rect 4709 25103 4767 25109
rect 5902 25100 5908 25152
rect 5960 25140 5966 25152
rect 6549 25143 6607 25149
rect 6549 25140 6561 25143
rect 5960 25112 6561 25140
rect 5960 25100 5966 25112
rect 6549 25109 6561 25112
rect 6595 25140 6607 25143
rect 6748 25140 6776 25239
rect 8478 25236 8484 25248
rect 8536 25236 8542 25288
rect 11793 25279 11851 25285
rect 11793 25245 11805 25279
rect 11839 25276 11851 25279
rect 12066 25276 12072 25288
rect 11839 25248 12072 25276
rect 11839 25245 11851 25248
rect 11793 25239 11851 25245
rect 12066 25236 12072 25248
rect 12124 25236 12130 25288
rect 9490 25168 9496 25220
rect 9548 25208 9554 25220
rect 13679 25211 13737 25217
rect 13679 25208 13691 25211
rect 9548 25180 13691 25208
rect 9548 25168 9554 25180
rect 13679 25177 13691 25180
rect 13725 25177 13737 25211
rect 13679 25171 13737 25177
rect 6595 25112 6776 25140
rect 6595 25109 6607 25112
rect 6549 25103 6607 25109
rect 7282 25100 7288 25152
rect 7340 25140 7346 25152
rect 7653 25143 7711 25149
rect 7653 25140 7665 25143
rect 7340 25112 7665 25140
rect 7340 25100 7346 25112
rect 7653 25109 7665 25112
rect 7699 25140 7711 25143
rect 7929 25143 7987 25149
rect 7929 25140 7941 25143
rect 7699 25112 7941 25140
rect 7699 25109 7711 25112
rect 7653 25103 7711 25109
rect 7929 25109 7941 25112
rect 7975 25109 7987 25143
rect 7929 25103 7987 25109
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 2501 24939 2559 24945
rect 2501 24905 2513 24939
rect 2547 24936 2559 24939
rect 2682 24936 2688 24948
rect 2547 24908 2688 24936
rect 2547 24905 2559 24908
rect 2501 24899 2559 24905
rect 2682 24896 2688 24908
rect 2740 24896 2746 24948
rect 2866 24936 2872 24948
rect 2827 24908 2872 24936
rect 2866 24896 2872 24908
rect 2924 24896 2930 24948
rect 4985 24939 5043 24945
rect 4985 24905 4997 24939
rect 5031 24936 5043 24939
rect 5258 24936 5264 24948
rect 5031 24908 5264 24936
rect 5031 24905 5043 24908
rect 4985 24899 5043 24905
rect 5258 24896 5264 24908
rect 5316 24936 5322 24948
rect 6641 24939 6699 24945
rect 6641 24936 6653 24939
rect 5316 24908 6653 24936
rect 5316 24896 5322 24908
rect 6641 24905 6653 24908
rect 6687 24936 6699 24939
rect 6730 24936 6736 24948
rect 6687 24908 6736 24936
rect 6687 24905 6699 24908
rect 6641 24899 6699 24905
rect 6730 24896 6736 24908
rect 6788 24896 6794 24948
rect 8205 24939 8263 24945
rect 8205 24905 8217 24939
rect 8251 24936 8263 24939
rect 8478 24936 8484 24948
rect 8251 24908 8484 24936
rect 8251 24905 8263 24908
rect 8205 24899 8263 24905
rect 3970 24760 3976 24812
rect 4028 24800 4034 24812
rect 4157 24803 4215 24809
rect 4157 24800 4169 24803
rect 4028 24772 4169 24800
rect 4028 24760 4034 24772
rect 4157 24769 4169 24772
rect 4203 24769 4215 24803
rect 5902 24800 5908 24812
rect 5863 24772 5908 24800
rect 4157 24763 4215 24769
rect 5902 24760 5908 24772
rect 5960 24760 5966 24812
rect 7193 24803 7251 24809
rect 7193 24769 7205 24803
rect 7239 24800 7251 24803
rect 8220 24800 8248 24899
rect 8478 24896 8484 24908
rect 8536 24896 8542 24948
rect 10045 24939 10103 24945
rect 10045 24905 10057 24939
rect 10091 24936 10103 24939
rect 10226 24936 10232 24948
rect 10091 24908 10232 24936
rect 10091 24905 10103 24908
rect 10045 24899 10103 24905
rect 10226 24896 10232 24908
rect 10284 24936 10290 24948
rect 10410 24936 10416 24948
rect 10284 24908 10416 24936
rect 10284 24896 10290 24908
rect 10410 24896 10416 24908
rect 10468 24936 10474 24948
rect 10686 24936 10692 24948
rect 10468 24908 10692 24936
rect 10468 24896 10474 24908
rect 10686 24896 10692 24908
rect 10744 24896 10750 24948
rect 11790 24936 11796 24948
rect 11751 24908 11796 24936
rect 11790 24896 11796 24908
rect 11848 24896 11854 24948
rect 13538 24936 13544 24948
rect 13499 24908 13544 24936
rect 13538 24896 13544 24908
rect 13596 24896 13602 24948
rect 8846 24800 8852 24812
rect 7239 24772 8248 24800
rect 8807 24772 8852 24800
rect 7239 24769 7251 24772
rect 7193 24763 7251 24769
rect 8846 24760 8852 24772
rect 8904 24760 8910 24812
rect 9493 24803 9551 24809
rect 9493 24769 9505 24803
rect 9539 24800 9551 24803
rect 11238 24800 11244 24812
rect 9539 24772 11244 24800
rect 9539 24769 9551 24772
rect 9493 24763 9551 24769
rect 11238 24760 11244 24772
rect 11296 24760 11302 24812
rect 13078 24800 13084 24812
rect 12728 24772 13084 24800
rect 3605 24735 3663 24741
rect 3605 24732 3617 24735
rect 3436 24704 3617 24732
rect 3436 24608 3464 24704
rect 3605 24701 3617 24704
rect 3651 24701 3663 24735
rect 3605 24695 3663 24701
rect 4065 24735 4123 24741
rect 4065 24701 4077 24735
rect 4111 24732 4123 24735
rect 5445 24735 5503 24741
rect 4111 24704 4200 24732
rect 4111 24701 4123 24704
rect 4065 24695 4123 24701
rect 4172 24676 4200 24704
rect 5445 24701 5457 24735
rect 5491 24701 5503 24735
rect 5626 24732 5632 24744
rect 5587 24704 5632 24732
rect 5445 24695 5503 24701
rect 4154 24624 4160 24676
rect 4212 24624 4218 24676
rect 5460 24664 5488 24695
rect 5626 24692 5632 24704
rect 5684 24692 5690 24744
rect 10502 24732 10508 24744
rect 10463 24704 10508 24732
rect 10502 24692 10508 24704
rect 10560 24692 10566 24744
rect 12728 24741 12756 24772
rect 13078 24760 13084 24772
rect 13136 24760 13142 24812
rect 12253 24735 12311 24741
rect 12253 24732 12265 24735
rect 10612 24704 12265 24732
rect 6273 24667 6331 24673
rect 6273 24664 6285 24667
rect 5460 24636 6285 24664
rect 6273 24633 6285 24636
rect 6319 24664 6331 24667
rect 6638 24664 6644 24676
rect 6319 24636 6644 24664
rect 6319 24633 6331 24636
rect 6273 24627 6331 24633
rect 6638 24624 6644 24636
rect 6696 24664 6702 24676
rect 6696 24636 7230 24664
rect 6696 24624 6702 24636
rect 3418 24596 3424 24608
rect 3379 24568 3424 24596
rect 3418 24556 3424 24568
rect 3476 24556 3482 24608
rect 7202 24596 7230 24636
rect 7282 24624 7288 24676
rect 7340 24664 7346 24676
rect 7340 24636 7385 24664
rect 7340 24624 7346 24636
rect 7650 24624 7656 24676
rect 7708 24664 7714 24676
rect 7837 24667 7895 24673
rect 7837 24664 7849 24667
rect 7708 24636 7849 24664
rect 7708 24624 7714 24636
rect 7837 24633 7849 24636
rect 7883 24633 7895 24667
rect 7837 24627 7895 24633
rect 8665 24667 8723 24673
rect 8665 24633 8677 24667
rect 8711 24664 8723 24667
rect 8941 24667 8999 24673
rect 8941 24664 8953 24667
rect 8711 24636 8953 24664
rect 8711 24633 8723 24636
rect 8665 24627 8723 24633
rect 8941 24633 8953 24636
rect 8987 24664 8999 24667
rect 9306 24664 9312 24676
rect 8987 24636 9312 24664
rect 8987 24633 8999 24636
rect 8941 24627 8999 24633
rect 9306 24624 9312 24636
rect 9364 24624 9370 24676
rect 10410 24624 10416 24676
rect 10468 24664 10474 24676
rect 10612 24664 10640 24704
rect 12253 24701 12265 24704
rect 12299 24732 12311 24735
rect 12713 24735 12771 24741
rect 12713 24732 12725 24735
rect 12299 24704 12725 24732
rect 12299 24701 12311 24704
rect 12253 24695 12311 24701
rect 12713 24701 12725 24704
rect 12759 24701 12771 24735
rect 12894 24732 12900 24744
rect 12855 24704 12900 24732
rect 12713 24695 12771 24701
rect 12894 24692 12900 24704
rect 12952 24692 12958 24744
rect 10468 24636 10640 24664
rect 10468 24624 10474 24636
rect 10686 24624 10692 24676
rect 10744 24664 10750 24676
rect 10826 24667 10884 24673
rect 10826 24664 10838 24667
rect 10744 24636 10838 24664
rect 10744 24624 10750 24636
rect 10826 24633 10838 24636
rect 10872 24633 10884 24667
rect 10826 24627 10884 24633
rect 8110 24596 8116 24608
rect 7202 24568 8116 24596
rect 8110 24556 8116 24568
rect 8168 24556 8174 24608
rect 11422 24596 11428 24608
rect 11383 24568 11428 24596
rect 11422 24556 11428 24568
rect 11480 24556 11486 24608
rect 12526 24596 12532 24608
rect 12487 24568 12532 24596
rect 12526 24556 12532 24568
rect 12584 24556 12590 24608
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 6086 24352 6092 24404
rect 6144 24392 6150 24404
rect 8754 24392 8760 24404
rect 6144 24364 8760 24392
rect 6144 24352 6150 24364
rect 8754 24352 8760 24364
rect 8812 24352 8818 24404
rect 9674 24352 9680 24404
rect 9732 24392 9738 24404
rect 10137 24395 10195 24401
rect 10137 24392 10149 24395
rect 9732 24364 10149 24392
rect 9732 24352 9738 24364
rect 10137 24361 10149 24364
rect 10183 24361 10195 24395
rect 10137 24355 10195 24361
rect 10502 24352 10508 24404
rect 10560 24392 10566 24404
rect 10965 24395 11023 24401
rect 10965 24392 10977 24395
rect 10560 24364 10977 24392
rect 10560 24352 10566 24364
rect 10965 24361 10977 24364
rect 11011 24392 11023 24395
rect 12526 24392 12532 24404
rect 11011 24364 12532 24392
rect 11011 24361 11023 24364
rect 10965 24355 11023 24361
rect 12526 24352 12532 24364
rect 12584 24352 12590 24404
rect 4798 24324 4804 24336
rect 4759 24296 4804 24324
rect 4798 24284 4804 24296
rect 4856 24284 4862 24336
rect 6549 24327 6607 24333
rect 6549 24293 6561 24327
rect 6595 24324 6607 24327
rect 7193 24327 7251 24333
rect 7193 24324 7205 24327
rect 6595 24296 7205 24324
rect 6595 24293 6607 24296
rect 6549 24287 6607 24293
rect 7193 24293 7205 24296
rect 7239 24324 7251 24327
rect 7282 24324 7288 24336
rect 7239 24296 7288 24324
rect 7239 24293 7251 24296
rect 7193 24287 7251 24293
rect 7282 24284 7288 24296
rect 7340 24284 7346 24336
rect 11241 24327 11299 24333
rect 11241 24293 11253 24327
rect 11287 24324 11299 24327
rect 11422 24324 11428 24336
rect 11287 24296 11428 24324
rect 11287 24293 11299 24296
rect 11241 24287 11299 24293
rect 11422 24284 11428 24296
rect 11480 24284 11486 24336
rect 2958 24256 2964 24268
rect 2919 24228 2964 24256
rect 2958 24216 2964 24228
rect 3016 24216 3022 24268
rect 3970 24216 3976 24268
rect 4028 24256 4034 24268
rect 4065 24259 4123 24265
rect 4065 24256 4077 24259
rect 4028 24228 4077 24256
rect 4028 24216 4034 24228
rect 4065 24225 4077 24228
rect 4111 24225 4123 24259
rect 4065 24219 4123 24225
rect 4080 24188 4108 24219
rect 4154 24216 4160 24268
rect 4212 24256 4218 24268
rect 4525 24259 4583 24265
rect 4525 24256 4537 24259
rect 4212 24228 4537 24256
rect 4212 24216 4218 24228
rect 4525 24225 4537 24228
rect 4571 24225 4583 24259
rect 5994 24256 6000 24268
rect 5955 24228 6000 24256
rect 4525 24219 4583 24225
rect 5994 24216 6000 24228
rect 6052 24216 6058 24268
rect 8570 24256 8576 24268
rect 8531 24228 8576 24256
rect 8570 24216 8576 24228
rect 8628 24216 8634 24268
rect 9677 24259 9735 24265
rect 9677 24225 9689 24259
rect 9723 24256 9735 24259
rect 9766 24256 9772 24268
rect 9723 24228 9772 24256
rect 9723 24225 9735 24228
rect 9677 24219 9735 24225
rect 9766 24216 9772 24228
rect 9824 24216 9830 24268
rect 10042 24216 10048 24268
rect 10100 24256 10106 24268
rect 10505 24259 10563 24265
rect 10505 24256 10517 24259
rect 10100 24228 10517 24256
rect 10100 24216 10106 24228
rect 10505 24225 10517 24228
rect 10551 24225 10563 24259
rect 12618 24256 12624 24268
rect 12579 24228 12624 24256
rect 10505 24219 10563 24225
rect 12618 24216 12624 24228
rect 12676 24216 12682 24268
rect 7101 24191 7159 24197
rect 4080 24160 4154 24188
rect 4126 24120 4154 24160
rect 7101 24157 7113 24191
rect 7147 24188 7159 24191
rect 7926 24188 7932 24200
rect 7147 24160 7932 24188
rect 7147 24157 7159 24160
rect 7101 24151 7159 24157
rect 7926 24148 7932 24160
rect 7984 24148 7990 24200
rect 11149 24191 11207 24197
rect 11149 24157 11161 24191
rect 11195 24188 11207 24191
rect 11238 24188 11244 24200
rect 11195 24160 11244 24188
rect 11195 24157 11207 24160
rect 11149 24151 11207 24157
rect 11238 24148 11244 24160
rect 11296 24148 11302 24200
rect 11514 24148 11520 24200
rect 11572 24188 11578 24200
rect 11790 24188 11796 24200
rect 11572 24160 11796 24188
rect 11572 24148 11578 24160
rect 11790 24148 11796 24160
rect 11848 24148 11854 24200
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 12529 24191 12587 24197
rect 12529 24188 12541 24191
rect 11931 24160 12541 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 12529 24157 12541 24160
rect 12575 24188 12587 24191
rect 12894 24188 12900 24200
rect 12575 24160 12900 24188
rect 12575 24157 12587 24160
rect 12529 24151 12587 24157
rect 12894 24148 12900 24160
rect 12952 24148 12958 24200
rect 4890 24120 4896 24132
rect 4126 24092 4896 24120
rect 4890 24080 4896 24092
rect 4948 24080 4954 24132
rect 5534 24080 5540 24132
rect 5592 24120 5598 24132
rect 6181 24123 6239 24129
rect 6181 24120 6193 24123
rect 5592 24092 6193 24120
rect 5592 24080 5598 24092
rect 6181 24089 6193 24092
rect 6227 24089 6239 24123
rect 7650 24120 7656 24132
rect 7611 24092 7656 24120
rect 6181 24083 6239 24089
rect 7650 24080 7656 24092
rect 7708 24080 7714 24132
rect 8202 24080 8208 24132
rect 8260 24120 8266 24132
rect 8260 24092 9260 24120
rect 8260 24080 8266 24092
rect 2406 24012 2412 24064
rect 2464 24052 2470 24064
rect 3145 24055 3203 24061
rect 3145 24052 3157 24055
rect 2464 24024 3157 24052
rect 2464 24012 2470 24024
rect 3145 24021 3157 24024
rect 3191 24052 3203 24055
rect 3418 24052 3424 24064
rect 3191 24024 3424 24052
rect 3191 24021 3203 24024
rect 3145 24015 3203 24021
rect 3418 24012 3424 24024
rect 3476 24012 3482 24064
rect 3697 24055 3755 24061
rect 3697 24021 3709 24055
rect 3743 24052 3755 24055
rect 4154 24052 4160 24064
rect 3743 24024 4160 24052
rect 3743 24021 3755 24024
rect 3697 24015 3755 24021
rect 4154 24012 4160 24024
rect 4212 24012 4218 24064
rect 5261 24055 5319 24061
rect 5261 24021 5273 24055
rect 5307 24052 5319 24055
rect 5626 24052 5632 24064
rect 5307 24024 5632 24052
rect 5307 24021 5319 24024
rect 5261 24015 5319 24021
rect 5626 24012 5632 24024
rect 5684 24012 5690 24064
rect 6822 24052 6828 24064
rect 6783 24024 6828 24052
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 7190 24012 7196 24064
rect 7248 24052 7254 24064
rect 8757 24055 8815 24061
rect 8757 24052 8769 24055
rect 7248 24024 8769 24052
rect 7248 24012 7254 24024
rect 8757 24021 8769 24024
rect 8803 24021 8815 24055
rect 8757 24015 8815 24021
rect 8846 24012 8852 24064
rect 8904 24052 8910 24064
rect 9033 24055 9091 24061
rect 9033 24052 9045 24055
rect 8904 24024 9045 24052
rect 8904 24012 8910 24024
rect 9033 24021 9045 24024
rect 9079 24021 9091 24055
rect 9232 24052 9260 24092
rect 9398 24080 9404 24132
rect 9456 24120 9462 24132
rect 12759 24123 12817 24129
rect 12759 24120 12771 24123
rect 9456 24092 12771 24120
rect 9456 24080 9462 24092
rect 12759 24089 12771 24092
rect 12805 24089 12817 24123
rect 12759 24083 12817 24089
rect 9582 24052 9588 24064
rect 9232 24024 9588 24052
rect 9033 24015 9091 24021
rect 9582 24012 9588 24024
rect 9640 24052 9646 24064
rect 9861 24055 9919 24061
rect 9861 24052 9873 24055
rect 9640 24024 9873 24052
rect 9640 24012 9646 24024
rect 9861 24021 9873 24024
rect 9907 24052 9919 24055
rect 11885 24055 11943 24061
rect 11885 24052 11897 24055
rect 9907 24024 11897 24052
rect 9907 24021 9919 24024
rect 9861 24015 9919 24021
rect 11885 24021 11897 24024
rect 11931 24021 11943 24055
rect 12066 24052 12072 24064
rect 12027 24024 12072 24052
rect 11885 24015 11943 24021
rect 12066 24012 12072 24024
rect 12124 24012 12130 24064
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 2777 23851 2835 23857
rect 2777 23817 2789 23851
rect 2823 23848 2835 23851
rect 3970 23848 3976 23860
rect 2823 23820 3976 23848
rect 2823 23817 2835 23820
rect 2777 23811 2835 23817
rect 3970 23808 3976 23820
rect 4028 23808 4034 23860
rect 8202 23848 8208 23860
rect 4126 23820 8208 23848
rect 4126 23792 4154 23820
rect 8202 23808 8208 23820
rect 8260 23808 8266 23860
rect 8386 23808 8392 23860
rect 8444 23848 8450 23860
rect 8481 23851 8539 23857
rect 8481 23848 8493 23851
rect 8444 23820 8493 23848
rect 8444 23808 8450 23820
rect 8481 23817 8493 23820
rect 8527 23848 8539 23851
rect 8570 23848 8576 23860
rect 8527 23820 8576 23848
rect 8527 23817 8539 23820
rect 8481 23811 8539 23817
rect 8570 23808 8576 23820
rect 8628 23808 8634 23860
rect 11241 23851 11299 23857
rect 11241 23817 11253 23851
rect 11287 23848 11299 23851
rect 11422 23848 11428 23860
rect 11287 23820 11428 23848
rect 11287 23817 11299 23820
rect 11241 23811 11299 23817
rect 11422 23808 11428 23820
rect 11480 23808 11486 23860
rect 2501 23783 2559 23789
rect 2501 23749 2513 23783
rect 2547 23780 2559 23783
rect 2958 23780 2964 23792
rect 2547 23752 2964 23780
rect 2547 23749 2559 23752
rect 2501 23743 2559 23749
rect 2958 23740 2964 23752
rect 3016 23740 3022 23792
rect 4062 23740 4068 23792
rect 4120 23752 4154 23792
rect 6641 23783 6699 23789
rect 4120 23740 4126 23752
rect 6641 23749 6653 23783
rect 6687 23780 6699 23783
rect 6730 23780 6736 23792
rect 6687 23752 6736 23780
rect 6687 23749 6699 23752
rect 6641 23743 6699 23749
rect 6730 23740 6736 23752
rect 6788 23780 6794 23792
rect 6788 23752 6960 23780
rect 6788 23740 6794 23752
rect 4338 23712 4344 23724
rect 4299 23684 4344 23712
rect 4338 23672 4344 23684
rect 4396 23672 4402 23724
rect 6822 23712 6828 23724
rect 6783 23684 6828 23712
rect 6822 23672 6828 23684
rect 6880 23672 6886 23724
rect 2593 23647 2651 23653
rect 2593 23613 2605 23647
rect 2639 23644 2651 23647
rect 3142 23644 3148 23656
rect 2639 23616 3148 23644
rect 2639 23613 2651 23616
rect 2593 23607 2651 23613
rect 3142 23604 3148 23616
rect 3200 23604 3206 23656
rect 3326 23604 3332 23656
rect 3384 23644 3390 23656
rect 3513 23647 3571 23653
rect 3513 23644 3525 23647
rect 3384 23616 3525 23644
rect 3384 23604 3390 23616
rect 3513 23613 3525 23616
rect 3559 23644 3571 23647
rect 3605 23647 3663 23653
rect 3605 23644 3617 23647
rect 3559 23616 3617 23644
rect 3559 23613 3571 23616
rect 3513 23607 3571 23613
rect 3605 23613 3617 23616
rect 3651 23613 3663 23647
rect 3605 23607 3663 23613
rect 4154 23604 4160 23656
rect 4212 23644 4218 23656
rect 5169 23647 5227 23653
rect 5169 23644 5181 23647
rect 4212 23616 4305 23644
rect 5000 23616 5181 23644
rect 4212 23604 4218 23616
rect 2958 23536 2964 23588
rect 3016 23576 3022 23588
rect 3418 23576 3424 23588
rect 3016 23548 3424 23576
rect 3016 23536 3022 23548
rect 3418 23536 3424 23548
rect 3476 23536 3482 23588
rect 4172 23576 4200 23604
rect 4338 23576 4344 23588
rect 4172 23548 4344 23576
rect 4338 23536 4344 23548
rect 4396 23536 4402 23588
rect 4430 23536 4436 23588
rect 4488 23576 4494 23588
rect 5000 23585 5028 23616
rect 5169 23613 5181 23616
rect 5215 23644 5227 23647
rect 5534 23644 5540 23656
rect 5215 23616 5540 23644
rect 5215 23613 5227 23616
rect 5169 23607 5227 23613
rect 5534 23604 5540 23616
rect 5592 23604 5598 23656
rect 5626 23604 5632 23656
rect 5684 23644 5690 23656
rect 5721 23647 5779 23653
rect 5721 23644 5733 23647
rect 5684 23616 5733 23644
rect 5684 23604 5690 23616
rect 5721 23613 5733 23616
rect 5767 23644 5779 23647
rect 6178 23644 6184 23656
rect 5767 23616 6184 23644
rect 5767 23613 5779 23616
rect 5721 23607 5779 23613
rect 6178 23604 6184 23616
rect 6236 23604 6242 23656
rect 6932 23588 6960 23752
rect 7650 23740 7656 23792
rect 7708 23780 7714 23792
rect 7708 23752 8984 23780
rect 7708 23740 7714 23752
rect 8662 23712 8668 23724
rect 8575 23684 8668 23712
rect 8662 23672 8668 23684
rect 8720 23712 8726 23724
rect 8846 23712 8852 23724
rect 8720 23684 8852 23712
rect 8720 23672 8726 23684
rect 8846 23672 8852 23684
rect 8904 23672 8910 23724
rect 8956 23721 8984 23752
rect 10594 23740 10600 23792
rect 10652 23780 10658 23792
rect 12618 23780 12624 23792
rect 10652 23752 12624 23780
rect 10652 23740 10658 23752
rect 12618 23740 12624 23752
rect 12676 23740 12682 23792
rect 8941 23715 8999 23721
rect 8941 23681 8953 23715
rect 8987 23681 8999 23715
rect 8941 23675 8999 23681
rect 10873 23715 10931 23721
rect 10873 23681 10885 23715
rect 10919 23712 10931 23715
rect 12066 23712 12072 23724
rect 10919 23684 12072 23712
rect 10919 23681 10931 23684
rect 10873 23675 10931 23681
rect 12066 23672 12072 23684
rect 12124 23672 12130 23724
rect 12250 23672 12256 23724
rect 12308 23712 12314 23724
rect 12434 23712 12440 23724
rect 12308 23684 12440 23712
rect 12308 23672 12314 23684
rect 12434 23672 12440 23684
rect 12492 23672 12498 23724
rect 10045 23647 10103 23653
rect 10045 23613 10057 23647
rect 10091 23644 10103 23647
rect 10410 23644 10416 23656
rect 10091 23616 10416 23644
rect 10091 23613 10103 23616
rect 10045 23607 10103 23613
rect 4985 23579 5043 23585
rect 4985 23576 4997 23579
rect 4488 23548 4997 23576
rect 4488 23536 4494 23548
rect 4985 23545 4997 23548
rect 5031 23545 5043 23579
rect 5902 23576 5908 23588
rect 5863 23548 5908 23576
rect 4985 23539 5043 23545
rect 5902 23536 5908 23548
rect 5960 23536 5966 23588
rect 5994 23536 6000 23588
rect 6052 23576 6058 23588
rect 6273 23579 6331 23585
rect 6273 23576 6285 23579
rect 6052 23548 6285 23576
rect 6052 23536 6058 23548
rect 6273 23545 6285 23548
rect 6319 23576 6331 23579
rect 6730 23576 6736 23588
rect 6319 23548 6736 23576
rect 6319 23545 6331 23548
rect 6273 23539 6331 23545
rect 6730 23536 6736 23548
rect 6788 23536 6794 23588
rect 6914 23576 6920 23588
rect 6827 23548 6920 23576
rect 6914 23536 6920 23548
rect 6972 23576 6978 23588
rect 7146 23579 7204 23585
rect 7146 23576 7158 23579
rect 6972 23548 7158 23576
rect 6972 23536 6978 23548
rect 7146 23545 7158 23548
rect 7192 23545 7204 23579
rect 7146 23539 7204 23545
rect 8757 23579 8815 23585
rect 8757 23545 8769 23579
rect 8803 23545 8815 23579
rect 8757 23539 8815 23545
rect 3142 23508 3148 23520
rect 3103 23480 3148 23508
rect 3142 23468 3148 23480
rect 3200 23468 3206 23520
rect 4709 23511 4767 23517
rect 4709 23477 4721 23511
rect 4755 23508 4767 23511
rect 4890 23508 4896 23520
rect 4755 23480 4896 23508
rect 4755 23477 4767 23480
rect 4709 23471 4767 23477
rect 4890 23468 4896 23480
rect 4948 23468 4954 23520
rect 7745 23511 7803 23517
rect 7745 23477 7757 23511
rect 7791 23508 7803 23511
rect 8021 23511 8079 23517
rect 8021 23508 8033 23511
rect 7791 23480 8033 23508
rect 7791 23477 7803 23480
rect 7745 23471 7803 23477
rect 8021 23477 8033 23480
rect 8067 23508 8079 23511
rect 8772 23508 8800 23539
rect 8846 23536 8852 23588
rect 8904 23576 8910 23588
rect 10060 23576 10088 23607
rect 10410 23604 10416 23616
rect 10468 23604 10474 23656
rect 10597 23647 10655 23653
rect 10597 23613 10609 23647
rect 10643 23613 10655 23647
rect 10597 23607 10655 23613
rect 8904 23548 10088 23576
rect 8904 23536 8910 23548
rect 8067 23480 8800 23508
rect 9677 23511 9735 23517
rect 8067 23477 8079 23480
rect 8021 23471 8079 23477
rect 9677 23477 9689 23511
rect 9723 23508 9735 23511
rect 9766 23508 9772 23520
rect 9723 23480 9772 23508
rect 9723 23477 9735 23480
rect 9677 23471 9735 23477
rect 9766 23468 9772 23480
rect 9824 23468 9830 23520
rect 10318 23468 10324 23520
rect 10376 23508 10382 23520
rect 10612 23508 10640 23607
rect 11238 23604 11244 23656
rect 11296 23644 11302 23656
rect 11517 23647 11575 23653
rect 11517 23644 11529 23647
rect 11296 23616 11529 23644
rect 11296 23604 11302 23616
rect 11517 23613 11529 23616
rect 11563 23613 11575 23647
rect 11517 23607 11575 23613
rect 11790 23536 11796 23588
rect 11848 23536 11854 23588
rect 10376 23480 10640 23508
rect 11808 23508 11836 23536
rect 12158 23508 12164 23520
rect 11808 23480 12164 23508
rect 10376 23468 10382 23480
rect 12158 23468 12164 23480
rect 12216 23468 12222 23520
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 4338 23304 4344 23316
rect 4299 23276 4344 23304
rect 4338 23264 4344 23276
rect 4396 23264 4402 23316
rect 5902 23264 5908 23316
rect 5960 23304 5966 23316
rect 6181 23307 6239 23313
rect 6181 23304 6193 23307
rect 5960 23276 6193 23304
rect 5960 23264 5966 23276
rect 6181 23273 6193 23276
rect 6227 23304 6239 23307
rect 7282 23304 7288 23316
rect 6227 23276 6408 23304
rect 7243 23276 7288 23304
rect 6227 23273 6239 23276
rect 6181 23267 6239 23273
rect 4982 23236 4988 23248
rect 4943 23208 4988 23236
rect 4982 23196 4988 23208
rect 5040 23196 5046 23248
rect 2866 23128 2872 23180
rect 2924 23168 2930 23180
rect 6380 23177 6408 23276
rect 7282 23264 7288 23276
rect 7340 23264 7346 23316
rect 7926 23304 7932 23316
rect 7887 23276 7932 23304
rect 7926 23264 7932 23276
rect 7984 23264 7990 23316
rect 9490 23264 9496 23316
rect 9548 23304 9554 23316
rect 9861 23307 9919 23313
rect 9861 23304 9873 23307
rect 9548 23276 9873 23304
rect 9548 23264 9554 23276
rect 9861 23273 9873 23276
rect 9907 23304 9919 23307
rect 10318 23304 10324 23316
rect 9907 23276 10324 23304
rect 9907 23273 9919 23276
rect 9861 23267 9919 23273
rect 10318 23264 10324 23276
rect 10376 23264 10382 23316
rect 10686 23264 10692 23316
rect 10744 23304 10750 23316
rect 12342 23304 12348 23316
rect 10744 23276 12348 23304
rect 10744 23264 10750 23276
rect 12342 23264 12348 23276
rect 12400 23264 12406 23316
rect 6727 23239 6785 23245
rect 6727 23205 6739 23239
rect 6773 23236 6785 23239
rect 6914 23236 6920 23248
rect 6773 23208 6920 23236
rect 6773 23205 6785 23208
rect 6727 23199 6785 23205
rect 6914 23196 6920 23208
rect 6972 23196 6978 23248
rect 7834 23196 7840 23248
rect 7892 23236 7898 23248
rect 8846 23236 8852 23248
rect 7892 23208 8852 23236
rect 7892 23196 7898 23208
rect 8846 23196 8852 23208
rect 8904 23196 8910 23248
rect 11241 23239 11299 23245
rect 11241 23205 11253 23239
rect 11287 23236 11299 23239
rect 11514 23236 11520 23248
rect 11287 23208 11520 23236
rect 11287 23205 11299 23208
rect 11241 23199 11299 23205
rect 11514 23196 11520 23208
rect 11572 23196 11578 23248
rect 11793 23239 11851 23245
rect 11793 23205 11805 23239
rect 11839 23236 11851 23239
rect 12158 23236 12164 23248
rect 11839 23208 12164 23236
rect 11839 23205 11851 23208
rect 11793 23199 11851 23205
rect 12158 23196 12164 23208
rect 12216 23196 12222 23248
rect 2961 23171 3019 23177
rect 2961 23168 2973 23171
rect 2924 23140 2973 23168
rect 2924 23128 2930 23140
rect 2961 23137 2973 23140
rect 3007 23137 3019 23171
rect 2961 23131 3019 23137
rect 6365 23171 6423 23177
rect 6365 23137 6377 23171
rect 6411 23137 6423 23171
rect 8110 23168 8116 23180
rect 8071 23140 8116 23168
rect 6365 23131 6423 23137
rect 8110 23128 8116 23140
rect 8168 23128 8174 23180
rect 9674 23168 9680 23180
rect 9635 23140 9680 23168
rect 9674 23128 9680 23140
rect 9732 23168 9738 23180
rect 10137 23171 10195 23177
rect 10137 23168 10149 23171
rect 9732 23140 10149 23168
rect 9732 23128 9738 23140
rect 10137 23137 10149 23140
rect 10183 23137 10195 23171
rect 10137 23131 10195 23137
rect 3510 23060 3516 23112
rect 3568 23100 3574 23112
rect 4893 23103 4951 23109
rect 4893 23100 4905 23103
rect 3568 23072 4905 23100
rect 3568 23060 3574 23072
rect 4893 23069 4905 23072
rect 4939 23100 4951 23103
rect 5350 23100 5356 23112
rect 4939 23072 5356 23100
rect 4939 23069 4951 23072
rect 4893 23063 4951 23069
rect 5350 23060 5356 23072
rect 5408 23060 5414 23112
rect 5534 23100 5540 23112
rect 5447 23072 5540 23100
rect 5534 23060 5540 23072
rect 5592 23100 5598 23112
rect 7190 23100 7196 23112
rect 5592 23072 7196 23100
rect 5592 23060 5598 23072
rect 7190 23060 7196 23072
rect 7248 23060 7254 23112
rect 11149 23103 11207 23109
rect 11149 23069 11161 23103
rect 11195 23100 11207 23103
rect 11422 23100 11428 23112
rect 11195 23072 11428 23100
rect 11195 23069 11207 23072
rect 11149 23063 11207 23069
rect 11422 23060 11428 23072
rect 11480 23100 11486 23112
rect 12621 23103 12679 23109
rect 12621 23100 12633 23103
rect 11480 23072 12633 23100
rect 11480 23060 11486 23072
rect 12621 23069 12633 23072
rect 12667 23069 12679 23103
rect 12621 23063 12679 23069
rect 3142 22964 3148 22976
rect 3103 22936 3148 22964
rect 3142 22924 3148 22936
rect 3200 22964 3206 22976
rect 3326 22964 3332 22976
rect 3200 22936 3332 22964
rect 3200 22924 3206 22936
rect 3326 22924 3332 22936
rect 3384 22924 3390 22976
rect 3697 22967 3755 22973
rect 3697 22933 3709 22967
rect 3743 22964 3755 22967
rect 4338 22964 4344 22976
rect 3743 22936 4344 22964
rect 3743 22933 3755 22936
rect 3697 22927 3755 22933
rect 4338 22924 4344 22936
rect 4396 22924 4402 22976
rect 4709 22967 4767 22973
rect 4709 22933 4721 22967
rect 4755 22964 4767 22967
rect 4798 22964 4804 22976
rect 4755 22936 4804 22964
rect 4755 22933 4767 22936
rect 4709 22927 4767 22933
rect 4798 22924 4804 22936
rect 4856 22924 4862 22976
rect 7006 22924 7012 22976
rect 7064 22964 7070 22976
rect 7561 22967 7619 22973
rect 7561 22964 7573 22967
rect 7064 22936 7573 22964
rect 7064 22924 7070 22936
rect 7561 22933 7573 22936
rect 7607 22933 7619 22967
rect 7561 22927 7619 22933
rect 8297 22967 8355 22973
rect 8297 22933 8309 22967
rect 8343 22964 8355 22967
rect 8478 22964 8484 22976
rect 8343 22936 8484 22964
rect 8343 22933 8355 22936
rect 8297 22927 8355 22933
rect 8478 22924 8484 22936
rect 8536 22964 8542 22976
rect 8573 22967 8631 22973
rect 8573 22964 8585 22967
rect 8536 22936 8585 22964
rect 8536 22924 8542 22936
rect 8573 22933 8585 22936
rect 8619 22933 8631 22967
rect 8573 22927 8631 22933
rect 8846 22924 8852 22976
rect 8904 22964 8910 22976
rect 9033 22967 9091 22973
rect 9033 22964 9045 22967
rect 8904 22936 9045 22964
rect 8904 22924 8910 22936
rect 9033 22933 9045 22936
rect 9079 22964 9091 22967
rect 9582 22964 9588 22976
rect 9079 22936 9588 22964
rect 9079 22933 9091 22936
rect 9033 22927 9091 22933
rect 9582 22924 9588 22936
rect 9640 22924 9646 22976
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 2866 22720 2872 22772
rect 2924 22760 2930 22772
rect 2961 22763 3019 22769
rect 2961 22760 2973 22763
rect 2924 22732 2973 22760
rect 2924 22720 2930 22732
rect 2961 22729 2973 22732
rect 3007 22729 3019 22763
rect 3510 22760 3516 22772
rect 3471 22732 3516 22760
rect 2961 22723 3019 22729
rect 3510 22720 3516 22732
rect 3568 22720 3574 22772
rect 4062 22760 4068 22772
rect 4023 22732 4068 22760
rect 4062 22720 4068 22732
rect 4120 22720 4126 22772
rect 4982 22720 4988 22772
rect 5040 22760 5046 22772
rect 5442 22760 5448 22772
rect 5040 22732 5448 22760
rect 5040 22720 5046 22732
rect 5442 22720 5448 22732
rect 5500 22760 5506 22772
rect 5813 22763 5871 22769
rect 5813 22760 5825 22763
rect 5500 22732 5825 22760
rect 5500 22720 5506 22732
rect 5813 22729 5825 22732
rect 5859 22729 5871 22763
rect 5813 22723 5871 22729
rect 6457 22763 6515 22769
rect 6457 22729 6469 22763
rect 6503 22760 6515 22763
rect 6549 22763 6607 22769
rect 6549 22760 6561 22763
rect 6503 22732 6561 22760
rect 6503 22729 6515 22732
rect 6457 22723 6515 22729
rect 6549 22729 6561 22732
rect 6595 22760 6607 22763
rect 6914 22760 6920 22772
rect 6595 22732 6920 22760
rect 6595 22729 6607 22732
rect 6549 22723 6607 22729
rect 6914 22720 6920 22732
rect 6972 22720 6978 22772
rect 11422 22760 11428 22772
rect 11383 22732 11428 22760
rect 11422 22720 11428 22732
rect 11480 22720 11486 22772
rect 12342 22720 12348 22772
rect 12400 22760 12406 22772
rect 12621 22763 12679 22769
rect 12621 22760 12633 22763
rect 12400 22732 12633 22760
rect 12400 22720 12406 22732
rect 12621 22729 12633 22732
rect 12667 22729 12679 22763
rect 12621 22723 12679 22729
rect 3789 22695 3847 22701
rect 3789 22661 3801 22695
rect 3835 22692 3847 22695
rect 4706 22692 4712 22704
rect 3835 22664 4712 22692
rect 3835 22661 3847 22664
rect 3789 22655 3847 22661
rect 4706 22652 4712 22664
rect 4764 22652 4770 22704
rect 5537 22695 5595 22701
rect 5537 22661 5549 22695
rect 5583 22692 5595 22695
rect 7006 22692 7012 22704
rect 5583 22664 7012 22692
rect 5583 22661 5595 22664
rect 5537 22655 5595 22661
rect 7006 22652 7012 22664
rect 7064 22652 7070 22704
rect 7466 22692 7472 22704
rect 7116 22664 7472 22692
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22624 6975 22627
rect 7116 22624 7144 22664
rect 7466 22652 7472 22664
rect 7524 22652 7530 22704
rect 8294 22652 8300 22704
rect 8352 22692 8358 22704
rect 13633 22695 13691 22701
rect 13633 22692 13645 22695
rect 8352 22664 13645 22692
rect 8352 22652 8358 22664
rect 13633 22661 13645 22664
rect 13679 22661 13691 22695
rect 13633 22655 13691 22661
rect 6963 22596 7144 22624
rect 6963 22593 6975 22596
rect 6917 22587 6975 22593
rect 7190 22584 7196 22636
rect 7248 22624 7254 22636
rect 7248 22596 7293 22624
rect 7248 22584 7254 22596
rect 8110 22584 8116 22636
rect 8168 22624 8174 22636
rect 8205 22627 8263 22633
rect 8205 22624 8217 22627
rect 8168 22596 8217 22624
rect 8168 22584 8174 22596
rect 8205 22593 8217 22596
rect 8251 22624 8263 22627
rect 9398 22624 9404 22636
rect 8251 22596 9404 22624
rect 8251 22593 8263 22596
rect 8205 22587 8263 22593
rect 9398 22584 9404 22596
rect 9456 22584 9462 22636
rect 9766 22584 9772 22636
rect 9824 22624 9830 22636
rect 10413 22627 10471 22633
rect 10413 22624 10425 22627
rect 9824 22596 10425 22624
rect 9824 22584 9830 22596
rect 10413 22593 10425 22596
rect 10459 22593 10471 22627
rect 10413 22587 10471 22593
rect 3605 22559 3663 22565
rect 3605 22525 3617 22559
rect 3651 22556 3663 22559
rect 4062 22556 4068 22568
rect 3651 22528 4068 22556
rect 3651 22525 3663 22528
rect 3605 22519 3663 22525
rect 4062 22516 4068 22528
rect 4120 22516 4126 22568
rect 4617 22559 4675 22565
rect 4617 22525 4629 22559
rect 4663 22556 4675 22559
rect 4798 22556 4804 22568
rect 4663 22528 4804 22556
rect 4663 22525 4675 22528
rect 4617 22519 4675 22525
rect 4798 22516 4804 22528
rect 4856 22516 4862 22568
rect 8389 22559 8447 22565
rect 8389 22525 8401 22559
rect 8435 22556 8447 22559
rect 8478 22556 8484 22568
rect 8435 22528 8484 22556
rect 8435 22525 8447 22528
rect 8389 22519 8447 22525
rect 4982 22497 4988 22500
rect 4525 22491 4583 22497
rect 4525 22457 4537 22491
rect 4571 22488 4583 22491
rect 4979 22488 4988 22497
rect 4571 22460 4988 22488
rect 4571 22457 4583 22460
rect 4525 22451 4583 22457
rect 4979 22451 4988 22460
rect 5040 22488 5046 22500
rect 6549 22491 6607 22497
rect 6549 22488 6561 22491
rect 5040 22460 6561 22488
rect 4982 22448 4988 22451
rect 5040 22448 5046 22460
rect 6549 22457 6561 22460
rect 6595 22457 6607 22491
rect 6549 22451 6607 22457
rect 7006 22448 7012 22500
rect 7064 22488 7070 22500
rect 7064 22460 7109 22488
rect 7064 22448 7070 22460
rect 7190 22448 7196 22500
rect 7248 22488 7254 22500
rect 8404 22488 8432 22519
rect 8478 22516 8484 22528
rect 8536 22516 8542 22568
rect 8941 22559 8999 22565
rect 8941 22525 8953 22559
rect 8987 22556 8999 22559
rect 9582 22556 9588 22568
rect 8987 22528 9588 22556
rect 8987 22525 8999 22528
rect 8941 22519 8999 22525
rect 9582 22516 9588 22528
rect 9640 22516 9646 22568
rect 9858 22516 9864 22568
rect 9916 22556 9922 22568
rect 9953 22559 10011 22565
rect 9953 22556 9965 22559
rect 9916 22528 9965 22556
rect 9916 22516 9922 22528
rect 9953 22525 9965 22528
rect 9999 22525 10011 22559
rect 9953 22519 10011 22525
rect 10042 22516 10048 22568
rect 10100 22556 10106 22568
rect 10226 22556 10232 22568
rect 10100 22528 10145 22556
rect 10187 22528 10232 22556
rect 10100 22516 10106 22528
rect 10226 22516 10232 22528
rect 10284 22556 10290 22568
rect 10965 22559 11023 22565
rect 10965 22556 10977 22559
rect 10284 22528 10977 22556
rect 10284 22516 10290 22528
rect 10965 22525 10977 22528
rect 11011 22556 11023 22559
rect 12066 22556 12072 22568
rect 11011 22528 12072 22556
rect 11011 22525 11023 22528
rect 10965 22519 11023 22525
rect 12066 22516 12072 22528
rect 12124 22516 12130 22568
rect 12437 22559 12495 22565
rect 12437 22525 12449 22559
rect 12483 22556 12495 22559
rect 12526 22556 12532 22568
rect 12483 22528 12532 22556
rect 12483 22525 12495 22528
rect 12437 22519 12495 22525
rect 12526 22516 12532 22528
rect 12584 22556 12590 22568
rect 12897 22559 12955 22565
rect 12897 22556 12909 22559
rect 12584 22528 12909 22556
rect 12584 22516 12590 22528
rect 12897 22525 12909 22528
rect 12943 22525 12955 22559
rect 13446 22556 13452 22568
rect 13407 22528 13452 22556
rect 12897 22519 12955 22525
rect 13446 22516 13452 22528
rect 13504 22556 13510 22568
rect 13909 22559 13967 22565
rect 13909 22556 13921 22559
rect 13504 22528 13921 22556
rect 13504 22516 13510 22528
rect 13909 22525 13921 22528
rect 13955 22525 13967 22559
rect 13909 22519 13967 22525
rect 9122 22488 9128 22500
rect 7248 22460 8432 22488
rect 9083 22460 9128 22488
rect 7248 22448 7254 22460
rect 9122 22448 9128 22460
rect 9180 22448 9186 22500
rect 9398 22448 9404 22500
rect 9456 22488 9462 22500
rect 12618 22488 12624 22500
rect 9456 22460 12624 22488
rect 9456 22448 9462 22460
rect 12618 22448 12624 22460
rect 12676 22448 12682 22500
rect 9490 22420 9496 22432
rect 9451 22392 9496 22420
rect 9490 22380 9496 22392
rect 9548 22380 9554 22432
rect 9766 22420 9772 22432
rect 9727 22392 9772 22420
rect 9766 22380 9772 22392
rect 9824 22420 9830 22432
rect 10042 22420 10048 22432
rect 9824 22392 10048 22420
rect 9824 22380 9830 22392
rect 10042 22380 10048 22392
rect 10100 22380 10106 22432
rect 11514 22380 11520 22432
rect 11572 22420 11578 22432
rect 11701 22423 11759 22429
rect 11701 22420 11713 22423
rect 11572 22392 11713 22420
rect 11572 22380 11578 22392
rect 11701 22389 11713 22392
rect 11747 22389 11759 22423
rect 11701 22383 11759 22389
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 4338 22216 4344 22228
rect 4299 22188 4344 22216
rect 4338 22176 4344 22188
rect 4396 22176 4402 22228
rect 5442 22216 5448 22228
rect 5403 22188 5448 22216
rect 5442 22176 5448 22188
rect 5500 22176 5506 22228
rect 7466 22176 7472 22228
rect 7524 22216 7530 22228
rect 7653 22219 7711 22225
rect 7653 22216 7665 22219
rect 7524 22188 7665 22216
rect 7524 22176 7530 22188
rect 7653 22185 7665 22188
rect 7699 22185 7711 22219
rect 7653 22179 7711 22185
rect 9122 22176 9128 22228
rect 9180 22216 9186 22228
rect 9401 22219 9459 22225
rect 9401 22216 9413 22219
rect 9180 22188 9413 22216
rect 9180 22176 9186 22188
rect 9401 22185 9413 22188
rect 9447 22216 9459 22219
rect 10410 22216 10416 22228
rect 9447 22188 10088 22216
rect 10371 22188 10416 22216
rect 9447 22185 9459 22188
rect 9401 22179 9459 22185
rect 4887 22151 4945 22157
rect 4887 22117 4899 22151
rect 4933 22148 4945 22151
rect 4982 22148 4988 22160
rect 4933 22120 4988 22148
rect 4933 22117 4945 22120
rect 4887 22111 4945 22117
rect 4982 22108 4988 22120
rect 5040 22108 5046 22160
rect 6178 22108 6184 22160
rect 6236 22148 6242 22160
rect 6236 22120 6776 22148
rect 6236 22108 6242 22120
rect 5902 22040 5908 22092
rect 5960 22080 5966 22092
rect 6748 22089 6776 22120
rect 6273 22083 6331 22089
rect 6273 22080 6285 22083
rect 5960 22052 6285 22080
rect 5960 22040 5966 22052
rect 6273 22049 6285 22052
rect 6319 22049 6331 22083
rect 6273 22043 6331 22049
rect 6733 22083 6791 22089
rect 6733 22049 6745 22083
rect 6779 22049 6791 22083
rect 6733 22043 6791 22049
rect 8478 22040 8484 22092
rect 8536 22080 8542 22092
rect 8665 22083 8723 22089
rect 8665 22080 8677 22083
rect 8536 22052 8677 22080
rect 8536 22040 8542 22052
rect 8665 22049 8677 22052
rect 8711 22080 8723 22083
rect 9766 22080 9772 22092
rect 8711 22052 9772 22080
rect 8711 22049 8723 22052
rect 8665 22043 8723 22049
rect 9766 22040 9772 22052
rect 9824 22040 9830 22092
rect 10060 22089 10088 22188
rect 10410 22176 10416 22188
rect 10468 22176 10474 22228
rect 10965 22219 11023 22225
rect 10965 22185 10977 22219
rect 11011 22216 11023 22219
rect 11514 22216 11520 22228
rect 11011 22188 11520 22216
rect 11011 22185 11023 22188
rect 10965 22179 11023 22185
rect 11514 22176 11520 22188
rect 11572 22176 11578 22228
rect 12526 22148 12532 22160
rect 12487 22120 12532 22148
rect 12526 22108 12532 22120
rect 12584 22108 12590 22160
rect 10045 22083 10103 22089
rect 10045 22049 10057 22083
rect 10091 22049 10103 22083
rect 10045 22043 10103 22049
rect 11514 22040 11520 22092
rect 11572 22080 11578 22092
rect 11793 22083 11851 22089
rect 11793 22080 11805 22083
rect 11572 22052 11805 22080
rect 11572 22040 11578 22052
rect 11793 22049 11805 22052
rect 11839 22049 11851 22083
rect 12066 22080 12072 22092
rect 12027 22052 12072 22080
rect 11793 22043 11851 22049
rect 12066 22040 12072 22052
rect 12124 22040 12130 22092
rect 4522 22012 4528 22024
rect 4483 21984 4528 22012
rect 4522 21972 4528 21984
rect 4580 21972 4586 22024
rect 6822 22012 6828 22024
rect 6783 21984 6828 22012
rect 6822 21972 6828 21984
rect 6880 21972 6886 22024
rect 6914 21972 6920 22024
rect 6972 22012 6978 22024
rect 7377 22015 7435 22021
rect 7377 22012 7389 22015
rect 6972 21984 7389 22012
rect 6972 21972 6978 21984
rect 7377 21981 7389 21984
rect 7423 22012 7435 22015
rect 8754 22012 8760 22024
rect 7423 21984 8760 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 8754 21972 8760 21984
rect 8812 21972 8818 22024
rect 11885 21947 11943 21953
rect 11885 21913 11897 21947
rect 11931 21944 11943 21947
rect 12158 21944 12164 21956
rect 11931 21916 12164 21944
rect 11931 21913 11943 21916
rect 11885 21907 11943 21913
rect 12158 21904 12164 21916
rect 12216 21904 12222 21956
rect 9858 21876 9864 21888
rect 9819 21848 9864 21876
rect 9858 21836 9864 21848
rect 9916 21836 9922 21888
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 4982 21632 4988 21684
rect 5040 21672 5046 21684
rect 5261 21675 5319 21681
rect 5261 21672 5273 21675
rect 5040 21644 5273 21672
rect 5040 21632 5046 21644
rect 5261 21641 5273 21644
rect 5307 21672 5319 21675
rect 5626 21672 5632 21684
rect 5307 21644 5632 21672
rect 5307 21641 5319 21644
rect 5261 21635 5319 21641
rect 5626 21632 5632 21644
rect 5684 21632 5690 21684
rect 5902 21672 5908 21684
rect 5863 21644 5908 21672
rect 5902 21632 5908 21644
rect 5960 21632 5966 21684
rect 7929 21675 7987 21681
rect 7929 21641 7941 21675
rect 7975 21672 7987 21675
rect 8846 21672 8852 21684
rect 7975 21644 8852 21672
rect 7975 21641 7987 21644
rect 7929 21635 7987 21641
rect 6914 21604 6920 21616
rect 6875 21576 6920 21604
rect 6914 21564 6920 21576
rect 6972 21564 6978 21616
rect 7944 21604 7972 21635
rect 8846 21632 8852 21644
rect 8904 21632 8910 21684
rect 10410 21632 10416 21684
rect 10468 21672 10474 21684
rect 10965 21675 11023 21681
rect 10965 21672 10977 21675
rect 10468 21644 10977 21672
rect 10468 21632 10474 21644
rect 10965 21641 10977 21644
rect 11011 21641 11023 21675
rect 12618 21672 12624 21684
rect 12579 21644 12624 21672
rect 10965 21635 11023 21641
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 8478 21604 8484 21616
rect 7484 21576 7972 21604
rect 8439 21576 8484 21604
rect 4430 21536 4436 21548
rect 4172 21508 4436 21536
rect 4172 21477 4200 21508
rect 4430 21496 4436 21508
rect 4488 21496 4494 21548
rect 4798 21536 4804 21548
rect 4759 21508 4804 21536
rect 4798 21496 4804 21508
rect 4856 21496 4862 21548
rect 6273 21539 6331 21545
rect 6273 21505 6285 21539
rect 6319 21536 6331 21539
rect 6319 21508 7144 21536
rect 6319 21505 6331 21508
rect 6273 21499 6331 21505
rect 4157 21471 4215 21477
rect 4157 21437 4169 21471
rect 4203 21437 4215 21471
rect 4157 21431 4215 21437
rect 4338 21428 4344 21480
rect 4396 21468 4402 21480
rect 7116 21477 7144 21508
rect 4709 21471 4767 21477
rect 4709 21468 4721 21471
rect 4396 21440 4721 21468
rect 4396 21428 4402 21440
rect 4709 21437 4721 21440
rect 4755 21437 4767 21471
rect 4709 21431 4767 21437
rect 6825 21471 6883 21477
rect 6825 21437 6837 21471
rect 6871 21437 6883 21471
rect 6825 21431 6883 21437
rect 7101 21471 7159 21477
rect 7101 21437 7113 21471
rect 7147 21468 7159 21471
rect 7484 21468 7512 21576
rect 8478 21564 8484 21576
rect 8536 21564 8542 21616
rect 8754 21564 8760 21616
rect 8812 21604 8818 21616
rect 10045 21607 10103 21613
rect 10045 21604 10057 21607
rect 8812 21576 10057 21604
rect 8812 21564 8818 21576
rect 10045 21573 10057 21576
rect 10091 21604 10103 21607
rect 11333 21607 11391 21613
rect 11333 21604 11345 21607
rect 10091 21576 11345 21604
rect 10091 21573 10103 21576
rect 10045 21567 10103 21573
rect 11333 21573 11345 21576
rect 11379 21573 11391 21607
rect 11333 21567 11391 21573
rect 7561 21539 7619 21545
rect 7561 21505 7573 21539
rect 7607 21536 7619 21539
rect 9674 21536 9680 21548
rect 7607 21508 9680 21536
rect 7607 21505 7619 21508
rect 7561 21499 7619 21505
rect 9674 21496 9680 21508
rect 9732 21496 9738 21548
rect 8389 21471 8447 21477
rect 8389 21468 8401 21471
rect 7147 21440 7512 21468
rect 8312 21440 8401 21468
rect 7147 21437 7159 21440
rect 7101 21431 7159 21437
rect 3418 21360 3424 21412
rect 3476 21400 3482 21412
rect 4065 21403 4123 21409
rect 4065 21400 4077 21403
rect 3476 21372 4077 21400
rect 3476 21360 3482 21372
rect 4065 21369 4077 21372
rect 4111 21369 4123 21403
rect 4065 21363 4123 21369
rect 6641 21403 6699 21409
rect 6641 21369 6653 21403
rect 6687 21400 6699 21403
rect 6840 21400 6868 21431
rect 8312 21400 8340 21440
rect 8389 21437 8401 21440
rect 8435 21437 8447 21471
rect 8389 21431 8447 21437
rect 8665 21471 8723 21477
rect 8665 21437 8677 21471
rect 8711 21468 8723 21471
rect 8754 21468 8760 21480
rect 8711 21440 8760 21468
rect 8711 21437 8723 21440
rect 8665 21431 8723 21437
rect 8754 21428 8760 21440
rect 8812 21428 8818 21480
rect 9490 21428 9496 21480
rect 9548 21468 9554 21480
rect 9858 21468 9864 21480
rect 9548 21440 9864 21468
rect 9548 21428 9554 21440
rect 9858 21428 9864 21440
rect 9916 21468 9922 21480
rect 9953 21471 10011 21477
rect 9953 21468 9965 21471
rect 9916 21440 9965 21468
rect 9916 21428 9922 21440
rect 9953 21437 9965 21440
rect 9999 21437 10011 21471
rect 9953 21431 10011 21437
rect 10042 21428 10048 21480
rect 10100 21468 10106 21480
rect 10229 21471 10287 21477
rect 10229 21468 10241 21471
rect 10100 21440 10241 21468
rect 10100 21428 10106 21440
rect 10229 21437 10241 21440
rect 10275 21437 10287 21471
rect 10229 21431 10287 21437
rect 10689 21471 10747 21477
rect 10689 21437 10701 21471
rect 10735 21468 10747 21471
rect 12437 21471 12495 21477
rect 12437 21468 12449 21471
rect 10735 21440 12449 21468
rect 10735 21437 10747 21440
rect 10689 21431 10747 21437
rect 12437 21437 12449 21440
rect 12483 21468 12495 21471
rect 12897 21471 12955 21477
rect 12897 21468 12909 21471
rect 12483 21440 12909 21468
rect 12483 21437 12495 21440
rect 12437 21431 12495 21437
rect 12897 21437 12909 21440
rect 12943 21437 12955 21471
rect 12897 21431 12955 21437
rect 6687 21372 8340 21400
rect 6687 21369 6699 21372
rect 6641 21363 6699 21369
rect 8312 21344 8340 21372
rect 9125 21403 9183 21409
rect 9125 21369 9137 21403
rect 9171 21400 9183 21403
rect 13446 21400 13452 21412
rect 9171 21372 13452 21400
rect 9171 21369 9183 21372
rect 9125 21363 9183 21369
rect 13446 21360 13452 21372
rect 13504 21360 13510 21412
rect 3786 21332 3792 21344
rect 3747 21304 3792 21332
rect 3786 21292 3792 21304
rect 3844 21292 3850 21344
rect 8294 21332 8300 21344
rect 8255 21304 8300 21332
rect 8294 21292 8300 21304
rect 8352 21292 8358 21344
rect 9493 21335 9551 21341
rect 9493 21301 9505 21335
rect 9539 21332 9551 21335
rect 9674 21332 9680 21344
rect 9539 21304 9680 21332
rect 9539 21301 9551 21304
rect 9493 21295 9551 21301
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 9861 21335 9919 21341
rect 9861 21301 9873 21335
rect 9907 21332 9919 21335
rect 9950 21332 9956 21344
rect 9907 21304 9956 21332
rect 9907 21301 9919 21304
rect 9861 21295 9919 21301
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 10042 21292 10048 21344
rect 10100 21332 10106 21344
rect 11514 21332 11520 21344
rect 10100 21304 11520 21332
rect 10100 21292 10106 21304
rect 11514 21292 11520 21304
rect 11572 21332 11578 21344
rect 11793 21335 11851 21341
rect 11793 21332 11805 21335
rect 11572 21304 11805 21332
rect 11572 21292 11578 21304
rect 11793 21301 11805 21304
rect 11839 21301 11851 21335
rect 12158 21332 12164 21344
rect 12119 21304 12164 21332
rect 11793 21295 11851 21301
rect 12158 21292 12164 21304
rect 12216 21292 12222 21344
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 3786 21088 3792 21140
rect 3844 21128 3850 21140
rect 4249 21131 4307 21137
rect 4249 21128 4261 21131
rect 3844 21100 4261 21128
rect 3844 21088 3850 21100
rect 4249 21097 4261 21100
rect 4295 21128 4307 21131
rect 4522 21128 4528 21140
rect 4295 21100 4528 21128
rect 4295 21097 4307 21100
rect 4249 21091 4307 21097
rect 4522 21088 4528 21100
rect 4580 21088 4586 21140
rect 6178 21088 6184 21140
rect 6236 21128 6242 21140
rect 6273 21131 6331 21137
rect 6273 21128 6285 21131
rect 6236 21100 6285 21128
rect 6236 21088 6242 21100
rect 6273 21097 6285 21100
rect 6319 21097 6331 21131
rect 6273 21091 6331 21097
rect 8294 21088 8300 21140
rect 8352 21128 8358 21140
rect 10042 21128 10048 21140
rect 8352 21100 10048 21128
rect 8352 21088 8358 21100
rect 10042 21088 10048 21100
rect 10100 21088 10106 21140
rect 10137 21131 10195 21137
rect 10137 21097 10149 21131
rect 10183 21128 10195 21131
rect 10226 21128 10232 21140
rect 10183 21100 10232 21128
rect 10183 21097 10195 21100
rect 10137 21091 10195 21097
rect 10226 21088 10232 21100
rect 10284 21088 10290 21140
rect 10781 21131 10839 21137
rect 10781 21097 10793 21131
rect 10827 21128 10839 21131
rect 11146 21128 11152 21140
rect 10827 21100 11152 21128
rect 10827 21097 10839 21100
rect 10781 21091 10839 21097
rect 11146 21088 11152 21100
rect 11204 21088 11210 21140
rect 12066 21088 12072 21140
rect 12124 21128 12130 21140
rect 12253 21131 12311 21137
rect 12253 21128 12265 21131
rect 12124 21100 12265 21128
rect 12124 21088 12130 21100
rect 12253 21097 12265 21100
rect 12299 21097 12311 21131
rect 12253 21091 12311 21097
rect 4706 21060 4712 21072
rect 4264 21032 4712 21060
rect 4264 21001 4292 21032
rect 4706 21020 4712 21032
rect 4764 21060 4770 21072
rect 5902 21060 5908 21072
rect 4764 21032 5908 21060
rect 4764 21020 4770 21032
rect 5902 21020 5908 21032
rect 5960 21020 5966 21072
rect 6638 21020 6644 21072
rect 6696 21060 6702 21072
rect 6733 21063 6791 21069
rect 6733 21060 6745 21063
rect 6696 21032 6745 21060
rect 6696 21020 6702 21032
rect 6733 21029 6745 21032
rect 6779 21029 6791 21063
rect 6733 21023 6791 21029
rect 7285 21063 7343 21069
rect 7285 21029 7297 21063
rect 7331 21060 7343 21063
rect 7466 21060 7472 21072
rect 7331 21032 7472 21060
rect 7331 21029 7343 21032
rect 7285 21023 7343 21029
rect 7466 21020 7472 21032
rect 7524 21060 7530 21072
rect 8662 21060 8668 21072
rect 7524 21032 8668 21060
rect 7524 21020 7530 21032
rect 8662 21020 8668 21032
rect 8720 21020 8726 21072
rect 8754 21020 8760 21072
rect 8812 21060 8818 21072
rect 9950 21060 9956 21072
rect 8812 21032 9956 21060
rect 8812 21020 8818 21032
rect 9784 21004 9812 21032
rect 9950 21020 9956 21032
rect 10008 21060 10014 21072
rect 10008 21032 11560 21060
rect 10008 21020 10014 21032
rect 11532 21004 11560 21032
rect 4249 20995 4307 21001
rect 4249 20961 4261 20995
rect 4295 20961 4307 20995
rect 4249 20955 4307 20961
rect 4338 20952 4344 21004
rect 4396 20992 4402 21004
rect 4617 20995 4675 21001
rect 4617 20992 4629 20995
rect 4396 20964 4629 20992
rect 4396 20952 4402 20964
rect 4617 20961 4629 20964
rect 4663 20961 4675 20995
rect 4617 20955 4675 20961
rect 7558 20952 7564 21004
rect 7616 20992 7622 21004
rect 7834 20992 7840 21004
rect 7616 20964 7840 20992
rect 7616 20952 7622 20964
rect 7834 20952 7840 20964
rect 7892 20992 7898 21004
rect 8148 20995 8206 21001
rect 8148 20992 8160 20995
rect 7892 20964 8160 20992
rect 7892 20952 7898 20964
rect 8148 20961 8160 20964
rect 8194 20961 8206 20995
rect 9766 20992 9772 21004
rect 9679 20964 9772 20992
rect 8148 20955 8206 20961
rect 9766 20952 9772 20964
rect 9824 20952 9830 21004
rect 9858 20952 9864 21004
rect 9916 20992 9922 21004
rect 11238 20992 11244 21004
rect 9916 20964 11244 20992
rect 9916 20952 9922 20964
rect 11238 20952 11244 20964
rect 11296 20952 11302 21004
rect 11514 20992 11520 21004
rect 11475 20964 11520 20992
rect 11514 20952 11520 20964
rect 11572 20952 11578 21004
rect 3970 20884 3976 20936
rect 4028 20924 4034 20936
rect 4356 20924 4384 20952
rect 4028 20896 4384 20924
rect 4028 20884 4034 20896
rect 6270 20884 6276 20936
rect 6328 20924 6334 20936
rect 6641 20927 6699 20933
rect 6641 20924 6653 20927
rect 6328 20896 6653 20924
rect 6328 20884 6334 20896
rect 6641 20893 6653 20896
rect 6687 20924 6699 20927
rect 8251 20927 8309 20933
rect 8251 20924 8263 20927
rect 6687 20896 8263 20924
rect 6687 20893 6699 20896
rect 6641 20887 6699 20893
rect 8251 20893 8263 20896
rect 8297 20893 8309 20927
rect 8251 20887 8309 20893
rect 8386 20884 8392 20936
rect 8444 20924 8450 20936
rect 11701 20927 11759 20933
rect 11701 20924 11713 20927
rect 8444 20896 11713 20924
rect 8444 20884 8450 20896
rect 11701 20893 11713 20896
rect 11747 20893 11759 20927
rect 11701 20887 11759 20893
rect 4338 20816 4344 20868
rect 4396 20856 4402 20868
rect 7742 20856 7748 20868
rect 4396 20828 7748 20856
rect 4396 20816 4402 20828
rect 7742 20816 7748 20828
rect 7800 20856 7806 20868
rect 8018 20856 8024 20868
rect 7800 20828 8024 20856
rect 7800 20816 7806 20828
rect 8018 20816 8024 20828
rect 8076 20816 8082 20868
rect 8665 20859 8723 20865
rect 8665 20825 8677 20859
rect 8711 20856 8723 20859
rect 9674 20856 9680 20868
rect 8711 20828 9680 20856
rect 8711 20825 8723 20828
rect 8665 20819 8723 20825
rect 9674 20816 9680 20828
rect 9732 20856 9738 20868
rect 11333 20859 11391 20865
rect 11333 20856 11345 20859
rect 9732 20828 11345 20856
rect 9732 20816 9738 20828
rect 11333 20825 11345 20828
rect 11379 20856 11391 20859
rect 12066 20856 12072 20868
rect 11379 20828 12072 20856
rect 11379 20825 11391 20828
rect 11333 20819 11391 20825
rect 12066 20816 12072 20828
rect 12124 20816 12130 20868
rect 6730 20748 6736 20800
rect 6788 20788 6794 20800
rect 7561 20791 7619 20797
rect 7561 20788 7573 20791
rect 6788 20760 7573 20788
rect 6788 20748 6794 20760
rect 7561 20757 7573 20760
rect 7607 20757 7619 20791
rect 7561 20751 7619 20757
rect 9493 20791 9551 20797
rect 9493 20757 9505 20791
rect 9539 20788 9551 20791
rect 9950 20788 9956 20800
rect 9539 20760 9956 20788
rect 9539 20757 9551 20760
rect 9493 20751 9551 20757
rect 9950 20748 9956 20760
rect 10008 20748 10014 20800
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 3510 20544 3516 20596
rect 3568 20584 3574 20596
rect 3605 20587 3663 20593
rect 3605 20584 3617 20587
rect 3568 20556 3617 20584
rect 3568 20544 3574 20556
rect 3605 20553 3617 20556
rect 3651 20584 3663 20587
rect 3970 20584 3976 20596
rect 3651 20556 3976 20584
rect 3651 20553 3663 20556
rect 3605 20547 3663 20553
rect 3970 20544 3976 20556
rect 4028 20544 4034 20596
rect 4617 20587 4675 20593
rect 4617 20553 4629 20587
rect 4663 20584 4675 20587
rect 4706 20584 4712 20596
rect 4663 20556 4712 20584
rect 4663 20553 4675 20556
rect 4617 20547 4675 20553
rect 3835 20451 3893 20457
rect 3835 20417 3847 20451
rect 3881 20448 3893 20451
rect 4522 20448 4528 20460
rect 3881 20420 4528 20448
rect 3881 20417 3893 20420
rect 3835 20411 3893 20417
rect 4522 20408 4528 20420
rect 4580 20408 4586 20460
rect 3748 20383 3806 20389
rect 3748 20349 3760 20383
rect 3794 20349 3806 20383
rect 3748 20343 3806 20349
rect 3763 20244 3791 20343
rect 4062 20272 4068 20324
rect 4120 20312 4126 20324
rect 4632 20312 4660 20547
rect 4706 20544 4712 20556
rect 4764 20544 4770 20596
rect 6270 20584 6276 20596
rect 6231 20556 6276 20584
rect 6270 20544 6276 20556
rect 6328 20544 6334 20596
rect 9766 20584 9772 20596
rect 9727 20556 9772 20584
rect 9766 20544 9772 20556
rect 9824 20544 9830 20596
rect 11238 20544 11244 20596
rect 11296 20584 11302 20596
rect 11977 20587 12035 20593
rect 11977 20584 11989 20587
rect 11296 20556 11989 20584
rect 11296 20544 11302 20556
rect 11977 20553 11989 20556
rect 12023 20553 12035 20587
rect 11977 20547 12035 20553
rect 7466 20516 7472 20528
rect 7427 20488 7472 20516
rect 7466 20476 7472 20488
rect 7524 20476 7530 20528
rect 9490 20476 9496 20528
rect 9548 20516 9554 20528
rect 10045 20519 10103 20525
rect 10045 20516 10057 20519
rect 9548 20488 10057 20516
rect 9548 20476 9554 20488
rect 10045 20485 10057 20488
rect 10091 20516 10103 20519
rect 11054 20516 11060 20528
rect 10091 20488 11060 20516
rect 10091 20485 10103 20488
rect 10045 20479 10103 20485
rect 11054 20476 11060 20488
rect 11112 20516 11118 20528
rect 14734 20516 14740 20528
rect 11112 20488 14740 20516
rect 11112 20476 11118 20488
rect 14734 20476 14740 20488
rect 14792 20476 14798 20528
rect 5445 20451 5503 20457
rect 5445 20417 5457 20451
rect 5491 20448 5503 20451
rect 5534 20448 5540 20460
rect 5491 20420 5540 20448
rect 5491 20417 5503 20420
rect 5445 20411 5503 20417
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 5994 20408 6000 20460
rect 6052 20448 6058 20460
rect 7834 20448 7840 20460
rect 6052 20420 7840 20448
rect 6052 20408 6058 20420
rect 7834 20408 7840 20420
rect 7892 20408 7898 20460
rect 8478 20408 8484 20460
rect 8536 20448 8542 20460
rect 9125 20451 9183 20457
rect 9125 20448 9137 20451
rect 8536 20420 9137 20448
rect 8536 20408 8542 20420
rect 9125 20417 9137 20420
rect 9171 20448 9183 20451
rect 9398 20448 9404 20460
rect 9171 20420 9404 20448
rect 9171 20417 9183 20420
rect 9125 20411 9183 20417
rect 9398 20408 9404 20420
rect 9456 20408 9462 20460
rect 8294 20380 8300 20392
rect 8207 20352 8300 20380
rect 8294 20340 8300 20352
rect 8352 20380 8358 20392
rect 8754 20380 8760 20392
rect 8352 20352 8760 20380
rect 8352 20340 8358 20352
rect 8754 20340 8760 20352
rect 8812 20340 8818 20392
rect 9950 20380 9956 20392
rect 9911 20352 9956 20380
rect 9950 20340 9956 20352
rect 10008 20340 10014 20392
rect 10134 20340 10140 20392
rect 10192 20380 10198 20392
rect 10229 20383 10287 20389
rect 10229 20380 10241 20383
rect 10192 20352 10241 20380
rect 10192 20340 10198 20352
rect 10229 20349 10241 20352
rect 10275 20380 10287 20383
rect 11146 20380 11152 20392
rect 10275 20352 11152 20380
rect 10275 20349 10287 20352
rect 10229 20343 10287 20349
rect 11146 20340 11152 20352
rect 11204 20340 11210 20392
rect 4798 20312 4804 20324
rect 4120 20284 4660 20312
rect 4759 20284 4804 20312
rect 4120 20272 4126 20284
rect 4798 20272 4804 20284
rect 4856 20272 4862 20324
rect 4890 20272 4896 20324
rect 4948 20312 4954 20324
rect 4948 20284 4993 20312
rect 4948 20272 4954 20284
rect 6730 20272 6736 20324
rect 6788 20312 6794 20324
rect 6917 20315 6975 20321
rect 6917 20312 6929 20315
rect 6788 20284 6929 20312
rect 6788 20272 6794 20284
rect 6917 20281 6929 20284
rect 6963 20281 6975 20315
rect 6917 20275 6975 20281
rect 7006 20272 7012 20324
rect 7064 20312 7070 20324
rect 10686 20312 10692 20324
rect 7064 20284 7109 20312
rect 10647 20284 10692 20312
rect 7064 20272 7070 20284
rect 10686 20272 10692 20284
rect 10744 20272 10750 20324
rect 11333 20315 11391 20321
rect 11333 20281 11345 20315
rect 11379 20312 11391 20315
rect 11514 20312 11520 20324
rect 11379 20284 11520 20312
rect 11379 20281 11391 20284
rect 11333 20275 11391 20281
rect 11514 20272 11520 20284
rect 11572 20312 11578 20324
rect 12250 20312 12256 20324
rect 11572 20284 12256 20312
rect 11572 20272 11578 20284
rect 12250 20272 12256 20284
rect 12308 20272 12314 20324
rect 4246 20244 4252 20256
rect 3763 20216 4252 20244
rect 4246 20204 4252 20216
rect 4304 20244 4310 20256
rect 5074 20244 5080 20256
rect 4304 20216 5080 20244
rect 4304 20204 4310 20216
rect 5074 20204 5080 20216
rect 5132 20204 5138 20256
rect 6638 20244 6644 20256
rect 6599 20216 6644 20244
rect 6638 20204 6644 20216
rect 6696 20204 6702 20256
rect 11701 20247 11759 20253
rect 11701 20213 11713 20247
rect 11747 20244 11759 20247
rect 12066 20244 12072 20256
rect 11747 20216 12072 20244
rect 11747 20213 11759 20216
rect 11701 20207 11759 20213
rect 12066 20204 12072 20216
rect 12124 20204 12130 20256
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 4798 20040 4804 20052
rect 4126 20012 4804 20040
rect 2961 19975 3019 19981
rect 2961 19941 2973 19975
rect 3007 19972 3019 19975
rect 4126 19972 4154 20012
rect 4798 20000 4804 20012
rect 4856 20000 4862 20052
rect 4890 20000 4896 20052
rect 4948 20040 4954 20052
rect 5077 20043 5135 20049
rect 5077 20040 5089 20043
rect 4948 20012 5089 20040
rect 4948 20000 4954 20012
rect 5077 20009 5089 20012
rect 5123 20009 5135 20043
rect 5077 20003 5135 20009
rect 6457 20043 6515 20049
rect 6457 20009 6469 20043
rect 6503 20009 6515 20043
rect 9490 20040 9496 20052
rect 9451 20012 9496 20040
rect 6457 20003 6515 20009
rect 5534 19972 5540 19984
rect 3007 19944 4154 19972
rect 4310 19944 5540 19972
rect 3007 19941 3019 19944
rect 2961 19935 3019 19941
rect 3970 19864 3976 19916
rect 4028 19904 4034 19916
rect 4310 19913 4338 19944
rect 5534 19932 5540 19944
rect 5592 19932 5598 19984
rect 5626 19932 5632 19984
rect 5684 19972 5690 19984
rect 5902 19981 5908 19984
rect 5858 19975 5908 19981
rect 5858 19972 5870 19975
rect 5684 19944 5870 19972
rect 5684 19932 5690 19944
rect 5858 19941 5870 19944
rect 5904 19941 5908 19975
rect 5858 19935 5908 19941
rect 5902 19932 5908 19935
rect 5960 19932 5966 19984
rect 6472 19972 6500 20003
rect 9490 20000 9496 20012
rect 9548 20000 9554 20052
rect 9582 20000 9588 20052
rect 9640 20040 9646 20052
rect 11609 20043 11667 20049
rect 11609 20040 11621 20043
rect 9640 20012 11621 20040
rect 9640 20000 9646 20012
rect 11609 20009 11621 20012
rect 11655 20009 11667 20043
rect 11609 20003 11667 20009
rect 6638 19972 6644 19984
rect 6472 19944 6644 19972
rect 6638 19932 6644 19944
rect 6696 19972 6702 19984
rect 7469 19975 7527 19981
rect 7469 19972 7481 19975
rect 6696 19944 7481 19972
rect 6696 19932 6702 19944
rect 7469 19941 7481 19944
rect 7515 19972 7527 19975
rect 7834 19972 7840 19984
rect 7515 19944 7840 19972
rect 7515 19941 7527 19944
rect 7469 19935 7527 19941
rect 7834 19932 7840 19944
rect 7892 19932 7898 19984
rect 10597 19975 10655 19981
rect 10597 19941 10609 19975
rect 10643 19972 10655 19975
rect 10962 19972 10968 19984
rect 10643 19944 10968 19972
rect 10643 19941 10655 19944
rect 10597 19935 10655 19941
rect 10962 19932 10968 19944
rect 11020 19932 11026 19984
rect 4295 19907 4353 19913
rect 4295 19904 4307 19907
rect 4028 19876 4307 19904
rect 4028 19864 4034 19876
rect 4295 19873 4307 19876
rect 4341 19873 4353 19907
rect 4295 19867 4353 19873
rect 4522 19864 4528 19916
rect 4580 19904 4586 19916
rect 9861 19907 9919 19913
rect 4580 19876 7189 19904
rect 4580 19864 4586 19876
rect 4154 19796 4160 19848
rect 4212 19836 4218 19848
rect 4387 19839 4445 19845
rect 4387 19836 4399 19839
rect 4212 19808 4399 19836
rect 4212 19796 4218 19808
rect 4387 19805 4399 19808
rect 4433 19805 4445 19839
rect 5534 19836 5540 19848
rect 5495 19808 5540 19836
rect 4387 19799 4445 19805
rect 5534 19796 5540 19808
rect 5592 19796 5598 19848
rect 7161 19836 7189 19876
rect 9861 19873 9873 19907
rect 9907 19904 9919 19907
rect 9950 19904 9956 19916
rect 9907 19876 9956 19904
rect 9907 19873 9919 19876
rect 9861 19867 9919 19873
rect 7377 19839 7435 19845
rect 7377 19836 7389 19839
rect 7161 19808 7389 19836
rect 7377 19805 7389 19808
rect 7423 19836 7435 19839
rect 8294 19836 8300 19848
rect 7423 19808 8300 19836
rect 7423 19805 7435 19808
rect 7377 19799 7435 19805
rect 8294 19796 8300 19808
rect 8352 19796 8358 19848
rect 9876 19836 9904 19867
rect 9950 19864 9956 19876
rect 10008 19864 10014 19916
rect 10134 19904 10140 19916
rect 10095 19876 10140 19904
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 10686 19864 10692 19916
rect 10744 19904 10750 19916
rect 11425 19907 11483 19913
rect 11425 19904 11437 19907
rect 10744 19876 11437 19904
rect 10744 19864 10750 19876
rect 11425 19873 11437 19876
rect 11471 19904 11483 19907
rect 11514 19904 11520 19916
rect 11471 19876 11520 19904
rect 11471 19873 11483 19876
rect 11425 19867 11483 19873
rect 11514 19864 11520 19876
rect 11572 19864 11578 19916
rect 10594 19836 10600 19848
rect 9876 19808 10600 19836
rect 10594 19796 10600 19808
rect 10652 19796 10658 19848
rect 7926 19768 7932 19780
rect 7887 19740 7932 19768
rect 7926 19728 7932 19740
rect 7984 19728 7990 19780
rect 9950 19768 9956 19780
rect 9911 19740 9956 19768
rect 9950 19728 9956 19740
rect 10008 19728 10014 19780
rect 6914 19700 6920 19712
rect 6875 19672 6920 19700
rect 6914 19660 6920 19672
rect 6972 19660 6978 19712
rect 7374 19660 7380 19712
rect 7432 19700 7438 19712
rect 8297 19703 8355 19709
rect 8297 19700 8309 19703
rect 7432 19672 8309 19700
rect 7432 19660 7438 19672
rect 8297 19669 8309 19672
rect 8343 19669 8355 19703
rect 8297 19663 8355 19669
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 3789 19499 3847 19505
rect 3789 19465 3801 19499
rect 3835 19496 3847 19499
rect 3970 19496 3976 19508
rect 3835 19468 3976 19496
rect 3835 19465 3847 19468
rect 3789 19459 3847 19465
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 4890 19456 4896 19508
rect 4948 19496 4954 19508
rect 5169 19499 5227 19505
rect 5169 19496 5181 19499
rect 4948 19468 5181 19496
rect 4948 19456 4954 19468
rect 5169 19465 5181 19468
rect 5215 19465 5227 19499
rect 7834 19496 7840 19508
rect 7795 19468 7840 19496
rect 5169 19459 5227 19465
rect 7834 19456 7840 19468
rect 7892 19456 7898 19508
rect 9677 19499 9735 19505
rect 9677 19465 9689 19499
rect 9723 19496 9735 19499
rect 10134 19496 10140 19508
rect 9723 19468 10140 19496
rect 9723 19465 9735 19468
rect 9677 19459 9735 19465
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 10597 19499 10655 19505
rect 10597 19465 10609 19499
rect 10643 19496 10655 19499
rect 10873 19499 10931 19505
rect 10873 19496 10885 19499
rect 10643 19468 10885 19496
rect 10643 19465 10655 19468
rect 10597 19459 10655 19465
rect 10873 19465 10885 19468
rect 10919 19496 10931 19499
rect 11054 19496 11060 19508
rect 10919 19468 11060 19496
rect 10919 19465 10931 19468
rect 10873 19459 10931 19465
rect 11054 19456 11060 19468
rect 11112 19456 11118 19508
rect 11514 19496 11520 19508
rect 11475 19468 11520 19496
rect 11514 19456 11520 19468
rect 11572 19456 11578 19508
rect 3326 19388 3332 19440
rect 3384 19428 3390 19440
rect 6730 19428 6736 19440
rect 3384 19400 6736 19428
rect 3384 19388 3390 19400
rect 6730 19388 6736 19400
rect 6788 19388 6794 19440
rect 9309 19431 9367 19437
rect 9309 19428 9321 19431
rect 8588 19400 9321 19428
rect 4065 19363 4123 19369
rect 4065 19329 4077 19363
rect 4111 19360 4123 19363
rect 4522 19360 4528 19372
rect 4111 19332 4528 19360
rect 4111 19329 4123 19332
rect 4065 19323 4123 19329
rect 4522 19320 4528 19332
rect 4580 19320 4586 19372
rect 7374 19360 7380 19372
rect 6748 19332 7380 19360
rect 2685 19295 2743 19301
rect 2685 19261 2697 19295
rect 2731 19261 2743 19295
rect 2685 19255 2743 19261
rect 3237 19295 3295 19301
rect 3237 19261 3249 19295
rect 3283 19292 3295 19295
rect 3510 19292 3516 19304
rect 3283 19264 3516 19292
rect 3283 19261 3295 19264
rect 3237 19255 3295 19261
rect 2406 19116 2412 19168
rect 2464 19156 2470 19168
rect 2501 19159 2559 19165
rect 2501 19156 2513 19159
rect 2464 19128 2513 19156
rect 2464 19116 2470 19128
rect 2501 19125 2513 19128
rect 2547 19156 2559 19159
rect 2700 19156 2728 19255
rect 3510 19252 3516 19264
rect 3568 19252 3574 19304
rect 4246 19292 4252 19304
rect 4207 19264 4252 19292
rect 4246 19252 4252 19264
rect 4304 19252 4310 19304
rect 5534 19292 5540 19304
rect 4448 19264 5540 19292
rect 3421 19227 3479 19233
rect 3421 19193 3433 19227
rect 3467 19224 3479 19227
rect 4448 19224 4476 19264
rect 5534 19252 5540 19264
rect 5592 19292 5598 19304
rect 5905 19295 5963 19301
rect 5905 19292 5917 19295
rect 5592 19264 5917 19292
rect 5592 19252 5598 19264
rect 5905 19261 5917 19264
rect 5951 19261 5963 19295
rect 5905 19255 5963 19261
rect 3467 19196 4476 19224
rect 3467 19193 3479 19196
rect 3421 19187 3479 19193
rect 5626 19184 5632 19236
rect 5684 19224 5690 19236
rect 6748 19224 6776 19332
rect 7374 19320 7380 19332
rect 7432 19320 7438 19372
rect 7561 19363 7619 19369
rect 7561 19329 7573 19363
rect 7607 19360 7619 19363
rect 7926 19360 7932 19372
rect 7607 19332 7932 19360
rect 7607 19329 7619 19332
rect 7561 19323 7619 19329
rect 7926 19320 7932 19332
rect 7984 19320 7990 19372
rect 8588 19301 8616 19400
rect 9309 19397 9321 19400
rect 9355 19428 9367 19431
rect 11422 19428 11428 19440
rect 9355 19400 11428 19428
rect 9355 19397 9367 19400
rect 9309 19391 9367 19397
rect 11422 19388 11428 19400
rect 11480 19388 11486 19440
rect 8941 19363 8999 19369
rect 8941 19329 8953 19363
rect 8987 19360 8999 19363
rect 12434 19360 12440 19372
rect 8987 19332 12440 19360
rect 8987 19329 8999 19332
rect 8941 19323 8999 19329
rect 12434 19320 12440 19332
rect 12492 19320 12498 19372
rect 8573 19295 8631 19301
rect 8573 19261 8585 19295
rect 8619 19261 8631 19295
rect 8573 19255 8631 19261
rect 9766 19252 9772 19304
rect 9824 19292 9830 19304
rect 10413 19295 10471 19301
rect 10413 19292 10425 19295
rect 9824 19264 10425 19292
rect 9824 19252 9830 19264
rect 10413 19261 10425 19264
rect 10459 19292 10471 19295
rect 10597 19295 10655 19301
rect 10597 19292 10609 19295
rect 10459 19264 10609 19292
rect 10459 19261 10471 19264
rect 10413 19255 10471 19261
rect 10597 19261 10609 19264
rect 10643 19261 10655 19295
rect 10597 19255 10655 19261
rect 6917 19227 6975 19233
rect 6917 19224 6929 19227
rect 5684 19196 6929 19224
rect 5684 19184 5690 19196
rect 6917 19193 6929 19196
rect 6963 19193 6975 19227
rect 6917 19187 6975 19193
rect 7009 19227 7067 19233
rect 7009 19193 7021 19227
rect 7055 19193 7067 19227
rect 7009 19187 7067 19193
rect 2547 19128 2728 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 4522 19116 4528 19168
rect 4580 19156 4586 19168
rect 4617 19159 4675 19165
rect 4617 19156 4629 19159
rect 4580 19128 4629 19156
rect 4580 19116 4586 19128
rect 4617 19125 4629 19128
rect 4663 19156 4675 19159
rect 5537 19159 5595 19165
rect 5537 19156 5549 19159
rect 4663 19128 5549 19156
rect 4663 19125 4675 19128
rect 4617 19119 4675 19125
rect 5537 19125 5549 19128
rect 5583 19156 5595 19159
rect 5902 19156 5908 19168
rect 5583 19128 5908 19156
rect 5583 19125 5595 19128
rect 5537 19119 5595 19125
rect 5902 19116 5908 19128
rect 5960 19116 5966 19168
rect 6638 19156 6644 19168
rect 6551 19128 6644 19156
rect 6638 19116 6644 19128
rect 6696 19156 6702 19168
rect 7024 19156 7052 19187
rect 7650 19184 7656 19236
rect 7708 19224 7714 19236
rect 8297 19227 8355 19233
rect 8297 19224 8309 19227
rect 7708 19196 8309 19224
rect 7708 19184 7714 19196
rect 8297 19193 8309 19196
rect 8343 19224 8355 19227
rect 8389 19227 8447 19233
rect 8389 19224 8401 19227
rect 8343 19196 8401 19224
rect 8343 19193 8355 19196
rect 8297 19187 8355 19193
rect 8389 19193 8401 19196
rect 8435 19193 8447 19227
rect 8389 19187 8447 19193
rect 9950 19184 9956 19236
rect 10008 19224 10014 19236
rect 10505 19227 10563 19233
rect 10505 19224 10517 19227
rect 10008 19196 10517 19224
rect 10008 19184 10014 19196
rect 10505 19193 10517 19196
rect 10551 19224 10563 19227
rect 11149 19227 11207 19233
rect 11149 19224 11161 19227
rect 10551 19196 11161 19224
rect 10551 19193 10563 19196
rect 10505 19187 10563 19193
rect 11149 19193 11161 19196
rect 11195 19193 11207 19227
rect 11149 19187 11207 19193
rect 6696 19128 7052 19156
rect 6696 19116 6702 19128
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 3237 18955 3295 18961
rect 3237 18921 3249 18955
rect 3283 18952 3295 18955
rect 3326 18952 3332 18964
rect 3283 18924 3332 18952
rect 3283 18921 3295 18924
rect 3237 18915 3295 18921
rect 3326 18912 3332 18924
rect 3384 18912 3390 18964
rect 3510 18912 3516 18964
rect 3568 18952 3574 18964
rect 4246 18952 4252 18964
rect 3568 18924 4154 18952
rect 4207 18924 4252 18952
rect 3568 18912 3574 18924
rect 2774 18884 2780 18896
rect 2687 18856 2780 18884
rect 2774 18844 2780 18856
rect 2832 18884 2838 18896
rect 3528 18884 3556 18912
rect 2832 18856 3556 18884
rect 4126 18884 4154 18924
rect 4246 18912 4252 18924
rect 4304 18912 4310 18964
rect 5445 18955 5503 18961
rect 5445 18952 5457 18955
rect 4626 18924 5457 18952
rect 4626 18884 4654 18924
rect 5445 18921 5457 18924
rect 5491 18952 5503 18955
rect 5534 18952 5540 18964
rect 5491 18924 5540 18952
rect 5491 18921 5503 18924
rect 5445 18915 5503 18921
rect 5534 18912 5540 18924
rect 5592 18952 5598 18964
rect 6178 18952 6184 18964
rect 5592 18924 6184 18952
rect 5592 18912 5598 18924
rect 6178 18912 6184 18924
rect 6236 18912 6242 18964
rect 6457 18955 6515 18961
rect 6457 18921 6469 18955
rect 6503 18921 6515 18955
rect 8294 18952 8300 18964
rect 8255 18924 8300 18952
rect 6457 18915 6515 18921
rect 4126 18856 4654 18884
rect 2832 18844 2838 18856
rect 5166 18844 5172 18896
rect 5224 18884 5230 18896
rect 5718 18884 5724 18896
rect 5224 18856 5724 18884
rect 5224 18844 5230 18856
rect 5718 18844 5724 18856
rect 5776 18844 5782 18896
rect 5902 18893 5908 18896
rect 5899 18884 5908 18893
rect 5863 18856 5908 18884
rect 5899 18847 5908 18856
rect 5902 18844 5908 18847
rect 5960 18844 5966 18896
rect 6472 18884 6500 18915
rect 8294 18912 8300 18924
rect 8352 18912 8358 18964
rect 9401 18955 9459 18961
rect 9401 18921 9413 18955
rect 9447 18952 9459 18955
rect 9582 18952 9588 18964
rect 9447 18924 9588 18952
rect 9447 18921 9459 18924
rect 9401 18915 9459 18921
rect 9582 18912 9588 18924
rect 9640 18952 9646 18964
rect 9950 18952 9956 18964
rect 9640 18924 9956 18952
rect 9640 18912 9646 18924
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 10594 18912 10600 18964
rect 10652 18952 10658 18964
rect 10689 18955 10747 18961
rect 10689 18952 10701 18955
rect 10652 18924 10701 18952
rect 10652 18912 10658 18924
rect 10689 18921 10701 18924
rect 10735 18921 10747 18955
rect 10689 18915 10747 18921
rect 6914 18884 6920 18896
rect 6472 18856 6920 18884
rect 6914 18844 6920 18856
rect 6972 18884 6978 18896
rect 7469 18887 7527 18893
rect 7469 18884 7481 18887
rect 6972 18856 7481 18884
rect 6972 18844 6978 18856
rect 7469 18853 7481 18856
rect 7515 18884 7527 18887
rect 8018 18884 8024 18896
rect 7515 18856 8024 18884
rect 7515 18853 7527 18856
rect 7469 18847 7527 18853
rect 8018 18844 8024 18856
rect 8076 18844 8082 18896
rect 1949 18819 2007 18825
rect 1949 18785 1961 18819
rect 1995 18816 2007 18819
rect 2038 18816 2044 18828
rect 1995 18788 2044 18816
rect 1995 18785 2007 18788
rect 1949 18779 2007 18785
rect 2038 18776 2044 18788
rect 2096 18776 2102 18828
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18816 2927 18819
rect 2958 18816 2964 18828
rect 2915 18788 2964 18816
rect 2915 18785 2927 18788
rect 2869 18779 2927 18785
rect 2958 18776 2964 18788
rect 3016 18776 3022 18828
rect 4592 18819 4650 18825
rect 4592 18785 4604 18819
rect 4638 18816 4650 18819
rect 4706 18816 4712 18828
rect 4638 18788 4712 18816
rect 4638 18785 4650 18788
rect 4592 18779 4650 18785
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 7190 18816 7196 18828
rect 5460 18788 7196 18816
rect 3326 18708 3332 18760
rect 3384 18748 3390 18760
rect 3513 18751 3571 18757
rect 3513 18748 3525 18751
rect 3384 18720 3525 18748
rect 3384 18708 3390 18720
rect 3513 18717 3525 18720
rect 3559 18748 3571 18751
rect 5460 18748 5488 18788
rect 7190 18776 7196 18788
rect 7248 18776 7254 18828
rect 9033 18819 9091 18825
rect 9033 18785 9045 18819
rect 9079 18816 9091 18819
rect 9665 18819 9723 18825
rect 9665 18816 9677 18819
rect 9079 18788 9677 18816
rect 9079 18785 9091 18788
rect 9033 18779 9091 18785
rect 9646 18785 9677 18788
rect 9711 18785 9723 18819
rect 9646 18779 9723 18785
rect 9953 18819 10011 18825
rect 9953 18785 9965 18819
rect 9999 18816 10011 18819
rect 10134 18816 10140 18828
rect 9999 18788 10140 18816
rect 9999 18785 10011 18788
rect 9953 18779 10011 18785
rect 3559 18720 5488 18748
rect 5537 18751 5595 18757
rect 3559 18717 3571 18720
rect 3513 18711 3571 18717
rect 5537 18717 5549 18751
rect 5583 18748 5595 18751
rect 5718 18748 5724 18760
rect 5583 18720 5724 18748
rect 5583 18717 5595 18720
rect 5537 18711 5595 18717
rect 5718 18708 5724 18720
rect 5776 18708 5782 18760
rect 7374 18748 7380 18760
rect 7335 18720 7380 18748
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 9646 18692 9674 18779
rect 10134 18776 10140 18788
rect 10192 18776 10198 18828
rect 11422 18776 11428 18828
rect 11480 18816 11486 18828
rect 11885 18819 11943 18825
rect 11885 18816 11897 18819
rect 11480 18788 11897 18816
rect 11480 18776 11486 18788
rect 11885 18785 11897 18788
rect 11931 18816 11943 18819
rect 13078 18816 13084 18828
rect 11931 18788 13084 18816
rect 11931 18785 11943 18788
rect 11885 18779 11943 18785
rect 13078 18776 13084 18788
rect 13136 18776 13142 18828
rect 9766 18748 9772 18760
rect 9727 18720 9772 18748
rect 9766 18708 9772 18720
rect 9824 18708 9830 18760
rect 10410 18748 10416 18760
rect 10371 18720 10416 18748
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 10686 18708 10692 18760
rect 10744 18748 10750 18760
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 10744 18720 11253 18748
rect 10744 18708 10750 18720
rect 11241 18717 11253 18720
rect 11287 18717 11299 18751
rect 11241 18711 11299 18717
rect 4663 18683 4721 18689
rect 4663 18649 4675 18683
rect 4709 18680 4721 18683
rect 6730 18680 6736 18692
rect 4709 18652 6736 18680
rect 4709 18649 4721 18652
rect 4663 18643 4721 18649
rect 6730 18640 6736 18652
rect 6788 18640 6794 18692
rect 7926 18680 7932 18692
rect 7887 18652 7932 18680
rect 7926 18640 7932 18652
rect 7984 18640 7990 18692
rect 9646 18652 9680 18692
rect 9674 18640 9680 18652
rect 9732 18640 9738 18692
rect 10226 18640 10232 18692
rect 10284 18680 10290 18692
rect 10778 18680 10784 18692
rect 10284 18652 10784 18680
rect 10284 18640 10290 18652
rect 10778 18640 10784 18652
rect 10836 18640 10842 18692
rect 2087 18615 2145 18621
rect 2087 18581 2099 18615
rect 2133 18612 2145 18615
rect 2590 18612 2596 18624
rect 2133 18584 2596 18612
rect 2133 18581 2145 18584
rect 2087 18575 2145 18581
rect 2590 18572 2596 18584
rect 2648 18572 2654 18624
rect 4982 18612 4988 18624
rect 4943 18584 4988 18612
rect 4982 18572 4988 18584
rect 5040 18572 5046 18624
rect 6822 18612 6828 18624
rect 6783 18584 6828 18612
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 2038 18408 2044 18420
rect 1951 18380 2044 18408
rect 2038 18368 2044 18380
rect 2096 18408 2102 18420
rect 4338 18408 4344 18420
rect 2096 18380 4344 18408
rect 2096 18368 2102 18380
rect 4338 18368 4344 18380
rect 4396 18368 4402 18420
rect 4617 18411 4675 18417
rect 4617 18377 4629 18411
rect 4663 18408 4675 18411
rect 4706 18408 4712 18420
rect 4663 18380 4712 18408
rect 4663 18377 4675 18380
rect 4617 18371 4675 18377
rect 4706 18368 4712 18380
rect 4764 18368 4770 18420
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 5997 18411 6055 18417
rect 5997 18408 6009 18411
rect 5960 18380 6009 18408
rect 5960 18368 5966 18380
rect 5997 18377 6009 18380
rect 6043 18408 6055 18411
rect 6549 18411 6607 18417
rect 6549 18408 6561 18411
rect 6043 18380 6561 18408
rect 6043 18377 6055 18380
rect 5997 18371 6055 18377
rect 6549 18377 6561 18380
rect 6595 18377 6607 18411
rect 8018 18408 8024 18420
rect 7979 18380 8024 18408
rect 6549 18371 6607 18377
rect 2593 18343 2651 18349
rect 2593 18309 2605 18343
rect 2639 18340 2651 18343
rect 2774 18340 2780 18352
rect 2639 18312 2780 18340
rect 2639 18309 2651 18312
rect 2593 18303 2651 18309
rect 2774 18300 2780 18312
rect 2832 18300 2838 18352
rect 2958 18340 2964 18352
rect 2919 18312 2964 18340
rect 2958 18300 2964 18312
rect 3016 18340 3022 18352
rect 5442 18340 5448 18352
rect 3016 18312 5448 18340
rect 3016 18300 3022 18312
rect 5442 18300 5448 18312
rect 5500 18300 5506 18352
rect 4157 18275 4215 18281
rect 4157 18241 4169 18275
rect 4203 18272 4215 18275
rect 4246 18272 4252 18284
rect 4203 18244 4252 18272
rect 4203 18241 4215 18244
rect 4157 18235 4215 18241
rect 4246 18232 4252 18244
rect 4304 18232 4310 18284
rect 6564 18272 6592 18371
rect 8018 18368 8024 18380
rect 8076 18368 8082 18420
rect 8478 18408 8484 18420
rect 8439 18380 8484 18408
rect 8478 18368 8484 18380
rect 8536 18368 8542 18420
rect 9582 18408 9588 18420
rect 9543 18380 9588 18408
rect 9582 18368 9588 18380
rect 9640 18368 9646 18420
rect 10134 18368 10140 18420
rect 10192 18408 10198 18420
rect 10321 18411 10379 18417
rect 10321 18408 10333 18411
rect 10192 18380 10333 18408
rect 10192 18368 10198 18380
rect 10321 18377 10333 18380
rect 10367 18377 10379 18411
rect 11422 18408 11428 18420
rect 11383 18380 11428 18408
rect 10321 18371 10379 18377
rect 11422 18368 11428 18380
rect 11480 18368 11486 18420
rect 6638 18300 6644 18352
rect 6696 18340 6702 18352
rect 7745 18343 7803 18349
rect 7745 18340 7757 18343
rect 6696 18312 7757 18340
rect 6696 18300 6702 18312
rect 7745 18309 7757 18312
rect 7791 18309 7803 18343
rect 7745 18303 7803 18309
rect 8849 18343 8907 18349
rect 8849 18309 8861 18343
rect 8895 18340 8907 18343
rect 9766 18340 9772 18352
rect 8895 18312 9772 18340
rect 8895 18309 8907 18312
rect 8849 18303 8907 18309
rect 9766 18300 9772 18312
rect 9824 18300 9830 18352
rect 6564 18244 6960 18272
rect 2409 18207 2467 18213
rect 2409 18173 2421 18207
rect 2455 18204 2467 18207
rect 2498 18204 2504 18216
rect 2455 18176 2504 18204
rect 2455 18173 2467 18176
rect 2409 18167 2467 18173
rect 2498 18164 2504 18176
rect 2556 18164 2562 18216
rect 2682 18164 2688 18216
rect 2740 18204 2746 18216
rect 3326 18204 3332 18216
rect 2740 18176 3332 18204
rect 2740 18164 2746 18176
rect 3326 18164 3332 18176
rect 3384 18204 3390 18216
rect 3421 18207 3479 18213
rect 3421 18204 3433 18207
rect 3384 18176 3433 18204
rect 3384 18164 3390 18176
rect 3421 18173 3433 18176
rect 3467 18173 3479 18207
rect 3421 18167 3479 18173
rect 3510 18164 3516 18216
rect 3568 18204 3574 18216
rect 3881 18207 3939 18213
rect 3881 18204 3893 18207
rect 3568 18176 3893 18204
rect 3568 18164 3574 18176
rect 3881 18173 3893 18176
rect 3927 18173 3939 18207
rect 3881 18167 3939 18173
rect 4338 18164 4344 18216
rect 4396 18204 4402 18216
rect 4982 18204 4988 18216
rect 4396 18176 4988 18204
rect 4396 18164 4402 18176
rect 4982 18164 4988 18176
rect 5040 18164 5046 18216
rect 5534 18204 5540 18216
rect 5495 18176 5540 18204
rect 5534 18164 5540 18176
rect 5592 18164 5598 18216
rect 5810 18164 5816 18216
rect 5868 18204 5874 18216
rect 6822 18204 6828 18216
rect 5868 18176 6828 18204
rect 5868 18164 5874 18176
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 5718 18136 5724 18148
rect 5679 18108 5724 18136
rect 5718 18096 5724 18108
rect 5776 18096 5782 18148
rect 6932 18136 6960 18244
rect 7098 18232 7104 18284
rect 7156 18272 7162 18284
rect 8018 18272 8024 18284
rect 7156 18244 8024 18272
rect 7156 18232 7162 18244
rect 8018 18232 8024 18244
rect 8076 18232 8082 18284
rect 9456 18275 9514 18281
rect 9456 18241 9468 18275
rect 9502 18272 9514 18275
rect 9582 18272 9588 18284
rect 9502 18244 9588 18272
rect 9502 18241 9514 18244
rect 9456 18235 9514 18241
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18272 9735 18275
rect 9858 18272 9864 18284
rect 9723 18244 9864 18272
rect 9723 18241 9735 18244
rect 9677 18235 9735 18241
rect 9858 18232 9864 18244
rect 9916 18272 9922 18284
rect 10152 18272 10180 18368
rect 11514 18272 11520 18284
rect 9916 18244 11520 18272
rect 9916 18232 9922 18244
rect 11514 18232 11520 18244
rect 11572 18232 11578 18284
rect 8570 18164 8576 18216
rect 8628 18204 8634 18216
rect 10045 18207 10103 18213
rect 10045 18204 10057 18207
rect 8628 18176 10057 18204
rect 8628 18164 8634 18176
rect 10045 18173 10057 18176
rect 10091 18173 10103 18207
rect 10045 18167 10103 18173
rect 10410 18164 10416 18216
rect 10468 18204 10474 18216
rect 10873 18207 10931 18213
rect 10873 18204 10885 18207
rect 10468 18176 10885 18204
rect 10468 18164 10474 18176
rect 10873 18173 10885 18176
rect 10919 18204 10931 18207
rect 11701 18207 11759 18213
rect 11701 18204 11713 18207
rect 10919 18176 11713 18204
rect 10919 18173 10931 18176
rect 10873 18167 10931 18173
rect 11701 18173 11713 18176
rect 11747 18173 11759 18207
rect 12434 18204 12440 18216
rect 12395 18176 12440 18204
rect 11701 18167 11759 18173
rect 12434 18164 12440 18176
rect 12492 18204 12498 18216
rect 12897 18207 12955 18213
rect 12897 18204 12909 18207
rect 12492 18176 12909 18204
rect 12492 18164 12498 18176
rect 12897 18173 12909 18176
rect 12943 18173 12955 18207
rect 12897 18167 12955 18173
rect 7146 18139 7204 18145
rect 7146 18136 7158 18139
rect 6932 18108 7158 18136
rect 7146 18105 7158 18108
rect 7192 18105 7204 18139
rect 9306 18136 9312 18148
rect 9219 18108 9312 18136
rect 7146 18099 7204 18105
rect 9306 18096 9312 18108
rect 9364 18136 9370 18148
rect 9364 18108 11836 18136
rect 9364 18096 9370 18108
rect 1394 18028 1400 18080
rect 1452 18068 1458 18080
rect 3326 18068 3332 18080
rect 1452 18040 3332 18068
rect 1452 18028 1458 18040
rect 3326 18028 3332 18040
rect 3384 18068 3390 18080
rect 4706 18068 4712 18080
rect 3384 18040 4712 18068
rect 3384 18028 3390 18040
rect 4706 18028 4712 18040
rect 4764 18028 4770 18080
rect 9217 18071 9275 18077
rect 9217 18037 9229 18071
rect 9263 18068 9275 18071
rect 9858 18068 9864 18080
rect 9263 18040 9864 18068
rect 9263 18037 9275 18040
rect 9217 18031 9275 18037
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 10778 18068 10784 18080
rect 10739 18040 10784 18068
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 10962 18028 10968 18080
rect 11020 18068 11026 18080
rect 11057 18071 11115 18077
rect 11057 18068 11069 18071
rect 11020 18040 11069 18068
rect 11020 18028 11026 18040
rect 11057 18037 11069 18040
rect 11103 18037 11115 18071
rect 11808 18068 11836 18108
rect 12621 18071 12679 18077
rect 12621 18068 12633 18071
rect 11808 18040 12633 18068
rect 11057 18031 11115 18037
rect 12621 18037 12633 18040
rect 12667 18037 12679 18071
rect 12621 18031 12679 18037
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 3145 17867 3203 17873
rect 3145 17833 3157 17867
rect 3191 17864 3203 17867
rect 3510 17864 3516 17876
rect 3191 17836 3516 17864
rect 3191 17833 3203 17836
rect 3145 17827 3203 17833
rect 3510 17824 3516 17836
rect 3568 17824 3574 17876
rect 4203 17867 4261 17873
rect 4203 17833 4215 17867
rect 4249 17864 4261 17867
rect 5626 17864 5632 17876
rect 4249 17836 5632 17864
rect 4249 17833 4261 17836
rect 4203 17827 4261 17833
rect 5626 17824 5632 17836
rect 5684 17824 5690 17876
rect 5718 17824 5724 17876
rect 5776 17864 5782 17876
rect 6089 17867 6147 17873
rect 6089 17864 6101 17867
rect 5776 17836 6101 17864
rect 5776 17824 5782 17836
rect 6089 17833 6101 17836
rect 6135 17833 6147 17867
rect 6089 17827 6147 17833
rect 6549 17867 6607 17873
rect 6549 17833 6561 17867
rect 6595 17864 6607 17867
rect 6638 17864 6644 17876
rect 6595 17836 6644 17864
rect 6595 17833 6607 17836
rect 6549 17827 6607 17833
rect 6638 17824 6644 17836
rect 6696 17864 6702 17876
rect 9306 17864 9312 17876
rect 6696 17836 6868 17864
rect 6696 17824 6702 17836
rect 2590 17756 2596 17808
rect 2648 17796 2654 17808
rect 5810 17796 5816 17808
rect 2648 17768 5028 17796
rect 5771 17768 5816 17796
rect 2648 17756 2654 17768
rect 2958 17728 2964 17740
rect 2919 17700 2964 17728
rect 2958 17688 2964 17700
rect 3016 17688 3022 17740
rect 4154 17737 4160 17740
rect 4132 17731 4160 17737
rect 4132 17697 4144 17731
rect 4132 17691 4160 17697
rect 4154 17688 4160 17691
rect 4212 17688 4218 17740
rect 5000 17669 5028 17768
rect 5810 17756 5816 17768
rect 5868 17756 5874 17808
rect 6730 17796 6736 17808
rect 6691 17768 6736 17796
rect 6730 17756 6736 17768
rect 6788 17756 6794 17808
rect 6840 17805 6868 17836
rect 8220 17836 9312 17864
rect 6825 17799 6883 17805
rect 6825 17765 6837 17799
rect 6871 17765 6883 17799
rect 6825 17759 6883 17765
rect 7377 17799 7435 17805
rect 7377 17765 7389 17799
rect 7423 17796 7435 17799
rect 7466 17796 7472 17808
rect 7423 17768 7472 17796
rect 7423 17765 7435 17768
rect 7377 17759 7435 17765
rect 7466 17756 7472 17768
rect 7524 17756 7530 17808
rect 8220 17805 8248 17836
rect 9306 17824 9312 17836
rect 9364 17824 9370 17876
rect 9674 17864 9680 17876
rect 9646 17824 9680 17864
rect 9732 17864 9738 17876
rect 9732 17836 10548 17864
rect 9732 17824 9738 17836
rect 8113 17799 8171 17805
rect 8113 17765 8125 17799
rect 8159 17796 8171 17799
rect 8205 17799 8263 17805
rect 8205 17796 8217 17799
rect 8159 17768 8217 17796
rect 8159 17765 8171 17768
rect 8113 17759 8171 17765
rect 8205 17765 8217 17768
rect 8251 17765 8263 17799
rect 8205 17759 8263 17765
rect 5258 17728 5264 17740
rect 5219 17700 5264 17728
rect 5258 17688 5264 17700
rect 5316 17688 5322 17740
rect 5534 17728 5540 17740
rect 5495 17700 5540 17728
rect 5534 17688 5540 17700
rect 5592 17688 5598 17740
rect 9646 17737 9674 17824
rect 10520 17796 10548 17836
rect 10594 17824 10600 17876
rect 10652 17864 10658 17876
rect 13265 17867 13323 17873
rect 13265 17864 13277 17867
rect 10652 17836 13277 17864
rect 10652 17824 10658 17836
rect 13265 17833 13277 17836
rect 13311 17833 13323 17867
rect 13265 17827 13323 17833
rect 10778 17796 10784 17808
rect 10520 17768 10784 17796
rect 10778 17756 10784 17768
rect 10836 17796 10842 17808
rect 10836 17768 12848 17796
rect 10836 17756 10842 17768
rect 12820 17740 12848 17768
rect 8389 17731 8447 17737
rect 8389 17697 8401 17731
rect 8435 17697 8447 17731
rect 9646 17731 9723 17737
rect 9646 17700 9677 17731
rect 8389 17691 8447 17697
rect 9665 17697 9677 17700
rect 9711 17697 9723 17731
rect 9665 17691 9723 17697
rect 4985 17663 5043 17669
rect 4985 17629 4997 17663
rect 5031 17660 5043 17663
rect 7374 17660 7380 17672
rect 5031 17632 7380 17660
rect 5031 17629 5043 17632
rect 4985 17623 5043 17629
rect 7374 17620 7380 17632
rect 7432 17620 7438 17672
rect 8294 17620 8300 17672
rect 8352 17660 8358 17672
rect 8404 17660 8432 17691
rect 9766 17688 9772 17740
rect 9824 17728 9830 17740
rect 9953 17731 10011 17737
rect 9824 17700 9869 17728
rect 9824 17688 9830 17700
rect 9953 17697 9965 17731
rect 9999 17728 10011 17731
rect 11514 17728 11520 17740
rect 9999 17700 11284 17728
rect 11475 17700 11520 17728
rect 9999 17697 10011 17700
rect 9953 17691 10011 17697
rect 11256 17672 11284 17700
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 12802 17728 12808 17740
rect 12763 17700 12808 17728
rect 12802 17688 12808 17700
rect 12860 17688 12866 17740
rect 13078 17728 13084 17740
rect 13039 17700 13084 17728
rect 13078 17688 13084 17700
rect 13136 17688 13142 17740
rect 10137 17663 10195 17669
rect 10137 17660 10149 17663
rect 8352 17632 10149 17660
rect 8352 17620 8358 17632
rect 10137 17629 10149 17632
rect 10183 17629 10195 17663
rect 11238 17660 11244 17672
rect 11199 17632 11244 17660
rect 10137 17623 10195 17629
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 2498 17592 2504 17604
rect 2411 17564 2504 17592
rect 2498 17552 2504 17564
rect 2556 17592 2562 17604
rect 6822 17592 6828 17604
rect 2556 17564 6828 17592
rect 2556 17552 2562 17564
rect 6822 17552 6828 17564
rect 6880 17552 6886 17604
rect 7745 17595 7803 17601
rect 7745 17561 7757 17595
rect 7791 17592 7803 17595
rect 8846 17592 8852 17604
rect 7791 17564 8852 17592
rect 7791 17561 7803 17564
rect 7745 17555 7803 17561
rect 8846 17552 8852 17564
rect 8904 17552 8910 17604
rect 12894 17592 12900 17604
rect 12855 17564 12900 17592
rect 12894 17552 12900 17564
rect 12952 17552 12958 17604
rect 4617 17527 4675 17533
rect 4617 17493 4629 17527
rect 4663 17524 4675 17527
rect 4706 17524 4712 17536
rect 4663 17496 4712 17524
rect 4663 17493 4675 17496
rect 4617 17487 4675 17493
rect 4706 17484 4712 17496
rect 4764 17484 4770 17536
rect 8478 17524 8484 17536
rect 8439 17496 8484 17524
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 5258 17320 5264 17332
rect 4126 17292 5264 17320
rect 3142 17212 3148 17264
rect 3200 17252 3206 17264
rect 3878 17252 3884 17264
rect 3200 17224 3884 17252
rect 3200 17212 3206 17224
rect 3878 17212 3884 17224
rect 3936 17252 3942 17264
rect 4126 17252 4154 17292
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 5629 17323 5687 17329
rect 5629 17320 5641 17323
rect 5592 17292 5641 17320
rect 5592 17280 5598 17292
rect 5629 17289 5641 17292
rect 5675 17289 5687 17323
rect 8294 17320 8300 17332
rect 8255 17292 8300 17320
rect 5629 17283 5687 17289
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 10045 17323 10103 17329
rect 10045 17320 10057 17323
rect 9824 17292 10057 17320
rect 9824 17280 9830 17292
rect 10045 17289 10057 17292
rect 10091 17320 10103 17323
rect 10413 17323 10471 17329
rect 10413 17320 10425 17323
rect 10091 17292 10425 17320
rect 10091 17289 10103 17292
rect 10045 17283 10103 17289
rect 10413 17289 10425 17292
rect 10459 17320 10471 17323
rect 10459 17292 10732 17320
rect 10459 17289 10471 17292
rect 10413 17283 10471 17289
rect 10704 17261 10732 17292
rect 11514 17280 11520 17332
rect 11572 17320 11578 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 11572 17292 11621 17320
rect 11572 17280 11578 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 11609 17283 11667 17289
rect 12802 17280 12808 17332
rect 12860 17320 12866 17332
rect 13541 17323 13599 17329
rect 13541 17320 13553 17323
rect 12860 17292 13553 17320
rect 12860 17280 12866 17292
rect 13541 17289 13553 17292
rect 13587 17289 13599 17323
rect 13541 17283 13599 17289
rect 3936 17224 4154 17252
rect 6273 17255 6331 17261
rect 3936 17212 3942 17224
rect 6273 17221 6285 17255
rect 6319 17252 6331 17255
rect 10689 17255 10747 17261
rect 6319 17224 7696 17252
rect 6319 17221 6331 17224
rect 6273 17215 6331 17221
rect 2958 17144 2964 17196
rect 3016 17184 3022 17196
rect 3053 17187 3111 17193
rect 3053 17184 3065 17187
rect 3016 17156 3065 17184
rect 3016 17144 3022 17156
rect 3053 17153 3065 17156
rect 3099 17184 3111 17187
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 3099 17156 7573 17184
rect 3099 17153 3111 17156
rect 3053 17147 3111 17153
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 3789 17119 3847 17125
rect 3789 17085 3801 17119
rect 3835 17116 3847 17119
rect 4062 17116 4068 17128
rect 3835 17088 4068 17116
rect 3835 17085 3847 17088
rect 3789 17079 3847 17085
rect 4062 17076 4068 17088
rect 4120 17116 4126 17128
rect 4249 17119 4307 17125
rect 4249 17116 4261 17119
rect 4120 17088 4261 17116
rect 4120 17076 4126 17088
rect 4249 17085 4261 17088
rect 4295 17085 4307 17119
rect 4706 17116 4712 17128
rect 4667 17088 4712 17116
rect 4249 17079 4307 17085
rect 4264 17048 4292 17079
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 6178 17116 6184 17128
rect 4816 17088 6184 17116
rect 4816 17048 4844 17088
rect 6178 17076 6184 17088
rect 6236 17076 6242 17128
rect 7101 17119 7159 17125
rect 7101 17085 7113 17119
rect 7147 17085 7159 17119
rect 7101 17079 7159 17085
rect 4982 17048 4988 17060
rect 4264 17020 4844 17048
rect 4943 17020 4988 17048
rect 4982 17008 4988 17020
rect 5040 17008 5046 17060
rect 6641 17051 6699 17057
rect 6641 17017 6653 17051
rect 6687 17048 6699 17051
rect 7116 17048 7144 17079
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 7377 17119 7435 17125
rect 7248 17088 7293 17116
rect 7248 17076 7254 17088
rect 7377 17085 7389 17119
rect 7423 17116 7435 17119
rect 7668 17116 7696 17224
rect 10689 17221 10701 17255
rect 10735 17221 10747 17255
rect 10689 17215 10747 17221
rect 13078 17212 13084 17264
rect 13136 17252 13142 17264
rect 13173 17255 13231 17261
rect 13173 17252 13185 17255
rect 13136 17224 13185 17252
rect 13136 17212 13142 17224
rect 13173 17221 13185 17224
rect 13219 17221 13231 17255
rect 13173 17215 13231 17221
rect 8570 17144 8576 17196
rect 8628 17184 8634 17196
rect 8628 17156 9536 17184
rect 8628 17144 8634 17156
rect 8202 17116 8208 17128
rect 7423 17088 8208 17116
rect 7423 17085 7435 17088
rect 7377 17079 7435 17085
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 8938 17116 8944 17128
rect 8899 17088 8944 17116
rect 8938 17076 8944 17088
rect 8996 17076 9002 17128
rect 9306 17116 9312 17128
rect 9267 17088 9312 17116
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 9508 17125 9536 17156
rect 11514 17144 11520 17196
rect 11572 17184 11578 17196
rect 11974 17184 11980 17196
rect 11572 17156 11980 17184
rect 11572 17144 11578 17156
rect 11974 17144 11980 17156
rect 12032 17144 12038 17196
rect 9493 17119 9551 17125
rect 9493 17085 9505 17119
rect 9539 17085 9551 17119
rect 10594 17116 10600 17128
rect 10555 17088 10600 17116
rect 9493 17079 9551 17085
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 10778 17076 10784 17128
rect 10836 17116 10842 17128
rect 10873 17119 10931 17125
rect 10873 17116 10885 17119
rect 10836 17088 10885 17116
rect 10836 17076 10842 17088
rect 10873 17085 10885 17088
rect 10919 17116 10931 17119
rect 11238 17116 11244 17128
rect 10919 17088 11244 17116
rect 10919 17085 10931 17088
rect 10873 17079 10931 17085
rect 11238 17076 11244 17088
rect 11296 17076 11302 17128
rect 7558 17048 7564 17060
rect 6687 17020 7564 17048
rect 6687 17017 6699 17020
rect 6641 17011 6699 17017
rect 7558 17008 7564 17020
rect 7616 17048 7622 17060
rect 8294 17048 8300 17060
rect 7616 17020 8300 17048
rect 7616 17008 7622 17020
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 11514 17048 11520 17060
rect 9324 17020 11520 17048
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 9324 16980 9352 17020
rect 11514 17008 11520 17020
rect 11572 17008 11578 17060
rect 12894 17048 12900 17060
rect 12807 17020 12900 17048
rect 12894 17008 12900 17020
rect 12952 17048 12958 17060
rect 14734 17048 14740 17060
rect 12952 17020 14740 17048
rect 12952 17008 12958 17020
rect 14734 17008 14740 17020
rect 14792 17008 14798 17060
rect 9766 16980 9772 16992
rect 4212 16952 9352 16980
rect 9727 16952 9772 16980
rect 4212 16940 4218 16952
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 11054 16980 11060 16992
rect 11015 16952 11060 16980
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 3878 16736 3884 16788
rect 3936 16776 3942 16788
rect 4062 16776 4068 16788
rect 3936 16748 4068 16776
rect 3936 16736 3942 16748
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 4982 16736 4988 16788
rect 5040 16776 5046 16788
rect 5261 16779 5319 16785
rect 5261 16776 5273 16779
rect 5040 16748 5273 16776
rect 5040 16736 5046 16748
rect 5261 16745 5273 16748
rect 5307 16745 5319 16779
rect 5261 16739 5319 16745
rect 5905 16779 5963 16785
rect 5905 16745 5917 16779
rect 5951 16776 5963 16779
rect 6730 16776 6736 16788
rect 5951 16748 6736 16776
rect 5951 16745 5963 16748
rect 5905 16739 5963 16745
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 8021 16779 8079 16785
rect 8021 16776 8033 16779
rect 6880 16748 8033 16776
rect 6880 16736 6886 16748
rect 8021 16745 8033 16748
rect 8067 16745 8079 16779
rect 8021 16739 8079 16745
rect 8757 16779 8815 16785
rect 8757 16745 8769 16779
rect 8803 16776 8815 16779
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 8803 16748 9137 16776
rect 8803 16745 8815 16748
rect 8757 16739 8815 16745
rect 9125 16745 9137 16748
rect 9171 16776 9183 16779
rect 9306 16776 9312 16788
rect 9171 16748 9312 16776
rect 9171 16745 9183 16748
rect 9125 16739 9183 16745
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 9493 16779 9551 16785
rect 9493 16745 9505 16779
rect 9539 16776 9551 16779
rect 10778 16776 10784 16788
rect 9539 16748 10784 16776
rect 9539 16745 9551 16748
rect 9493 16739 9551 16745
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 11330 16736 11336 16788
rect 11388 16776 11394 16788
rect 13679 16779 13737 16785
rect 13679 16776 13691 16779
rect 11388 16748 13691 16776
rect 11388 16736 11394 16748
rect 13679 16745 13691 16748
rect 13725 16745 13737 16779
rect 13679 16739 13737 16745
rect 8938 16668 8944 16720
rect 8996 16708 9002 16720
rect 10318 16708 10324 16720
rect 8996 16680 10324 16708
rect 8996 16668 9002 16680
rect 3418 16600 3424 16652
rect 3476 16640 3482 16652
rect 4246 16640 4252 16652
rect 3476 16612 4252 16640
rect 3476 16600 3482 16612
rect 4246 16600 4252 16612
rect 4304 16600 4310 16652
rect 4706 16640 4712 16652
rect 4619 16612 4712 16640
rect 4154 16532 4160 16584
rect 4212 16572 4218 16584
rect 4626 16572 4654 16612
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 6638 16640 6644 16652
rect 6551 16612 6644 16640
rect 6638 16600 6644 16612
rect 6696 16640 6702 16652
rect 7190 16640 7196 16652
rect 6696 16612 7196 16640
rect 6696 16600 6702 16612
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 7558 16640 7564 16652
rect 7519 16612 7564 16640
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 7650 16600 7656 16652
rect 7708 16640 7714 16652
rect 7837 16643 7895 16649
rect 7708 16612 7753 16640
rect 7708 16600 7714 16612
rect 7837 16609 7849 16643
rect 7883 16640 7895 16643
rect 8202 16640 8208 16652
rect 7883 16612 8208 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 9692 16649 9720 16680
rect 10318 16668 10324 16680
rect 10376 16708 10382 16720
rect 10962 16708 10968 16720
rect 10376 16680 10968 16708
rect 10376 16668 10382 16680
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 11977 16711 12035 16717
rect 11977 16677 11989 16711
rect 12023 16708 12035 16711
rect 12802 16708 12808 16720
rect 12023 16680 12808 16708
rect 12023 16677 12035 16680
rect 11977 16671 12035 16677
rect 12802 16668 12808 16680
rect 12860 16668 12866 16720
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 9950 16640 9956 16652
rect 9863 16612 9956 16640
rect 9677 16603 9735 16609
rect 9950 16600 9956 16612
rect 10008 16640 10014 16652
rect 10686 16640 10692 16652
rect 10008 16612 10692 16640
rect 10008 16600 10014 16612
rect 10686 16600 10692 16612
rect 10744 16600 10750 16652
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16640 11943 16643
rect 12342 16640 12348 16652
rect 11931 16612 12348 16640
rect 11931 16609 11943 16612
rect 11885 16603 11943 16609
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 13538 16640 13544 16652
rect 13499 16612 13544 16640
rect 13538 16600 13544 16612
rect 13596 16600 13602 16652
rect 4798 16572 4804 16584
rect 4212 16544 4654 16572
rect 4759 16544 4804 16572
rect 4212 16532 4218 16544
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 6733 16575 6791 16581
rect 6733 16541 6745 16575
rect 6779 16572 6791 16575
rect 7668 16572 7696 16600
rect 10134 16572 10140 16584
rect 6779 16544 7696 16572
rect 10095 16544 10140 16572
rect 6779 16541 6791 16544
rect 6733 16535 6791 16541
rect 10134 16532 10140 16544
rect 10192 16532 10198 16584
rect 10594 16532 10600 16584
rect 10652 16572 10658 16584
rect 11057 16575 11115 16581
rect 11057 16572 11069 16575
rect 10652 16544 11069 16572
rect 10652 16532 10658 16544
rect 11057 16541 11069 16544
rect 11103 16541 11115 16575
rect 11057 16535 11115 16541
rect 11238 16532 11244 16584
rect 11296 16572 11302 16584
rect 12710 16572 12716 16584
rect 11296 16544 12716 16572
rect 11296 16532 11302 16544
rect 12710 16532 12716 16544
rect 12768 16532 12774 16584
rect 7190 16504 7196 16516
rect 7103 16476 7196 16504
rect 7190 16464 7196 16476
rect 7248 16504 7254 16516
rect 9769 16507 9827 16513
rect 9769 16504 9781 16507
rect 7248 16476 9781 16504
rect 7248 16464 7254 16476
rect 9769 16473 9781 16476
rect 9815 16504 9827 16507
rect 10042 16504 10048 16516
rect 9815 16476 10048 16504
rect 9815 16473 9827 16476
rect 9769 16467 9827 16473
rect 10042 16464 10048 16476
rect 10100 16504 10106 16516
rect 12894 16504 12900 16516
rect 10100 16476 12900 16504
rect 10100 16464 10106 16476
rect 12894 16464 12900 16476
rect 12952 16464 12958 16516
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 3510 16192 3516 16244
rect 3568 16232 3574 16244
rect 3743 16235 3801 16241
rect 3743 16232 3755 16235
rect 3568 16204 3755 16232
rect 3568 16192 3574 16204
rect 3743 16201 3755 16204
rect 3789 16201 3801 16235
rect 4522 16232 4528 16244
rect 4483 16204 4528 16232
rect 3743 16195 3801 16201
rect 4522 16192 4528 16204
rect 4580 16192 4586 16244
rect 6089 16235 6147 16241
rect 6089 16201 6101 16235
rect 6135 16232 6147 16235
rect 6638 16232 6644 16244
rect 6135 16204 6644 16232
rect 6135 16201 6147 16204
rect 6089 16195 6147 16201
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 7650 16192 7656 16244
rect 7708 16232 7714 16244
rect 7837 16235 7895 16241
rect 7837 16232 7849 16235
rect 7708 16204 7849 16232
rect 7708 16192 7714 16204
rect 7837 16201 7849 16204
rect 7883 16201 7895 16235
rect 10042 16232 10048 16244
rect 10003 16204 10048 16232
rect 7837 16195 7895 16201
rect 10042 16192 10048 16204
rect 10100 16192 10106 16244
rect 4246 16124 4252 16176
rect 4304 16164 4310 16176
rect 6549 16167 6607 16173
rect 6549 16164 6561 16167
rect 4304 16136 6561 16164
rect 4304 16124 4310 16136
rect 6549 16133 6561 16136
rect 6595 16133 6607 16167
rect 12158 16164 12164 16176
rect 6549 16127 6607 16133
rect 9876 16136 12164 16164
rect 4617 16099 4675 16105
rect 4617 16065 4629 16099
rect 4663 16096 4675 16099
rect 4982 16096 4988 16108
rect 4663 16068 4988 16096
rect 4663 16065 4675 16068
rect 4617 16059 4675 16065
rect 4982 16056 4988 16068
rect 5040 16056 5046 16108
rect 3513 16031 3571 16037
rect 3513 15997 3525 16031
rect 3559 16028 3571 16031
rect 3640 16031 3698 16037
rect 3640 16028 3652 16031
rect 3559 16000 3652 16028
rect 3559 15997 3571 16000
rect 3513 15991 3571 15997
rect 3640 15997 3652 16000
rect 3686 16028 3698 16031
rect 5074 16028 5080 16040
rect 3686 16000 5080 16028
rect 3686 15997 3698 16000
rect 3640 15991 3698 15997
rect 5074 15988 5080 16000
rect 5132 15988 5138 16040
rect 6564 16028 6592 16127
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16096 8631 16099
rect 8754 16096 8760 16108
rect 8619 16068 8760 16096
rect 8619 16065 8631 16068
rect 8573 16059 8631 16065
rect 8754 16056 8760 16068
rect 8812 16096 8818 16108
rect 8812 16068 9536 16096
rect 8812 16056 8818 16068
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6564 16000 6837 16028
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 7374 16028 7380 16040
rect 7335 16000 7380 16028
rect 6825 15991 6883 15997
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 8846 16028 8852 16040
rect 8807 16000 8852 16028
rect 8846 15988 8852 16000
rect 8904 15988 8910 16040
rect 9306 16028 9312 16040
rect 9267 16000 9312 16028
rect 9306 15988 9312 16000
rect 9364 15988 9370 16040
rect 9508 16037 9536 16068
rect 9493 16031 9551 16037
rect 9493 15997 9505 16031
rect 9539 16028 9551 16031
rect 9876 16028 9904 16136
rect 12158 16124 12164 16136
rect 12216 16124 12222 16176
rect 10873 16099 10931 16105
rect 10873 16065 10885 16099
rect 10919 16096 10931 16099
rect 11146 16096 11152 16108
rect 10919 16068 11152 16096
rect 10919 16065 10931 16068
rect 10873 16059 10931 16065
rect 11146 16056 11152 16068
rect 11204 16096 11210 16108
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 11204 16068 12449 16096
rect 11204 16056 11210 16068
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 9539 16000 9904 16028
rect 9539 15997 9551 16000
rect 9493 15991 9551 15997
rect 4522 15920 4528 15972
rect 4580 15960 4586 15972
rect 4938 15963 4996 15969
rect 4938 15960 4950 15963
rect 4580 15932 4950 15960
rect 4580 15920 4586 15932
rect 4938 15929 4950 15932
rect 4984 15929 4996 15963
rect 4938 15923 4996 15929
rect 10962 15920 10968 15972
rect 11020 15960 11026 15972
rect 11517 15963 11575 15969
rect 11020 15932 11065 15960
rect 11020 15920 11026 15932
rect 11517 15929 11529 15963
rect 11563 15960 11575 15963
rect 11974 15960 11980 15972
rect 11563 15932 11980 15960
rect 11563 15929 11575 15932
rect 11517 15923 11575 15929
rect 11974 15920 11980 15932
rect 12032 15960 12038 15972
rect 13538 15960 13544 15972
rect 12032 15932 13544 15960
rect 12032 15920 12038 15932
rect 13538 15920 13544 15932
rect 13596 15920 13602 15972
rect 4157 15895 4215 15901
rect 4157 15861 4169 15895
rect 4203 15892 4215 15895
rect 4246 15892 4252 15904
rect 4203 15864 4252 15892
rect 4203 15861 4215 15864
rect 4157 15855 4215 15861
rect 4246 15852 4252 15864
rect 4304 15852 4310 15904
rect 5534 15892 5540 15904
rect 5495 15864 5540 15892
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 7101 15895 7159 15901
rect 7101 15861 7113 15895
rect 7147 15892 7159 15895
rect 7282 15892 7288 15904
rect 7147 15864 7288 15892
rect 7147 15861 7159 15864
rect 7101 15855 7159 15861
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 9582 15892 9588 15904
rect 9543 15864 9588 15892
rect 9582 15852 9588 15864
rect 9640 15852 9646 15904
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 10980 15892 11008 15920
rect 10735 15864 11008 15892
rect 11885 15895 11943 15901
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 11885 15861 11897 15895
rect 11931 15892 11943 15895
rect 12342 15892 12348 15904
rect 11931 15864 12348 15892
rect 11931 15861 11943 15864
rect 11885 15855 11943 15861
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 5074 15648 5080 15700
rect 5132 15688 5138 15700
rect 5132 15660 7144 15688
rect 5132 15648 5138 15660
rect 4522 15580 4528 15632
rect 4580 15620 4586 15632
rect 4982 15629 4988 15632
rect 4938 15623 4988 15629
rect 4938 15620 4950 15623
rect 4580 15592 4950 15620
rect 4580 15580 4586 15592
rect 4938 15589 4950 15592
rect 4984 15589 4988 15623
rect 4938 15583 4988 15589
rect 4982 15580 4988 15583
rect 5040 15580 5046 15632
rect 5534 15580 5540 15632
rect 5592 15620 5598 15632
rect 6546 15620 6552 15632
rect 5592 15592 6552 15620
rect 5592 15580 5598 15592
rect 6546 15580 6552 15592
rect 6604 15580 6610 15632
rect 7116 15629 7144 15660
rect 7558 15648 7564 15700
rect 7616 15688 7622 15700
rect 7745 15691 7803 15697
rect 7745 15688 7757 15691
rect 7616 15660 7757 15688
rect 7616 15648 7622 15660
rect 7745 15657 7757 15660
rect 7791 15657 7803 15691
rect 7745 15651 7803 15657
rect 9033 15691 9091 15697
rect 9033 15657 9045 15691
rect 9079 15688 9091 15691
rect 9398 15688 9404 15700
rect 9079 15660 9404 15688
rect 9079 15657 9091 15660
rect 9033 15651 9091 15657
rect 7101 15623 7159 15629
rect 7101 15589 7113 15623
rect 7147 15620 7159 15623
rect 7190 15620 7196 15632
rect 7147 15592 7196 15620
rect 7147 15589 7159 15592
rect 7101 15583 7159 15589
rect 7190 15580 7196 15592
rect 7248 15580 7254 15632
rect 8846 15620 8852 15632
rect 7944 15592 8852 15620
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15552 4675 15555
rect 4798 15552 4804 15564
rect 4663 15524 4804 15552
rect 4663 15521 4675 15524
rect 4617 15515 4675 15521
rect 4798 15512 4804 15524
rect 4856 15512 4862 15564
rect 7944 15561 7972 15592
rect 8846 15580 8852 15592
rect 8904 15580 8910 15632
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15521 7987 15555
rect 8202 15552 8208 15564
rect 8115 15524 8208 15552
rect 7929 15515 7987 15521
rect 8202 15512 8208 15524
rect 8260 15552 8266 15564
rect 9048 15552 9076 15651
rect 9398 15648 9404 15660
rect 9456 15688 9462 15700
rect 9493 15691 9551 15697
rect 9493 15688 9505 15691
rect 9456 15660 9505 15688
rect 9456 15648 9462 15660
rect 9493 15657 9505 15660
rect 9539 15688 9551 15691
rect 9950 15688 9956 15700
rect 9539 15660 9956 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 11146 15688 11152 15700
rect 11107 15660 11152 15688
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 10182 15623 10240 15629
rect 10182 15620 10194 15623
rect 9968 15592 10194 15620
rect 9968 15564 9996 15592
rect 10182 15589 10194 15592
rect 10228 15589 10240 15623
rect 11790 15620 11796 15632
rect 10182 15583 10240 15589
rect 10796 15592 11796 15620
rect 8260 15524 9076 15552
rect 8260 15512 8266 15524
rect 9766 15512 9772 15564
rect 9824 15552 9830 15564
rect 9861 15555 9919 15561
rect 9861 15552 9873 15555
rect 9824 15524 9873 15552
rect 9824 15512 9830 15524
rect 9861 15521 9873 15524
rect 9907 15521 9919 15555
rect 9861 15515 9919 15521
rect 9950 15512 9956 15564
rect 10008 15512 10014 15564
rect 10796 15561 10824 15592
rect 11790 15580 11796 15592
rect 11848 15580 11854 15632
rect 10781 15555 10839 15561
rect 10781 15521 10793 15555
rect 10827 15521 10839 15555
rect 10781 15515 10839 15521
rect 2958 15484 2964 15496
rect 2919 15456 2964 15484
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15453 6515 15487
rect 6457 15447 6515 15453
rect 4154 15308 4160 15360
rect 4212 15348 4218 15360
rect 4249 15351 4307 15357
rect 4249 15348 4261 15351
rect 4212 15320 4261 15348
rect 4212 15308 4218 15320
rect 4249 15317 4261 15320
rect 4295 15317 4307 15351
rect 5534 15348 5540 15360
rect 5495 15320 5540 15348
rect 4249 15311 4307 15317
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 5626 15308 5632 15360
rect 5684 15348 5690 15360
rect 6181 15351 6239 15357
rect 6181 15348 6193 15351
rect 5684 15320 6193 15348
rect 5684 15308 5690 15320
rect 6181 15317 6193 15320
rect 6227 15348 6239 15351
rect 6472 15348 6500 15447
rect 7650 15444 7656 15496
rect 7708 15484 7714 15496
rect 8021 15487 8079 15493
rect 8021 15484 8033 15487
rect 7708 15456 8033 15484
rect 7708 15444 7714 15456
rect 8021 15453 8033 15456
rect 8067 15453 8079 15487
rect 8021 15447 8079 15453
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 8389 15487 8447 15493
rect 8389 15484 8401 15487
rect 8352 15456 8401 15484
rect 8352 15444 8358 15456
rect 8389 15453 8401 15456
rect 8435 15453 8447 15487
rect 11698 15484 11704 15496
rect 11659 15456 11704 15484
rect 8389 15447 8447 15453
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 11974 15484 11980 15496
rect 11935 15456 11980 15484
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 6227 15320 6500 15348
rect 6227 15317 6239 15320
rect 6181 15311 6239 15317
rect 7374 15308 7380 15360
rect 7432 15348 7438 15360
rect 7469 15351 7527 15357
rect 7469 15348 7481 15351
rect 7432 15320 7481 15348
rect 7432 15308 7438 15320
rect 7469 15317 7481 15320
rect 7515 15348 7527 15351
rect 8570 15348 8576 15360
rect 7515 15320 8576 15348
rect 7515 15317 7527 15320
rect 7469 15311 7527 15317
rect 8570 15308 8576 15320
rect 8628 15308 8634 15360
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 4798 15104 4804 15156
rect 4856 15144 4862 15156
rect 5537 15147 5595 15153
rect 5537 15144 5549 15147
rect 4856 15116 5549 15144
rect 4856 15104 4862 15116
rect 5537 15113 5549 15116
rect 5583 15113 5595 15147
rect 6546 15144 6552 15156
rect 6507 15116 6552 15144
rect 5537 15107 5595 15113
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 7650 15104 7656 15156
rect 7708 15144 7714 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7708 15116 7849 15144
rect 7708 15104 7714 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 9398 15144 9404 15156
rect 9359 15116 9404 15144
rect 7837 15107 7895 15113
rect 9398 15104 9404 15116
rect 9456 15104 9462 15156
rect 10318 15144 10324 15156
rect 10279 15116 10324 15144
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 10962 15104 10968 15156
rect 11020 15144 11026 15156
rect 11057 15147 11115 15153
rect 11057 15144 11069 15147
rect 11020 15116 11069 15144
rect 11020 15104 11026 15116
rect 11057 15113 11069 15116
rect 11103 15113 11115 15147
rect 11790 15144 11796 15156
rect 11751 15116 11796 15144
rect 11057 15107 11115 15113
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 3881 15079 3939 15085
rect 3881 15045 3893 15079
rect 3927 15076 3939 15079
rect 4430 15076 4436 15088
rect 3927 15048 4436 15076
rect 3927 15045 3939 15048
rect 3881 15039 3939 15045
rect 4430 15036 4436 15048
rect 4488 15076 4494 15088
rect 4982 15076 4988 15088
rect 4488 15048 4988 15076
rect 4488 15036 4494 15048
rect 4982 15036 4988 15048
rect 5040 15076 5046 15088
rect 5169 15079 5227 15085
rect 5169 15076 5181 15079
rect 5040 15048 5181 15076
rect 5040 15036 5046 15048
rect 5169 15045 5181 15048
rect 5215 15045 5227 15079
rect 5169 15039 5227 15045
rect 5905 15079 5963 15085
rect 5905 15045 5917 15079
rect 5951 15045 5963 15079
rect 5905 15039 5963 15045
rect 6273 15079 6331 15085
rect 6273 15045 6285 15079
rect 6319 15076 6331 15079
rect 8478 15076 8484 15088
rect 6319 15048 8484 15076
rect 6319 15045 6331 15048
rect 6273 15039 6331 15045
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 15008 2375 15011
rect 4154 15008 4160 15020
rect 2363 14980 4160 15008
rect 2363 14977 2375 14980
rect 2317 14971 2375 14977
rect 2682 14940 2688 14952
rect 2643 14912 2688 14940
rect 2682 14900 2688 14912
rect 2740 14900 2746 14952
rect 2976 14949 3004 14980
rect 4154 14968 4160 14980
rect 4212 15008 4218 15020
rect 5920 15008 5948 15039
rect 4212 14980 5948 15008
rect 4212 14968 4218 14980
rect 2961 14943 3019 14949
rect 2961 14909 2973 14943
rect 3007 14909 3019 14943
rect 2961 14903 3019 14909
rect 3973 14943 4031 14949
rect 3973 14909 3985 14943
rect 4019 14909 4031 14943
rect 3973 14903 4031 14909
rect 5721 14943 5779 14949
rect 5721 14909 5733 14943
rect 5767 14940 5779 14943
rect 6288 14940 6316 15039
rect 8478 15036 8484 15048
rect 8536 15036 8542 15088
rect 7190 15008 7196 15020
rect 7151 14980 7196 15008
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 5767 14912 6316 14940
rect 5767 14909 5779 14912
rect 5721 14903 5779 14909
rect 3145 14875 3203 14881
rect 3145 14841 3157 14875
rect 3191 14872 3203 14875
rect 3421 14875 3479 14881
rect 3421 14872 3433 14875
rect 3191 14844 3433 14872
rect 3191 14841 3203 14844
rect 3145 14835 3203 14841
rect 3421 14841 3433 14844
rect 3467 14872 3479 14875
rect 3988 14872 4016 14903
rect 8202 14900 8208 14952
rect 8260 14940 8266 14952
rect 8389 14943 8447 14949
rect 8389 14940 8401 14943
rect 8260 14912 8401 14940
rect 8260 14900 8266 14912
rect 8389 14909 8401 14912
rect 8435 14909 8447 14943
rect 8389 14903 8447 14909
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 8849 14943 8907 14949
rect 8849 14940 8861 14943
rect 8628 14912 8861 14940
rect 8628 14900 8634 14912
rect 8849 14909 8861 14912
rect 8895 14909 8907 14943
rect 8849 14903 8907 14909
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14940 10747 14943
rect 11425 14943 11483 14949
rect 11425 14940 11437 14943
rect 10735 14912 11437 14940
rect 10735 14909 10747 14912
rect 10689 14903 10747 14909
rect 11425 14909 11437 14912
rect 11471 14940 11483 14943
rect 11790 14940 11796 14952
rect 11471 14912 11796 14940
rect 11471 14909 11483 14912
rect 11425 14903 11483 14909
rect 11790 14900 11796 14912
rect 11848 14900 11854 14952
rect 3467 14844 4016 14872
rect 4335 14875 4393 14881
rect 3467 14841 3479 14844
rect 3421 14835 3479 14841
rect 4335 14841 4347 14875
rect 4381 14872 4393 14875
rect 4430 14872 4436 14884
rect 4381 14844 4436 14872
rect 4381 14841 4393 14844
rect 4335 14835 4393 14841
rect 4430 14832 4436 14844
rect 4488 14832 4494 14884
rect 5534 14832 5540 14884
rect 5592 14872 5598 14884
rect 6914 14872 6920 14884
rect 5592 14844 6770 14872
rect 6875 14844 6920 14872
rect 5592 14832 5598 14844
rect 6742 14816 6770 14844
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 7009 14875 7067 14881
rect 7009 14841 7021 14875
rect 7055 14841 7067 14875
rect 7009 14835 7067 14841
rect 4890 14804 4896 14816
rect 4851 14776 4896 14804
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 6730 14804 6736 14816
rect 6643 14776 6736 14804
rect 6730 14764 6736 14776
rect 6788 14804 6794 14816
rect 7024 14804 7052 14835
rect 11698 14832 11704 14884
rect 11756 14832 11762 14884
rect 8202 14804 8208 14816
rect 6788 14776 7052 14804
rect 8163 14776 8208 14804
rect 6788 14764 6794 14776
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 8478 14804 8484 14816
rect 8439 14776 8484 14804
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 9858 14804 9864 14816
rect 9819 14776 9864 14804
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 11716 14804 11744 14832
rect 12161 14807 12219 14813
rect 12161 14804 12173 14807
rect 10652 14776 12173 14804
rect 10652 14764 10658 14776
rect 12161 14773 12173 14776
rect 12207 14773 12219 14807
rect 12161 14767 12219 14773
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 2501 14603 2559 14609
rect 2501 14569 2513 14603
rect 2547 14600 2559 14603
rect 2682 14600 2688 14612
rect 2547 14572 2688 14600
rect 2547 14569 2559 14572
rect 2501 14563 2559 14569
rect 2682 14560 2688 14572
rect 2740 14560 2746 14612
rect 5902 14560 5908 14612
rect 5960 14600 5966 14612
rect 6181 14603 6239 14609
rect 6181 14600 6193 14603
rect 5960 14572 6193 14600
rect 5960 14560 5966 14572
rect 6181 14569 6193 14572
rect 6227 14600 6239 14603
rect 6914 14600 6920 14612
rect 6227 14572 6920 14600
rect 6227 14569 6239 14572
rect 6181 14563 6239 14569
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 7193 14603 7251 14609
rect 7193 14569 7205 14603
rect 7239 14600 7251 14603
rect 8846 14600 8852 14612
rect 7239 14572 8852 14600
rect 7239 14569 7251 14572
rect 7193 14563 7251 14569
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 9493 14603 9551 14609
rect 9493 14569 9505 14603
rect 9539 14600 9551 14603
rect 9766 14600 9772 14612
rect 9539 14572 9772 14600
rect 9539 14569 9551 14572
rect 9493 14563 9551 14569
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 4706 14532 4712 14544
rect 4619 14504 4712 14532
rect 4706 14492 4712 14504
rect 4764 14532 4770 14544
rect 4890 14532 4896 14544
rect 4764 14504 4896 14532
rect 4764 14492 4770 14504
rect 4890 14492 4896 14504
rect 4948 14492 4954 14544
rect 4982 14492 4988 14544
rect 5040 14532 5046 14544
rect 6730 14532 6736 14544
rect 5040 14504 6592 14532
rect 6691 14504 6736 14532
rect 5040 14492 5046 14504
rect 6273 14467 6331 14473
rect 6273 14433 6285 14467
rect 6319 14433 6331 14467
rect 6564 14464 6592 14504
rect 6730 14492 6736 14504
rect 6788 14492 6794 14544
rect 7098 14532 7104 14544
rect 6840 14504 7104 14532
rect 6840 14464 6868 14504
rect 7098 14492 7104 14504
rect 7156 14532 7162 14544
rect 7606 14535 7664 14541
rect 7606 14532 7618 14535
rect 7156 14504 7618 14532
rect 7156 14492 7162 14504
rect 7606 14501 7618 14504
rect 7652 14532 7664 14535
rect 9858 14532 9864 14544
rect 7652 14504 9864 14532
rect 7652 14501 7664 14504
rect 7606 14495 7664 14501
rect 9858 14492 9864 14504
rect 9916 14532 9922 14544
rect 9998 14535 10056 14541
rect 9998 14532 10010 14535
rect 9916 14504 10010 14532
rect 9916 14492 9922 14504
rect 9998 14501 10010 14504
rect 10044 14501 10056 14535
rect 9998 14495 10056 14501
rect 6564 14436 6868 14464
rect 7285 14467 7343 14473
rect 6273 14427 6331 14433
rect 7285 14433 7297 14467
rect 7331 14464 7343 14467
rect 7742 14464 7748 14476
rect 7331 14436 7748 14464
rect 7331 14433 7343 14436
rect 7285 14427 7343 14433
rect 2958 14356 2964 14408
rect 3016 14396 3022 14408
rect 4614 14396 4620 14408
rect 3016 14368 4620 14396
rect 3016 14356 3022 14368
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 5074 14396 5080 14408
rect 5035 14368 5080 14396
rect 5074 14356 5080 14368
rect 5132 14356 5138 14408
rect 6288 14396 6316 14427
rect 7742 14424 7748 14436
rect 7800 14464 7806 14476
rect 8478 14464 8484 14476
rect 7800 14436 8484 14464
rect 7800 14424 7806 14436
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 9582 14424 9588 14476
rect 9640 14464 9646 14476
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 9640 14436 9689 14464
rect 9640 14424 9646 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 11330 14424 11336 14476
rect 11388 14464 11394 14476
rect 11460 14467 11518 14473
rect 11460 14464 11472 14467
rect 11388 14436 11472 14464
rect 11388 14424 11394 14436
rect 11460 14433 11472 14436
rect 11506 14433 11518 14467
rect 11460 14427 11518 14433
rect 6362 14396 6368 14408
rect 6275 14368 6368 14396
rect 6362 14356 6368 14368
rect 6420 14396 6426 14408
rect 11054 14396 11060 14408
rect 6420 14368 11060 14396
rect 6420 14356 6426 14368
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 4430 14288 4436 14340
rect 4488 14328 4494 14340
rect 6457 14331 6515 14337
rect 6457 14328 6469 14331
rect 4488 14300 6469 14328
rect 4488 14288 4494 14300
rect 6457 14297 6469 14300
rect 6503 14328 6515 14331
rect 7374 14328 7380 14340
rect 6503 14300 7380 14328
rect 6503 14297 6515 14300
rect 6457 14291 6515 14297
rect 7374 14288 7380 14300
rect 7432 14288 7438 14340
rect 11330 14288 11336 14340
rect 11388 14328 11394 14340
rect 13262 14328 13268 14340
rect 11388 14300 13268 14328
rect 11388 14288 11394 14300
rect 13262 14288 13268 14300
rect 13320 14288 13326 14340
rect 4246 14220 4252 14272
rect 4304 14260 4310 14272
rect 4798 14260 4804 14272
rect 4304 14232 4804 14260
rect 4304 14220 4310 14232
rect 4798 14220 4804 14232
rect 4856 14220 4862 14272
rect 5258 14220 5264 14272
rect 5316 14260 5322 14272
rect 5537 14263 5595 14269
rect 5537 14260 5549 14263
rect 5316 14232 5549 14260
rect 5316 14220 5322 14232
rect 5537 14229 5549 14232
rect 5583 14229 5595 14263
rect 8202 14260 8208 14272
rect 8163 14232 8208 14260
rect 5537 14223 5595 14229
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 8570 14260 8576 14272
rect 8531 14232 8576 14260
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 10597 14263 10655 14269
rect 10597 14229 10609 14263
rect 10643 14260 10655 14263
rect 10686 14260 10692 14272
rect 10643 14232 10692 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 11563 14263 11621 14269
rect 11563 14260 11575 14263
rect 11020 14232 11575 14260
rect 11020 14220 11026 14232
rect 11563 14229 11575 14232
rect 11609 14229 11621 14263
rect 11563 14223 11621 14229
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 4614 14056 4620 14068
rect 4575 14028 4620 14056
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 6362 14056 6368 14068
rect 6323 14028 6368 14056
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 7098 14056 7104 14068
rect 7059 14028 7104 14056
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 9033 14059 9091 14065
rect 9033 14025 9045 14059
rect 9079 14056 9091 14059
rect 9490 14056 9496 14068
rect 9079 14028 9496 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 9858 14056 9864 14068
rect 9815 14028 9864 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 10962 14056 10968 14068
rect 10923 14028 10968 14056
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11514 14056 11520 14068
rect 11112 14028 11520 14056
rect 11112 14016 11118 14028
rect 11514 14016 11520 14028
rect 11572 14016 11578 14068
rect 10134 13988 10140 14000
rect 9508 13960 10140 13988
rect 9508 13932 9536 13960
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 3513 13923 3571 13929
rect 3513 13889 3525 13923
rect 3559 13920 3571 13923
rect 4430 13920 4436 13932
rect 3559 13892 4436 13920
rect 3559 13889 3571 13892
rect 3513 13883 3571 13889
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 3602 13852 3608 13864
rect 2740 13824 3608 13852
rect 2740 13812 2746 13824
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 4172 13861 4200 13892
rect 4430 13880 4436 13892
rect 4488 13880 4494 13932
rect 7282 13920 7288 13932
rect 7243 13892 7288 13920
rect 7282 13880 7288 13892
rect 7340 13920 7346 13932
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 7340 13892 8493 13920
rect 7340 13880 7346 13892
rect 8481 13889 8493 13892
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 9490 13880 9496 13932
rect 9548 13880 9554 13932
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13920 10011 13923
rect 10980 13920 11008 14016
rect 9999 13892 11008 13920
rect 9999 13889 10011 13892
rect 9953 13883 10011 13889
rect 4157 13855 4215 13861
rect 4157 13821 4169 13855
rect 4203 13821 4215 13855
rect 4157 13815 4215 13821
rect 4341 13855 4399 13861
rect 4341 13821 4353 13855
rect 4387 13852 4399 13855
rect 5074 13852 5080 13864
rect 4387 13824 5080 13852
rect 4387 13821 4399 13824
rect 4341 13815 4399 13821
rect 5074 13812 5080 13824
rect 5132 13812 5138 13864
rect 5258 13784 5264 13796
rect 5219 13756 5264 13784
rect 5258 13744 5264 13756
rect 5316 13744 5322 13796
rect 5350 13744 5356 13796
rect 5408 13784 5414 13796
rect 5905 13787 5963 13793
rect 5408 13756 5453 13784
rect 5408 13744 5414 13756
rect 5905 13753 5917 13787
rect 5951 13753 5963 13787
rect 5905 13747 5963 13753
rect 5077 13719 5135 13725
rect 5077 13685 5089 13719
rect 5123 13716 5135 13719
rect 5368 13716 5396 13744
rect 5123 13688 5396 13716
rect 5123 13685 5135 13688
rect 5077 13679 5135 13685
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 5920 13716 5948 13747
rect 7098 13744 7104 13796
rect 7156 13784 7162 13796
rect 7606 13787 7664 13793
rect 7606 13784 7618 13787
rect 7156 13756 7618 13784
rect 7156 13744 7162 13756
rect 7606 13753 7618 13756
rect 7652 13753 7664 13787
rect 7606 13747 7664 13753
rect 8110 13744 8116 13796
rect 8168 13784 8174 13796
rect 9306 13784 9312 13796
rect 8168 13756 9312 13784
rect 8168 13744 8174 13756
rect 9306 13744 9312 13756
rect 9364 13744 9370 13796
rect 9401 13787 9459 13793
rect 9401 13753 9413 13787
rect 9447 13784 9459 13787
rect 10045 13787 10103 13793
rect 10045 13784 10057 13787
rect 9447 13756 10057 13784
rect 9447 13753 9459 13756
rect 9401 13747 9459 13753
rect 10045 13753 10057 13756
rect 10091 13753 10103 13787
rect 10594 13784 10600 13796
rect 10555 13756 10600 13784
rect 10045 13747 10103 13753
rect 5868 13688 5948 13716
rect 8205 13719 8263 13725
rect 5868 13676 5874 13688
rect 8205 13685 8217 13719
rect 8251 13716 8263 13719
rect 8386 13716 8392 13728
rect 8251 13688 8392 13716
rect 8251 13685 8263 13688
rect 8205 13679 8263 13685
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 10060 13716 10088 13747
rect 10594 13744 10600 13756
rect 10652 13744 10658 13796
rect 10686 13716 10692 13728
rect 10060 13688 10692 13716
rect 10686 13676 10692 13688
rect 10744 13676 10750 13728
rect 11422 13716 11428 13728
rect 11383 13688 11428 13716
rect 11422 13676 11428 13688
rect 11480 13676 11486 13728
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 3602 13512 3608 13524
rect 3563 13484 3608 13512
rect 3602 13472 3608 13484
rect 3660 13472 3666 13524
rect 4614 13512 4620 13524
rect 4575 13484 4620 13512
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7285 13515 7343 13521
rect 7285 13512 7297 13515
rect 7156 13484 7297 13512
rect 7156 13472 7162 13484
rect 7285 13481 7297 13484
rect 7331 13481 7343 13515
rect 7742 13512 7748 13524
rect 7703 13484 7748 13512
rect 7285 13475 7343 13481
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 3099 13447 3157 13453
rect 3099 13413 3111 13447
rect 3145 13444 3157 13447
rect 5258 13444 5264 13456
rect 3145 13416 5264 13444
rect 3145 13413 3157 13416
rect 3099 13407 3157 13413
rect 5258 13404 5264 13416
rect 5316 13404 5322 13456
rect 5439 13447 5497 13453
rect 5439 13413 5451 13447
rect 5485 13413 5497 13447
rect 8202 13444 8208 13456
rect 8163 13416 8208 13444
rect 5439 13407 5497 13413
rect 3012 13379 3070 13385
rect 3012 13345 3024 13379
rect 3058 13376 3070 13379
rect 3326 13376 3332 13388
rect 3058 13348 3332 13376
rect 3058 13345 3070 13348
rect 3012 13339 3070 13345
rect 3326 13336 3332 13348
rect 3384 13336 3390 13388
rect 4132 13379 4190 13385
rect 4132 13345 4144 13379
rect 4178 13376 4190 13379
rect 4246 13376 4252 13388
rect 4178 13348 4252 13376
rect 4178 13345 4190 13348
rect 4132 13339 4190 13345
rect 4246 13336 4252 13348
rect 4304 13336 4310 13388
rect 4982 13336 4988 13388
rect 5040 13376 5046 13388
rect 5454 13376 5482 13407
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 10042 13444 10048 13456
rect 10003 13416 10048 13444
rect 10042 13404 10048 13416
rect 10100 13404 10106 13456
rect 10594 13444 10600 13456
rect 10555 13416 10600 13444
rect 10594 13404 10600 13416
rect 10652 13404 10658 13456
rect 11422 13376 11428 13388
rect 5040 13348 5482 13376
rect 11383 13348 11428 13376
rect 5040 13336 5046 13348
rect 11422 13336 11428 13348
rect 11480 13336 11486 13388
rect 5077 13311 5135 13317
rect 5077 13308 5089 13311
rect 4908 13280 5089 13308
rect 4908 13184 4936 13280
rect 5077 13277 5089 13280
rect 5123 13277 5135 13311
rect 6822 13308 6828 13320
rect 6783 13280 6828 13308
rect 5077 13271 5135 13277
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13308 8171 13311
rect 8846 13308 8852 13320
rect 8159 13280 8852 13308
rect 8159 13277 8171 13280
rect 8113 13271 8171 13277
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 9490 13268 9496 13320
rect 9548 13308 9554 13320
rect 9953 13311 10011 13317
rect 9953 13308 9965 13311
rect 9548 13280 9965 13308
rect 9548 13268 9554 13280
rect 9953 13277 9965 13280
rect 9999 13308 10011 13311
rect 11563 13311 11621 13317
rect 11563 13308 11575 13311
rect 9999 13280 11575 13308
rect 9999 13277 10011 13280
rect 9953 13271 10011 13277
rect 11563 13277 11575 13280
rect 11609 13277 11621 13311
rect 11563 13271 11621 13277
rect 8018 13200 8024 13252
rect 8076 13240 8082 13252
rect 8665 13243 8723 13249
rect 8665 13240 8677 13243
rect 8076 13212 8677 13240
rect 8076 13200 8082 13212
rect 8665 13209 8677 13212
rect 8711 13209 8723 13243
rect 8665 13203 8723 13209
rect 4203 13175 4261 13181
rect 4203 13141 4215 13175
rect 4249 13172 4261 13175
rect 4706 13172 4712 13184
rect 4249 13144 4712 13172
rect 4249 13141 4261 13144
rect 4203 13135 4261 13141
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 4890 13172 4896 13184
rect 4851 13144 4896 13172
rect 4890 13132 4896 13144
rect 4948 13132 4954 13184
rect 5994 13172 6000 13184
rect 5955 13144 6000 13172
rect 5994 13132 6000 13144
rect 6052 13132 6058 13184
rect 8754 13132 8760 13184
rect 8812 13172 8818 13184
rect 9033 13175 9091 13181
rect 9033 13172 9045 13175
rect 8812 13144 9045 13172
rect 8812 13132 8818 13144
rect 9033 13141 9045 13144
rect 9079 13141 9091 13175
rect 9033 13135 9091 13141
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 5074 12928 5080 12980
rect 5132 12968 5138 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 5132 12940 6193 12968
rect 5132 12928 5138 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 6181 12931 6239 12937
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 7098 12968 7104 12980
rect 6687 12940 7104 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 4246 12860 4252 12912
rect 4304 12900 4310 12912
rect 4709 12903 4767 12909
rect 4709 12900 4721 12903
rect 4304 12872 4721 12900
rect 4304 12860 4310 12872
rect 4709 12869 4721 12872
rect 4755 12900 4767 12903
rect 5166 12900 5172 12912
rect 4755 12872 5172 12900
rect 4755 12869 4767 12872
rect 4709 12863 4767 12869
rect 5166 12860 5172 12872
rect 5224 12900 5230 12912
rect 5224 12872 5948 12900
rect 5224 12860 5230 12872
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12832 4399 12835
rect 4890 12832 4896 12844
rect 4387 12804 4896 12832
rect 4387 12801 4399 12804
rect 4341 12795 4399 12801
rect 4890 12792 4896 12804
rect 4948 12792 4954 12844
rect 5626 12832 5632 12844
rect 5587 12804 5632 12832
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12733 3939 12767
rect 3881 12727 3939 12733
rect 3513 12699 3571 12705
rect 3513 12665 3525 12699
rect 3559 12696 3571 12699
rect 3896 12696 3924 12727
rect 4154 12724 4160 12776
rect 4212 12764 4218 12776
rect 4212 12736 4257 12764
rect 4212 12724 4218 12736
rect 4522 12724 4528 12776
rect 4580 12764 4586 12776
rect 4982 12764 4988 12776
rect 4580 12736 4988 12764
rect 4580 12724 4586 12736
rect 4982 12724 4988 12736
rect 5040 12724 5046 12776
rect 5920 12764 5948 12872
rect 6196 12832 6224 12931
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 8113 12971 8171 12977
rect 8113 12937 8125 12971
rect 8159 12968 8171 12971
rect 8202 12968 8208 12980
rect 8159 12940 8208 12968
rect 8159 12937 8171 12940
rect 8113 12931 8171 12937
rect 8202 12928 8208 12940
rect 8260 12928 8266 12980
rect 8386 12968 8392 12980
rect 8347 12940 8392 12968
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 11422 12968 11428 12980
rect 11383 12940 11428 12968
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6196 12804 6837 12832
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 8018 12792 8024 12844
rect 8076 12832 8082 12844
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 8076 12804 8953 12832
rect 8076 12792 8082 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 9953 12835 10011 12841
rect 9953 12801 9965 12835
rect 9999 12832 10011 12835
rect 10042 12832 10048 12844
rect 9999 12804 10048 12832
rect 9999 12801 10011 12804
rect 9953 12795 10011 12801
rect 10042 12792 10048 12804
rect 10100 12832 10106 12844
rect 10137 12835 10195 12841
rect 10137 12832 10149 12835
rect 10100 12804 10149 12832
rect 10100 12792 10106 12804
rect 10137 12801 10149 12804
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 7834 12764 7840 12776
rect 5920 12736 7840 12764
rect 7834 12724 7840 12736
rect 7892 12724 7898 12776
rect 10686 12764 10692 12776
rect 10647 12736 10692 12764
rect 10686 12724 10692 12736
rect 10744 12724 10750 12776
rect 4062 12696 4068 12708
rect 3559 12668 4068 12696
rect 3559 12665 3571 12668
rect 3513 12659 3571 12665
rect 4062 12656 4068 12668
rect 4120 12656 4126 12708
rect 4706 12656 4712 12708
rect 4764 12696 4770 12708
rect 5261 12699 5319 12705
rect 5261 12696 5273 12699
rect 4764 12668 5273 12696
rect 4764 12656 4770 12668
rect 5261 12665 5273 12668
rect 5307 12665 5319 12699
rect 5261 12659 5319 12665
rect 5350 12656 5356 12708
rect 5408 12696 5414 12708
rect 5994 12696 6000 12708
rect 5408 12668 6000 12696
rect 5408 12656 5414 12668
rect 5994 12656 6000 12668
rect 6052 12656 6058 12708
rect 8662 12696 8668 12708
rect 8623 12668 8668 12696
rect 8662 12656 8668 12668
rect 8720 12656 8726 12708
rect 8757 12699 8815 12705
rect 8757 12665 8769 12699
rect 8803 12665 8815 12699
rect 8757 12659 8815 12665
rect 3053 12631 3111 12637
rect 3053 12597 3065 12631
rect 3099 12628 3111 12631
rect 3326 12628 3332 12640
rect 3099 12600 3332 12628
rect 3099 12597 3111 12600
rect 3053 12591 3111 12597
rect 3326 12588 3332 12600
rect 3384 12588 3390 12640
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 7193 12631 7251 12637
rect 7193 12628 7205 12631
rect 7156 12600 7205 12628
rect 7156 12588 7162 12600
rect 7193 12597 7205 12600
rect 7239 12597 7251 12631
rect 7742 12628 7748 12640
rect 7703 12600 7748 12628
rect 7193 12591 7251 12597
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 8386 12588 8392 12640
rect 8444 12628 8450 12640
rect 8772 12628 8800 12659
rect 8444 12600 8800 12628
rect 8444 12588 8450 12600
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 3697 12427 3755 12433
rect 3697 12393 3709 12427
rect 3743 12424 3755 12427
rect 4154 12424 4160 12436
rect 3743 12396 4160 12424
rect 3743 12393 3755 12396
rect 3697 12387 3755 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 4706 12424 4712 12436
rect 4667 12396 4712 12424
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 5994 12424 6000 12436
rect 5955 12396 6000 12424
rect 5994 12384 6000 12396
rect 6052 12384 6058 12436
rect 7650 12424 7656 12436
rect 7563 12396 7656 12424
rect 7650 12384 7656 12396
rect 7708 12424 7714 12436
rect 9769 12427 9827 12433
rect 9769 12424 9781 12427
rect 7708 12396 9781 12424
rect 7708 12384 7714 12396
rect 9769 12393 9781 12396
rect 9815 12393 9827 12427
rect 10686 12424 10692 12436
rect 10647 12396 10692 12424
rect 9769 12387 9827 12393
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 106 12316 112 12368
rect 164 12356 170 12368
rect 3099 12359 3157 12365
rect 3099 12356 3111 12359
rect 164 12328 3111 12356
rect 164 12316 170 12328
rect 3099 12325 3111 12328
rect 3145 12325 3157 12359
rect 5074 12356 5080 12368
rect 5035 12328 5080 12356
rect 3099 12319 3157 12325
rect 5074 12316 5080 12328
rect 5132 12316 5138 12368
rect 6641 12359 6699 12365
rect 6641 12325 6653 12359
rect 6687 12356 6699 12359
rect 7006 12356 7012 12368
rect 6687 12328 7012 12356
rect 6687 12325 6699 12328
rect 6641 12319 6699 12325
rect 7006 12316 7012 12328
rect 7064 12356 7070 12368
rect 7742 12356 7748 12368
rect 7064 12328 7748 12356
rect 7064 12316 7070 12328
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 8202 12356 8208 12368
rect 8163 12328 8208 12356
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 8846 12316 8852 12368
rect 8904 12356 8910 12368
rect 9033 12359 9091 12365
rect 9033 12356 9045 12359
rect 8904 12328 9045 12356
rect 8904 12316 8910 12328
rect 9033 12325 9045 12328
rect 9079 12325 9091 12359
rect 9490 12356 9496 12368
rect 9451 12328 9496 12356
rect 9033 12319 9091 12325
rect 9490 12316 9496 12328
rect 9548 12316 9554 12368
rect 2958 12288 2964 12300
rect 2922 12260 2964 12288
rect 2958 12248 2964 12260
rect 3016 12297 3022 12300
rect 3016 12291 3070 12297
rect 3016 12257 3024 12291
rect 3058 12288 3070 12291
rect 9950 12288 9956 12300
rect 3058 12260 4154 12288
rect 9911 12260 9956 12288
rect 3058 12257 3070 12260
rect 3016 12251 3070 12257
rect 3016 12248 3022 12251
rect 4126 12152 4154 12260
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 10134 12288 10140 12300
rect 10095 12260 10140 12288
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 11308 12291 11366 12297
rect 11308 12257 11320 12291
rect 11354 12288 11366 12291
rect 11422 12288 11428 12300
rect 11354 12260 11428 12288
rect 11354 12257 11366 12260
rect 11308 12251 11366 12257
rect 11422 12248 11428 12260
rect 11480 12248 11486 12300
rect 4982 12220 4988 12232
rect 4943 12192 4988 12220
rect 4982 12180 4988 12192
rect 5040 12180 5046 12232
rect 5626 12220 5632 12232
rect 5587 12192 5632 12220
rect 5626 12180 5632 12192
rect 5684 12180 5690 12232
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 6822 12220 6828 12232
rect 6595 12192 6828 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12220 8171 12223
rect 8570 12220 8576 12232
rect 8159 12192 8576 12220
rect 8159 12189 8171 12192
rect 8113 12183 8171 12189
rect 8570 12180 8576 12192
rect 8628 12220 8634 12232
rect 8628 12192 11059 12220
rect 8628 12180 8634 12192
rect 7101 12155 7159 12161
rect 7101 12152 7113 12155
rect 4126 12124 7113 12152
rect 7101 12121 7113 12124
rect 7147 12152 7159 12155
rect 8018 12152 8024 12164
rect 7147 12124 8024 12152
rect 7147 12121 7159 12124
rect 7101 12115 7159 12121
rect 8018 12112 8024 12124
rect 8076 12112 8082 12164
rect 8665 12155 8723 12161
rect 8665 12121 8677 12155
rect 8711 12152 8723 12155
rect 8754 12152 8760 12164
rect 8711 12124 8760 12152
rect 8711 12121 8723 12124
rect 8665 12115 8723 12121
rect 8754 12112 8760 12124
rect 8812 12112 8818 12164
rect 11031 12152 11059 12192
rect 11379 12155 11437 12161
rect 11379 12152 11391 12155
rect 11031 12124 11391 12152
rect 11379 12121 11391 12124
rect 11425 12121 11437 12155
rect 11379 12115 11437 12121
rect 6638 12044 6644 12096
rect 6696 12084 6702 12096
rect 10318 12084 10324 12096
rect 6696 12056 10324 12084
rect 6696 12044 6702 12056
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 2958 11880 2964 11892
rect 2919 11852 2964 11880
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 4617 11883 4675 11889
rect 4617 11849 4629 11883
rect 4663 11880 4675 11883
rect 4985 11883 5043 11889
rect 4985 11880 4997 11883
rect 4663 11852 4997 11880
rect 4663 11849 4675 11852
rect 4617 11843 4675 11849
rect 4985 11849 4997 11852
rect 5031 11880 5043 11883
rect 5074 11880 5080 11892
rect 5031 11852 5080 11880
rect 5031 11849 5043 11852
rect 4985 11843 5043 11849
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 6549 11883 6607 11889
rect 6549 11849 6561 11883
rect 6595 11880 6607 11883
rect 6822 11880 6828 11892
rect 6595 11852 6828 11880
rect 6595 11849 6607 11852
rect 6549 11843 6607 11849
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 7006 11880 7012 11892
rect 6967 11852 7012 11880
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 7098 11840 7104 11892
rect 7156 11880 7162 11892
rect 7469 11883 7527 11889
rect 7469 11880 7481 11883
rect 7156 11852 7481 11880
rect 7156 11840 7162 11852
rect 7469 11849 7481 11852
rect 7515 11849 7527 11883
rect 7469 11843 7527 11849
rect 8202 11840 8208 11892
rect 8260 11880 8266 11892
rect 8573 11883 8631 11889
rect 8573 11880 8585 11883
rect 8260 11852 8585 11880
rect 8260 11840 8266 11852
rect 8573 11849 8585 11852
rect 8619 11880 8631 11883
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 8619 11852 8861 11880
rect 8619 11849 8631 11852
rect 8573 11843 8631 11849
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 8849 11843 8907 11849
rect 6089 11747 6147 11753
rect 6089 11744 6101 11747
rect 5000 11716 6101 11744
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11676 3479 11679
rect 3510 11676 3516 11688
rect 3467 11648 3516 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11676 4123 11679
rect 4154 11676 4160 11688
rect 4111 11648 4160 11676
rect 4111 11645 4123 11648
rect 4065 11639 4123 11645
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 4246 11608 4252 11620
rect 4207 11580 4252 11608
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 4338 11568 4344 11620
rect 4396 11608 4402 11620
rect 5000 11608 5028 11716
rect 6089 11713 6101 11716
rect 6135 11713 6147 11747
rect 7650 11744 7656 11756
rect 7611 11716 7656 11744
rect 6089 11707 6147 11713
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 5169 11611 5227 11617
rect 5169 11608 5181 11611
rect 4396 11580 5181 11608
rect 4396 11568 4402 11580
rect 5169 11577 5181 11580
rect 5215 11577 5227 11611
rect 5169 11571 5227 11577
rect 5261 11611 5319 11617
rect 5261 11577 5273 11611
rect 5307 11577 5319 11611
rect 5810 11608 5816 11620
rect 5771 11580 5816 11608
rect 5261 11571 5319 11577
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5276 11540 5304 11571
rect 5810 11568 5816 11580
rect 5868 11568 5874 11620
rect 7098 11568 7104 11620
rect 7156 11608 7162 11620
rect 7974 11611 8032 11617
rect 7974 11608 7986 11611
rect 7156 11580 7986 11608
rect 7156 11568 7162 11580
rect 7974 11577 7986 11580
rect 8020 11577 8032 11611
rect 8864 11608 8892 11843
rect 8938 11772 8944 11824
rect 8996 11812 9002 11824
rect 10045 11815 10103 11821
rect 10045 11812 10057 11815
rect 8996 11784 10057 11812
rect 8996 11772 9002 11784
rect 10045 11781 10057 11784
rect 10091 11812 10103 11815
rect 10410 11812 10416 11824
rect 10091 11784 10416 11812
rect 10091 11781 10103 11784
rect 10045 11775 10103 11781
rect 10410 11772 10416 11784
rect 10468 11772 10474 11824
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11744 9551 11747
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 9539 11716 10793 11744
rect 9539 11713 9551 11716
rect 9493 11707 9551 11713
rect 10781 11713 10793 11716
rect 10827 11744 10839 11747
rect 11103 11747 11161 11753
rect 11103 11744 11115 11747
rect 10827 11716 11115 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 11103 11713 11115 11716
rect 11149 11713 11161 11747
rect 11103 11707 11161 11713
rect 11016 11679 11074 11685
rect 11016 11645 11028 11679
rect 11062 11676 11074 11679
rect 11238 11676 11244 11688
rect 11062 11648 11244 11676
rect 11062 11645 11074 11648
rect 11016 11639 11074 11645
rect 11238 11636 11244 11648
rect 11296 11676 11302 11688
rect 11296 11648 11376 11676
rect 11296 11636 11302 11648
rect 9490 11608 9496 11620
rect 8864 11580 9496 11608
rect 7974 11571 8032 11577
rect 9490 11568 9496 11580
rect 9548 11608 9554 11620
rect 9585 11611 9643 11617
rect 9585 11608 9597 11611
rect 9548 11580 9597 11608
rect 9548 11568 9554 11580
rect 9585 11577 9597 11580
rect 9631 11577 9643 11611
rect 9585 11571 9643 11577
rect 9950 11568 9956 11620
rect 10008 11608 10014 11620
rect 10413 11611 10471 11617
rect 10413 11608 10425 11611
rect 10008 11580 10425 11608
rect 10008 11568 10014 11580
rect 10413 11577 10425 11580
rect 10459 11577 10471 11611
rect 10413 11571 10471 11577
rect 11348 11552 11376 11648
rect 11422 11636 11428 11688
rect 11480 11676 11486 11688
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 11480 11648 11805 11676
rect 11480 11636 11486 11648
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 5132 11512 5304 11540
rect 5132 11500 5138 11512
rect 8662 11500 8668 11552
rect 8720 11540 8726 11552
rect 9217 11543 9275 11549
rect 9217 11540 9229 11543
rect 8720 11512 9229 11540
rect 8720 11500 8726 11512
rect 9217 11509 9229 11512
rect 9263 11540 9275 11543
rect 10134 11540 10140 11552
rect 9263 11512 10140 11540
rect 9263 11509 9275 11512
rect 9217 11503 9275 11509
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 11425 11543 11483 11549
rect 11425 11540 11437 11543
rect 11388 11512 11437 11540
rect 11388 11500 11394 11512
rect 11425 11509 11437 11512
rect 11471 11509 11483 11543
rect 11425 11503 11483 11509
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 3605 11339 3663 11345
rect 3605 11305 3617 11339
rect 3651 11336 3663 11339
rect 4154 11336 4160 11348
rect 3651 11308 4160 11336
rect 3651 11305 3663 11308
rect 3605 11299 3663 11305
rect 2406 11200 2412 11212
rect 2367 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 2866 11160 2872 11212
rect 2924 11200 2930 11212
rect 2961 11203 3019 11209
rect 2961 11200 2973 11203
rect 2924 11172 2973 11200
rect 2924 11160 2930 11172
rect 2961 11169 2973 11172
rect 3007 11200 3019 11203
rect 3620 11200 3648 11299
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 4522 11296 4528 11348
rect 4580 11336 4586 11348
rect 4617 11339 4675 11345
rect 4617 11336 4629 11339
rect 4580 11308 4629 11336
rect 4580 11296 4586 11308
rect 4617 11305 4629 11308
rect 4663 11305 4675 11339
rect 4617 11299 4675 11305
rect 5074 11296 5080 11348
rect 5132 11336 5138 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 5132 11308 5181 11336
rect 5132 11296 5138 11308
rect 5169 11305 5181 11308
rect 5215 11305 5227 11339
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 5169 11299 5227 11305
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 9490 11336 9496 11348
rect 9451 11308 9496 11336
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 7098 11228 7104 11280
rect 7156 11268 7162 11280
rect 7606 11271 7664 11277
rect 7606 11268 7618 11271
rect 7156 11240 7618 11268
rect 7156 11228 7162 11240
rect 7606 11237 7618 11240
rect 7652 11237 7664 11271
rect 7606 11231 7664 11237
rect 8110 11228 8116 11280
rect 8168 11268 8174 11280
rect 9861 11271 9919 11277
rect 9861 11268 9873 11271
rect 8168 11240 9873 11268
rect 8168 11228 8174 11240
rect 9861 11237 9873 11240
rect 9907 11268 9919 11271
rect 10226 11268 10232 11280
rect 9907 11240 10232 11268
rect 9907 11237 9919 11240
rect 9861 11231 9919 11237
rect 10226 11228 10232 11240
rect 10284 11228 10290 11280
rect 10410 11268 10416 11280
rect 10371 11240 10416 11268
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 11425 11271 11483 11277
rect 11425 11237 11437 11271
rect 11471 11268 11483 11271
rect 11606 11268 11612 11280
rect 11471 11240 11612 11268
rect 11471 11237 11483 11240
rect 11425 11231 11483 11237
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 3007 11172 3648 11200
rect 6340 11203 6398 11209
rect 3007 11169 3019 11172
rect 2961 11163 3019 11169
rect 6340 11169 6352 11203
rect 6386 11200 6398 11203
rect 6638 11200 6644 11212
rect 6386 11172 6644 11200
rect 6386 11169 6398 11172
rect 6340 11163 6398 11169
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 3142 11132 3148 11144
rect 3103 11104 3148 11132
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 4246 11132 4252 11144
rect 4207 11104 4252 11132
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 7282 11132 7288 11144
rect 7243 11104 7288 11132
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11132 9827 11135
rect 10594 11132 10600 11144
rect 9815 11104 10600 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11132 11391 11135
rect 11974 11132 11980 11144
rect 11379 11104 11980 11132
rect 11379 11101 11391 11104
rect 11333 11095 11391 11101
rect 11974 11092 11980 11104
rect 12032 11092 12038 11144
rect 8754 11024 8760 11076
rect 8812 11064 8818 11076
rect 11885 11067 11943 11073
rect 11885 11064 11897 11067
rect 8812 11036 11897 11064
rect 8812 11024 8818 11036
rect 11885 11033 11897 11036
rect 11931 11033 11943 11067
rect 11885 11027 11943 11033
rect 4154 10956 4160 11008
rect 4212 10996 4218 11008
rect 4982 10996 4988 11008
rect 4212 10968 4988 10996
rect 4212 10956 4218 10968
rect 4982 10956 4988 10968
rect 5040 10996 5046 11008
rect 5445 10999 5503 11005
rect 5445 10996 5457 10999
rect 5040 10968 5457 10996
rect 5040 10956 5046 10968
rect 5445 10965 5457 10968
rect 5491 10965 5503 10999
rect 5445 10959 5503 10965
rect 6411 10999 6469 11005
rect 6411 10965 6423 10999
rect 6457 10996 6469 10999
rect 7926 10996 7932 11008
rect 6457 10968 7932 10996
rect 6457 10965 6469 10968
rect 6411 10959 6469 10965
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 8110 10956 8116 11008
rect 8168 10996 8174 11008
rect 8205 10999 8263 11005
rect 8205 10996 8217 10999
rect 8168 10968 8217 10996
rect 8168 10956 8174 10968
rect 8205 10965 8217 10968
rect 8251 10965 8263 10999
rect 8205 10959 8263 10965
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 2406 10792 2412 10804
rect 2367 10764 2412 10792
rect 2406 10752 2412 10764
rect 2464 10752 2470 10804
rect 2866 10792 2872 10804
rect 2827 10764 2872 10792
rect 2866 10752 2872 10764
rect 2924 10752 2930 10804
rect 3559 10795 3617 10801
rect 3559 10761 3571 10795
rect 3605 10792 3617 10795
rect 4154 10792 4160 10804
rect 3605 10764 4160 10792
rect 3605 10761 3617 10764
rect 3559 10755 3617 10761
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4246 10752 4252 10804
rect 4304 10792 4310 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 4304 10764 5641 10792
rect 4304 10752 4310 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 5629 10755 5687 10761
rect 6365 10795 6423 10801
rect 6365 10761 6377 10795
rect 6411 10792 6423 10795
rect 6638 10792 6644 10804
rect 6411 10764 6644 10792
rect 6411 10761 6423 10764
rect 6365 10755 6423 10761
rect 6638 10752 6644 10764
rect 6696 10792 6702 10804
rect 7006 10792 7012 10804
rect 6696 10764 7012 10792
rect 6696 10752 6702 10764
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7285 10795 7343 10801
rect 7285 10792 7297 10795
rect 7156 10764 7297 10792
rect 7156 10752 7162 10764
rect 7285 10761 7297 10764
rect 7331 10761 7343 10795
rect 10226 10792 10232 10804
rect 10187 10764 10232 10792
rect 7285 10755 7343 10761
rect 10226 10752 10232 10764
rect 10284 10752 10290 10804
rect 10594 10792 10600 10804
rect 10555 10764 10600 10792
rect 10594 10752 10600 10764
rect 10652 10792 10658 10804
rect 10919 10795 10977 10801
rect 10919 10792 10931 10795
rect 10652 10764 10931 10792
rect 10652 10752 10658 10764
rect 10919 10761 10931 10764
rect 10965 10761 10977 10795
rect 11606 10792 11612 10804
rect 11567 10764 11612 10792
rect 10919 10755 10977 10761
rect 11606 10752 11612 10764
rect 11664 10752 11670 10804
rect 8389 10727 8447 10733
rect 8389 10693 8401 10727
rect 8435 10724 8447 10727
rect 9125 10727 9183 10733
rect 9125 10724 9137 10727
rect 8435 10696 9137 10724
rect 8435 10693 8447 10696
rect 8389 10687 8447 10693
rect 9125 10693 9137 10696
rect 9171 10724 9183 10727
rect 9398 10724 9404 10736
rect 9171 10696 9404 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 9398 10684 9404 10696
rect 9456 10724 9462 10736
rect 11624 10724 11652 10752
rect 9456 10696 11652 10724
rect 9456 10684 9462 10696
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 3200 10628 4154 10656
rect 3200 10616 3206 10628
rect 3488 10591 3546 10597
rect 3488 10557 3500 10591
rect 3534 10588 3546 10591
rect 4126 10588 4154 10628
rect 7282 10616 7288 10668
rect 7340 10656 7346 10668
rect 8665 10659 8723 10665
rect 8665 10656 8677 10659
rect 7340 10628 8677 10656
rect 7340 10616 7346 10628
rect 8665 10625 8677 10628
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10656 10011 10659
rect 10410 10656 10416 10668
rect 9999 10628 10416 10656
rect 9999 10625 10011 10628
rect 9953 10619 10011 10625
rect 10410 10616 10416 10628
rect 10468 10616 10474 10668
rect 4430 10588 4436 10600
rect 3534 10560 4016 10588
rect 4126 10560 4436 10588
rect 3534 10557 3546 10560
rect 3488 10551 3546 10557
rect 3988 10461 4016 10560
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10588 7527 10591
rect 7558 10588 7564 10600
rect 7515 10560 7564 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 7558 10548 7564 10560
rect 7616 10548 7622 10600
rect 10870 10597 10876 10600
rect 10848 10591 10876 10597
rect 10848 10588 10860 10591
rect 10783 10560 10860 10588
rect 10848 10557 10860 10560
rect 10928 10588 10934 10600
rect 11241 10591 11299 10597
rect 11241 10588 11253 10591
rect 10928 10560 11253 10588
rect 10848 10551 10876 10557
rect 10870 10548 10876 10551
rect 10928 10548 10934 10560
rect 11241 10557 11253 10560
rect 11287 10557 11299 10591
rect 11241 10551 11299 10557
rect 4341 10523 4399 10529
rect 4341 10489 4353 10523
rect 4387 10520 4399 10523
rect 4522 10520 4528 10532
rect 4387 10492 4528 10520
rect 4387 10489 4399 10492
rect 4341 10483 4399 10489
rect 4522 10480 4528 10492
rect 4580 10520 4586 10532
rect 4754 10523 4812 10529
rect 4754 10520 4766 10523
rect 4580 10492 4766 10520
rect 4580 10480 4586 10492
rect 4754 10489 4766 10492
rect 4800 10489 4812 10523
rect 4754 10483 4812 10489
rect 7098 10480 7104 10532
rect 7156 10520 7162 10532
rect 7790 10523 7848 10529
rect 7790 10520 7802 10523
rect 7156 10492 7802 10520
rect 7156 10480 7162 10492
rect 7790 10489 7802 10492
rect 7836 10489 7848 10523
rect 9306 10520 9312 10532
rect 9267 10492 9312 10520
rect 7790 10483 7848 10489
rect 9306 10480 9312 10492
rect 9364 10480 9370 10532
rect 9398 10480 9404 10532
rect 9456 10520 9462 10532
rect 9456 10492 9501 10520
rect 9456 10480 9462 10492
rect 3973 10455 4031 10461
rect 3973 10421 3985 10455
rect 4019 10452 4031 10455
rect 4062 10452 4068 10464
rect 4019 10424 4068 10452
rect 4019 10421 4031 10424
rect 3973 10415 4031 10421
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 5350 10452 5356 10464
rect 5311 10424 5356 10452
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 11974 10452 11980 10464
rect 11935 10424 11980 10452
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 3099 10251 3157 10257
rect 3099 10217 3111 10251
rect 3145 10248 3157 10251
rect 4338 10248 4344 10260
rect 3145 10220 4344 10248
rect 3145 10217 3157 10220
rect 3099 10211 3157 10217
rect 4338 10208 4344 10220
rect 4396 10208 4402 10260
rect 4430 10208 4436 10260
rect 4488 10248 4494 10260
rect 5077 10251 5135 10257
rect 5077 10248 5089 10251
rect 4488 10220 5089 10248
rect 4488 10208 4494 10220
rect 5077 10217 5089 10220
rect 5123 10217 5135 10251
rect 5077 10211 5135 10217
rect 7098 10208 7104 10260
rect 7156 10248 7162 10260
rect 7466 10248 7472 10260
rect 7156 10220 7472 10248
rect 7156 10208 7162 10220
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 9306 10248 9312 10260
rect 9267 10220 9312 10248
rect 9306 10208 9312 10220
rect 9364 10248 9370 10260
rect 9815 10251 9873 10257
rect 9815 10248 9827 10251
rect 9364 10220 9827 10248
rect 9364 10208 9370 10220
rect 9815 10217 9827 10220
rect 9861 10217 9873 10251
rect 9815 10211 9873 10217
rect 5350 10140 5356 10192
rect 5408 10180 5414 10192
rect 5445 10183 5503 10189
rect 5445 10180 5457 10183
rect 5408 10152 5457 10180
rect 5408 10140 5414 10152
rect 5445 10149 5457 10152
rect 5491 10149 5503 10183
rect 5445 10143 5503 10149
rect 8110 10140 8116 10192
rect 8168 10180 8174 10192
rect 8205 10183 8263 10189
rect 8205 10180 8217 10183
rect 8168 10152 8217 10180
rect 8168 10140 8174 10152
rect 8205 10149 8217 10152
rect 8251 10149 8263 10183
rect 8754 10180 8760 10192
rect 8715 10152 8760 10180
rect 8205 10143 8263 10149
rect 8754 10140 8760 10152
rect 8812 10140 8818 10192
rect 4300 10115 4358 10121
rect 4300 10081 4312 10115
rect 4346 10112 4358 10115
rect 4706 10112 4712 10124
rect 4346 10084 4712 10112
rect 4346 10081 4358 10084
rect 4300 10075 4358 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 9585 10115 9643 10121
rect 9585 10081 9597 10115
rect 9631 10112 9643 10115
rect 9674 10112 9680 10124
rect 9631 10084 9680 10112
rect 9631 10081 9643 10084
rect 9585 10075 9643 10081
rect 9674 10072 9680 10084
rect 9732 10112 9738 10124
rect 10042 10112 10048 10124
rect 9732 10084 10048 10112
rect 9732 10072 9738 10084
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4387 10047 4445 10053
rect 4387 10044 4399 10047
rect 4028 10016 4399 10044
rect 4028 10004 4034 10016
rect 4387 10013 4399 10016
rect 4433 10044 4445 10047
rect 5353 10047 5411 10053
rect 5353 10044 5365 10047
rect 4433 10016 5365 10044
rect 4433 10013 4445 10016
rect 4387 10007 4445 10013
rect 5353 10013 5365 10016
rect 5399 10013 5411 10047
rect 5626 10044 5632 10056
rect 5587 10016 5632 10044
rect 5353 10007 5411 10013
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 6822 10044 6828 10056
rect 6783 10016 6828 10044
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 8113 10047 8171 10053
rect 8113 10044 8125 10047
rect 7984 10016 8125 10044
rect 7984 10004 7990 10016
rect 8113 10013 8125 10016
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 2590 9936 2596 9988
rect 2648 9976 2654 9988
rect 8018 9976 8024 9988
rect 2648 9948 8024 9976
rect 2648 9936 2654 9948
rect 8018 9936 8024 9948
rect 8076 9936 8082 9988
rect 2869 9911 2927 9917
rect 2869 9877 2881 9911
rect 2915 9908 2927 9911
rect 2958 9908 2964 9920
rect 2915 9880 2964 9908
rect 2915 9877 2927 9880
rect 2869 9871 2927 9877
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 4522 9868 4528 9920
rect 4580 9908 4586 9920
rect 4709 9911 4767 9917
rect 4709 9908 4721 9911
rect 4580 9880 4721 9908
rect 4580 9868 4586 9880
rect 4709 9877 4721 9880
rect 4755 9877 4767 9911
rect 4709 9871 4767 9877
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 7837 9911 7895 9917
rect 7837 9908 7849 9911
rect 7616 9880 7849 9908
rect 7616 9868 7622 9880
rect 7837 9877 7849 9880
rect 7883 9877 7895 9911
rect 7837 9871 7895 9877
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 3970 9704 3976 9716
rect 3931 9676 3976 9704
rect 3970 9664 3976 9676
rect 4028 9664 4034 9716
rect 4706 9704 4712 9716
rect 4619 9676 4712 9704
rect 4706 9664 4712 9676
rect 4764 9704 4770 9716
rect 6086 9704 6092 9716
rect 4764 9676 6092 9704
rect 4764 9664 4770 9676
rect 6086 9664 6092 9676
rect 6144 9664 6150 9716
rect 8110 9704 8116 9716
rect 8071 9676 8116 9704
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8527 9707 8585 9713
rect 8527 9673 8539 9707
rect 8573 9704 8585 9707
rect 11974 9704 11980 9716
rect 8573 9676 11980 9704
rect 8573 9673 8585 9676
rect 8527 9667 8585 9673
rect 11974 9664 11980 9676
rect 12032 9664 12038 9716
rect 2682 9596 2688 9648
rect 2740 9636 2746 9648
rect 5810 9636 5816 9648
rect 2740 9608 5672 9636
rect 5771 9608 5816 9636
rect 2740 9596 2746 9608
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 3234 9568 3240 9580
rect 2464 9540 3240 9568
rect 2464 9528 2470 9540
rect 3234 9528 3240 9540
rect 3292 9568 3298 9580
rect 5442 9568 5448 9580
rect 3292 9540 5448 9568
rect 3292 9528 3298 9540
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5644 9568 5672 9608
rect 5810 9596 5816 9608
rect 5868 9596 5874 9648
rect 7926 9596 7932 9648
rect 7984 9636 7990 9648
rect 9217 9639 9275 9645
rect 9217 9636 9229 9639
rect 7984 9608 9229 9636
rect 7984 9596 7990 9608
rect 9217 9605 9229 9608
rect 9263 9605 9275 9639
rect 9217 9599 9275 9605
rect 7374 9568 7380 9580
rect 5644 9540 7380 9568
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 7558 9568 7564 9580
rect 7519 9540 7564 9568
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 8662 9568 8668 9580
rect 7668 9540 8668 9568
rect 4208 9503 4266 9509
rect 4208 9469 4220 9503
rect 4254 9500 4266 9503
rect 5074 9500 5080 9512
rect 4254 9472 5080 9500
rect 4254 9469 4266 9472
rect 4208 9463 4266 9469
rect 5074 9460 5080 9472
rect 5132 9460 5138 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 3697 9435 3755 9441
rect 3697 9401 3709 9435
rect 3743 9432 3755 9435
rect 4295 9435 4353 9441
rect 4295 9432 4307 9435
rect 3743 9404 4307 9432
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 4295 9401 4307 9404
rect 4341 9432 4353 9435
rect 5261 9435 5319 9441
rect 5261 9432 5273 9435
rect 4341 9404 5273 9432
rect 4341 9401 4353 9404
rect 4295 9395 4353 9401
rect 5261 9401 5273 9404
rect 5307 9401 5319 9435
rect 5261 9395 5319 9401
rect 5350 9392 5356 9444
rect 5408 9432 5414 9444
rect 6549 9435 6607 9441
rect 6549 9432 6561 9435
rect 5408 9404 5453 9432
rect 5638 9404 6561 9432
rect 5408 9392 5414 9404
rect 2958 9364 2964 9376
rect 2919 9336 2964 9364
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 5074 9364 5080 9376
rect 5035 9336 5080 9364
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 5638 9364 5666 9404
rect 6549 9401 6561 9404
rect 6595 9432 6607 9435
rect 6840 9432 6868 9463
rect 7098 9460 7104 9512
rect 7156 9500 7162 9512
rect 7285 9503 7343 9509
rect 7285 9500 7297 9503
rect 7156 9472 7297 9500
rect 7156 9460 7162 9472
rect 7285 9469 7297 9472
rect 7331 9500 7343 9503
rect 7668 9500 7696 9540
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 8478 9509 8484 9512
rect 8456 9503 8484 9509
rect 8456 9500 8468 9503
rect 7331 9472 7696 9500
rect 8391 9472 8468 9500
rect 7331 9469 7343 9472
rect 7285 9463 7343 9469
rect 8456 9469 8468 9472
rect 8536 9500 8542 9512
rect 8536 9472 8708 9500
rect 8456 9463 8484 9469
rect 8478 9460 8484 9463
rect 8536 9460 8542 9472
rect 7190 9432 7196 9444
rect 6595 9404 7196 9432
rect 6595 9401 6607 9404
rect 6549 9395 6607 9401
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 8680 9376 8708 9472
rect 5500 9336 5666 9364
rect 6273 9367 6331 9373
rect 5500 9324 5506 9336
rect 6273 9333 6285 9367
rect 6319 9364 6331 9367
rect 7098 9364 7104 9376
rect 6319 9336 7104 9364
rect 6319 9333 6331 9336
rect 6273 9327 6331 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 8849 9367 8907 9373
rect 8849 9364 8861 9367
rect 8720 9336 8861 9364
rect 8720 9324 8726 9336
rect 8849 9333 8861 9336
rect 8895 9333 8907 9367
rect 9674 9364 9680 9376
rect 9635 9336 9680 9364
rect 8849 9327 8907 9333
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 5408 9132 5641 9160
rect 5408 9120 5414 9132
rect 5629 9129 5641 9132
rect 5675 9160 5687 9163
rect 5997 9163 6055 9169
rect 5997 9160 6009 9163
rect 5675 9132 6009 9160
rect 5675 9129 5687 9132
rect 5629 9123 5687 9129
rect 5997 9129 6009 9132
rect 6043 9129 6055 9163
rect 5997 9123 6055 9129
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 8570 9160 8576 9172
rect 7432 9132 8576 9160
rect 7432 9120 7438 9132
rect 8570 9120 8576 9132
rect 8628 9160 8634 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 8628 9132 8953 9160
rect 8628 9120 8634 9132
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 8941 9123 8999 9129
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 6178 9092 6184 9104
rect 4120 9064 6184 9092
rect 4120 9052 4126 9064
rect 6178 9052 6184 9064
rect 6236 9092 6242 9104
rect 7282 9092 7288 9104
rect 6236 9064 6592 9092
rect 7243 9064 7288 9092
rect 6236 9052 6242 9064
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 4430 9024 4436 9036
rect 3568 8996 4436 9024
rect 3568 8984 3574 8996
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 4706 9024 4712 9036
rect 4667 8996 4712 9024
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 6564 9033 6592 9064
rect 7282 9052 7288 9064
rect 7340 9052 7346 9104
rect 7558 9052 7564 9104
rect 7616 9092 7622 9104
rect 9674 9092 9680 9104
rect 7616 9064 9680 9092
rect 7616 9052 7622 9064
rect 9674 9052 9680 9064
rect 9732 9052 9738 9104
rect 6549 9027 6607 9033
rect 6549 8993 6561 9027
rect 6595 8993 6607 9027
rect 7098 9024 7104 9036
rect 7059 8996 7104 9024
rect 6549 8987 6607 8993
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 8113 9027 8171 9033
rect 8113 8993 8125 9027
rect 8159 9024 8171 9027
rect 8294 9024 8300 9036
rect 8159 8996 8300 9024
rect 8159 8993 8171 8996
rect 8113 8987 8171 8993
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 4798 8956 4804 8968
rect 4759 8928 4804 8956
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8956 6515 8959
rect 7116 8956 7144 8984
rect 6503 8928 7144 8956
rect 6503 8925 6515 8928
rect 6457 8919 6515 8925
rect 8297 8891 8355 8897
rect 8297 8888 8309 8891
rect 5368 8860 8309 8888
rect 5368 8832 5396 8860
rect 8297 8857 8309 8860
rect 8343 8888 8355 8891
rect 8573 8891 8631 8897
rect 8573 8888 8585 8891
rect 8343 8860 8585 8888
rect 8343 8857 8355 8860
rect 8297 8851 8355 8857
rect 8573 8857 8585 8860
rect 8619 8888 8631 8891
rect 8846 8888 8852 8900
rect 8619 8860 8852 8888
rect 8619 8857 8631 8860
rect 8573 8851 8631 8857
rect 8846 8848 8852 8860
rect 8904 8848 8910 8900
rect 5350 8820 5356 8832
rect 5311 8792 5356 8820
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 7653 8823 7711 8829
rect 7653 8789 7665 8823
rect 7699 8820 7711 8823
rect 8202 8820 8208 8832
rect 7699 8792 8208 8820
rect 7699 8789 7711 8792
rect 7653 8783 7711 8789
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 4985 8619 5043 8625
rect 4985 8616 4997 8619
rect 4948 8588 4997 8616
rect 4948 8576 4954 8588
rect 4985 8585 4997 8588
rect 5031 8616 5043 8619
rect 6178 8616 6184 8628
rect 5031 8588 5120 8616
rect 6139 8588 6184 8616
rect 5031 8585 5043 8588
rect 4985 8579 5043 8585
rect 658 8508 664 8560
rect 716 8548 722 8560
rect 4614 8548 4620 8560
rect 716 8520 4620 8548
rect 716 8508 722 8520
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8480 3571 8483
rect 5092 8480 5120 8588
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 8205 8619 8263 8625
rect 8205 8585 8217 8619
rect 8251 8616 8263 8619
rect 8294 8616 8300 8628
rect 8251 8588 8300 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 9950 8548 9956 8560
rect 3559 8452 5120 8480
rect 3559 8449 3571 8452
rect 3513 8443 3571 8449
rect 3896 8421 3924 8452
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8381 3939 8415
rect 3881 8375 3939 8381
rect 4157 8415 4215 8421
rect 4157 8381 4169 8415
rect 4203 8412 4215 8415
rect 4246 8412 4252 8424
rect 4203 8384 4252 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 4246 8372 4252 8384
rect 4304 8412 4310 8424
rect 4706 8412 4712 8424
rect 4304 8384 4712 8412
rect 4304 8372 4310 8384
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 5092 8412 5120 8452
rect 5736 8520 9956 8548
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 5092 8384 5181 8412
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 5350 8372 5356 8424
rect 5408 8412 5414 8424
rect 5629 8415 5687 8421
rect 5629 8412 5641 8415
rect 5408 8384 5641 8412
rect 5408 8372 5414 8384
rect 5629 8381 5641 8384
rect 5675 8381 5687 8415
rect 5629 8375 5687 8381
rect 4338 8344 4344 8356
rect 4299 8316 4344 8344
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 4614 8304 4620 8356
rect 4672 8344 4678 8356
rect 5258 8344 5264 8356
rect 4672 8316 5264 8344
rect 4672 8304 4678 8316
rect 5258 8304 5264 8316
rect 5316 8304 5322 8356
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 4154 8276 4160 8288
rect 4028 8248 4160 8276
rect 4028 8236 4034 8248
rect 4154 8236 4160 8248
rect 4212 8236 4218 8288
rect 4430 8236 4436 8288
rect 4488 8276 4494 8288
rect 4709 8279 4767 8285
rect 4709 8276 4721 8279
rect 4488 8248 4721 8276
rect 4488 8236 4494 8248
rect 4709 8245 4721 8248
rect 4755 8276 4767 8279
rect 5736 8276 5764 8520
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 8202 8480 8208 8492
rect 6871 8452 8208 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 7466 8412 7472 8424
rect 6687 8384 7472 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 5905 8347 5963 8353
rect 5905 8313 5917 8347
rect 5951 8344 5963 8347
rect 7006 8344 7012 8356
rect 5951 8316 7012 8344
rect 5951 8313 5963 8316
rect 5905 8307 5963 8313
rect 7006 8304 7012 8316
rect 7064 8304 7070 8356
rect 7161 8353 7189 8384
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 8570 8412 8576 8424
rect 8531 8384 8576 8412
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 9033 8415 9091 8421
rect 9033 8412 9045 8415
rect 8904 8384 9045 8412
rect 8904 8372 8910 8384
rect 9033 8381 9045 8384
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 7146 8347 7204 8353
rect 7146 8344 7158 8347
rect 7124 8316 7158 8344
rect 7146 8313 7158 8316
rect 7192 8313 7204 8347
rect 7146 8307 7204 8313
rect 4755 8248 5764 8276
rect 4755 8245 4767 8248
rect 4709 8239 4767 8245
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 7745 8279 7803 8285
rect 7745 8276 7757 8279
rect 6696 8248 7757 8276
rect 6696 8236 6702 8248
rect 7745 8245 7757 8248
rect 7791 8245 7803 8279
rect 7745 8239 7803 8245
rect 8202 8236 8208 8288
rect 8260 8276 8266 8288
rect 8665 8279 8723 8285
rect 8665 8276 8677 8279
rect 8260 8248 8677 8276
rect 8260 8236 8266 8248
rect 8665 8245 8677 8248
rect 8711 8245 8723 8279
rect 8665 8239 8723 8245
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 3237 8075 3295 8081
rect 3237 8041 3249 8075
rect 3283 8072 3295 8075
rect 3697 8075 3755 8081
rect 3697 8072 3709 8075
rect 3283 8044 3709 8072
rect 3283 8041 3295 8044
rect 3237 8035 3295 8041
rect 3697 8041 3709 8044
rect 3743 8072 3755 8075
rect 3970 8072 3976 8084
rect 3743 8044 3976 8072
rect 3743 8041 3755 8044
rect 3697 8035 3755 8041
rect 3970 8032 3976 8044
rect 4028 8072 4034 8084
rect 4246 8072 4252 8084
rect 4028 8044 4252 8072
rect 4028 8032 4034 8044
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4798 8072 4804 8084
rect 4759 8044 4804 8072
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 7558 8072 7564 8084
rect 5092 8044 7564 8072
rect 3050 7964 3056 8016
rect 3108 8004 3114 8016
rect 5092 8004 5120 8044
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7708 8044 7757 8072
rect 7708 8032 7714 8044
rect 7745 8041 7757 8044
rect 7791 8072 7803 8075
rect 9769 8075 9827 8081
rect 9769 8072 9781 8075
rect 7791 8044 9781 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 9769 8041 9781 8044
rect 9815 8041 9827 8075
rect 9769 8035 9827 8041
rect 6086 8004 6092 8016
rect 3108 7976 5120 8004
rect 5184 7976 6092 8004
rect 3108 7964 3114 7976
rect 4982 7896 4988 7948
rect 5040 7936 5046 7948
rect 5184 7945 5212 7976
rect 6086 7964 6092 7976
rect 6144 7964 6150 8016
rect 6638 8004 6644 8016
rect 6599 7976 6644 8004
rect 6638 7964 6644 7976
rect 6696 7964 6702 8016
rect 8202 8004 8208 8016
rect 8163 7976 8208 8004
rect 8202 7964 8208 7976
rect 8260 7964 8266 8016
rect 8846 7964 8852 8016
rect 8904 8004 8910 8016
rect 8904 7976 10180 8004
rect 8904 7964 8910 7976
rect 5169 7939 5227 7945
rect 5169 7936 5181 7939
rect 5040 7908 5181 7936
rect 5040 7896 5046 7908
rect 5169 7905 5181 7908
rect 5215 7905 5227 7939
rect 5350 7936 5356 7948
rect 5263 7908 5356 7936
rect 5169 7899 5227 7905
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 9950 7936 9956 7948
rect 9911 7908 9956 7936
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 10152 7945 10180 7976
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7905 10195 7939
rect 10137 7899 10195 7905
rect 4430 7828 4436 7880
rect 4488 7868 4494 7880
rect 5368 7868 5396 7896
rect 4488 7840 5396 7868
rect 5629 7871 5687 7877
rect 4488 7828 4494 7840
rect 5629 7837 5641 7871
rect 5675 7868 5687 7871
rect 6086 7868 6092 7880
rect 5675 7840 6092 7868
rect 5675 7837 5687 7840
rect 5629 7831 5687 7837
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 6822 7868 6828 7880
rect 6595 7840 6828 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7868 8171 7871
rect 8478 7868 8484 7880
rect 8159 7840 8484 7868
rect 8159 7837 8171 7840
rect 8113 7831 8171 7837
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 9306 7868 9312 7880
rect 8803 7840 9312 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 4154 7760 4160 7812
rect 4212 7800 4218 7812
rect 7101 7803 7159 7809
rect 7101 7800 7113 7803
rect 4212 7772 7113 7800
rect 4212 7760 4218 7772
rect 7101 7769 7113 7772
rect 7147 7800 7159 7803
rect 9858 7800 9864 7812
rect 7147 7772 9864 7800
rect 7147 7769 7159 7772
rect 7101 7763 7159 7769
rect 9858 7760 9864 7772
rect 9916 7760 9922 7812
rect 9490 7732 9496 7744
rect 9451 7704 9496 7732
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 6638 7488 6644 7540
rect 6696 7528 6702 7540
rect 7009 7531 7067 7537
rect 7009 7528 7021 7531
rect 6696 7500 7021 7528
rect 6696 7488 6702 7500
rect 7009 7497 7021 7500
rect 7055 7497 7067 7531
rect 7009 7491 7067 7497
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8573 7531 8631 7537
rect 8573 7528 8585 7531
rect 8260 7500 8585 7528
rect 8260 7488 8266 7500
rect 8573 7497 8585 7500
rect 8619 7528 8631 7531
rect 8849 7531 8907 7537
rect 8849 7528 8861 7531
rect 8619 7500 8861 7528
rect 8619 7497 8631 7500
rect 8573 7491 8631 7497
rect 8849 7497 8861 7500
rect 8895 7497 8907 7531
rect 8849 7491 8907 7497
rect 6549 7463 6607 7469
rect 6549 7429 6561 7463
rect 6595 7460 6607 7463
rect 6822 7460 6828 7472
rect 6595 7432 6828 7460
rect 6595 7429 6607 7432
rect 6549 7423 6607 7429
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 4062 7392 4068 7404
rect 3099 7364 4068 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 3436 7333 3464 7364
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7392 4767 7395
rect 4798 7392 4804 7404
rect 4755 7364 4804 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 7650 7392 7656 7404
rect 7611 7364 7656 7392
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 3421 7327 3479 7333
rect 3421 7293 3433 7327
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3697 7327 3755 7333
rect 3697 7293 3709 7327
rect 3743 7324 3755 7327
rect 3970 7324 3976 7336
rect 3743 7296 3976 7324
rect 3743 7293 3755 7296
rect 3697 7287 3755 7293
rect 3970 7284 3976 7296
rect 4028 7284 4034 7336
rect 4522 7284 4528 7336
rect 4580 7324 4586 7336
rect 4617 7327 4675 7333
rect 4617 7324 4629 7327
rect 4580 7296 4629 7324
rect 4580 7284 4586 7296
rect 4617 7293 4629 7296
rect 4663 7324 4675 7327
rect 4663 7296 5114 7324
rect 4663 7293 4675 7296
rect 4617 7287 4675 7293
rect 3881 7259 3939 7265
rect 3881 7225 3893 7259
rect 3927 7256 3939 7259
rect 4890 7256 4896 7268
rect 3927 7228 4896 7256
rect 3927 7225 3939 7228
rect 3881 7219 3939 7225
rect 4890 7216 4896 7228
rect 4948 7216 4954 7268
rect 5086 7265 5114 7296
rect 5071 7259 5129 7265
rect 5071 7225 5083 7259
rect 5117 7256 5129 7259
rect 5442 7256 5448 7268
rect 5117 7228 5448 7256
rect 5117 7225 5129 7228
rect 5071 7219 5129 7225
rect 5442 7216 5448 7228
rect 5500 7216 5506 7268
rect 7974 7259 8032 7265
rect 7974 7256 7986 7259
rect 7484 7228 7986 7256
rect 7484 7200 7512 7228
rect 7974 7225 7986 7228
rect 8020 7225 8032 7259
rect 8864 7256 8892 7491
rect 9950 7488 9956 7540
rect 10008 7528 10014 7540
rect 10413 7531 10471 7537
rect 10413 7528 10425 7531
rect 10008 7500 10425 7528
rect 10008 7488 10014 7500
rect 10413 7497 10425 7500
rect 10459 7497 10471 7531
rect 10413 7491 10471 7497
rect 8938 7420 8944 7472
rect 8996 7460 9002 7472
rect 9217 7463 9275 7469
rect 9217 7460 9229 7463
rect 8996 7432 9229 7460
rect 8996 7420 9002 7432
rect 9217 7429 9229 7432
rect 9263 7429 9275 7463
rect 9217 7423 9275 7429
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 11425 7463 11483 7469
rect 11425 7460 11437 7463
rect 9732 7432 11437 7460
rect 9732 7420 9738 7432
rect 9490 7392 9496 7404
rect 9403 7364 9496 7392
rect 9490 7352 9496 7364
rect 9548 7392 9554 7404
rect 11103 7395 11161 7401
rect 11103 7392 11115 7395
rect 9548 7364 11115 7392
rect 9548 7352 9554 7364
rect 11103 7361 11115 7364
rect 11149 7361 11161 7395
rect 11103 7355 11161 7361
rect 11016 7327 11074 7333
rect 11016 7293 11028 7327
rect 11062 7324 11074 7327
rect 11256 7324 11284 7432
rect 11425 7429 11437 7432
rect 11471 7429 11483 7463
rect 11425 7423 11483 7429
rect 11062 7296 11284 7324
rect 11062 7293 11074 7296
rect 11016 7287 11074 7293
rect 9490 7256 9496 7268
rect 8864 7228 9496 7256
rect 7974 7219 8032 7225
rect 9490 7216 9496 7228
rect 9548 7256 9554 7268
rect 9585 7259 9643 7265
rect 9585 7256 9597 7259
rect 9548 7228 9597 7256
rect 9548 7216 9554 7228
rect 9585 7225 9597 7228
rect 9631 7225 9643 7259
rect 9585 7219 9643 7225
rect 9766 7216 9772 7268
rect 9824 7256 9830 7268
rect 10137 7259 10195 7265
rect 10137 7256 10149 7259
rect 9824 7228 10149 7256
rect 9824 7216 9830 7228
rect 10137 7225 10149 7228
rect 10183 7225 10195 7259
rect 10137 7219 10195 7225
rect 4249 7191 4307 7197
rect 4249 7157 4261 7191
rect 4295 7188 4307 7191
rect 4430 7188 4436 7200
rect 4295 7160 4436 7188
rect 4295 7157 4307 7160
rect 4249 7151 4307 7157
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 5626 7188 5632 7200
rect 5587 7160 5632 7188
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 7466 7188 7472 7200
rect 7427 7160 7472 7188
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 4338 6944 4344 6996
rect 4396 6984 4402 6996
rect 6457 6987 6515 6993
rect 6457 6984 6469 6987
rect 4396 6956 6469 6984
rect 4396 6944 4402 6956
rect 6457 6953 6469 6956
rect 6503 6953 6515 6987
rect 9490 6984 9496 6996
rect 9451 6956 9496 6984
rect 6457 6947 6515 6953
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 2682 6916 2688 6928
rect 2424 6888 2688 6916
rect 2424 6857 2452 6888
rect 2682 6876 2688 6888
rect 2740 6876 2746 6928
rect 4982 6916 4988 6928
rect 4943 6888 4988 6916
rect 4982 6876 4988 6888
rect 5040 6876 5046 6928
rect 5442 6876 5448 6928
rect 5500 6916 5506 6928
rect 5582 6919 5640 6925
rect 5582 6916 5594 6919
rect 5500 6888 5594 6916
rect 5500 6876 5506 6888
rect 5582 6885 5594 6888
rect 5628 6885 5640 6919
rect 5582 6879 5640 6885
rect 7558 6876 7564 6928
rect 7616 6916 7622 6928
rect 7790 6919 7848 6925
rect 7790 6916 7802 6919
rect 7616 6888 7802 6916
rect 7616 6876 7622 6888
rect 7790 6885 7802 6888
rect 7836 6885 7848 6919
rect 7790 6879 7848 6885
rect 9861 6919 9919 6925
rect 9861 6885 9873 6919
rect 9907 6916 9919 6919
rect 9950 6916 9956 6928
rect 9907 6888 9956 6916
rect 9907 6885 9919 6888
rect 9861 6879 9919 6885
rect 9950 6876 9956 6888
rect 10008 6876 10014 6928
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6817 2467 6851
rect 2409 6811 2467 6817
rect 2498 6808 2504 6860
rect 2556 6848 2562 6860
rect 2961 6851 3019 6857
rect 2961 6848 2973 6851
rect 2556 6820 2973 6848
rect 2556 6808 2562 6820
rect 2961 6817 2973 6820
rect 3007 6848 3019 6851
rect 3970 6848 3976 6860
rect 3007 6820 3976 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6817 4307 6851
rect 4249 6811 4307 6817
rect 3142 6780 3148 6792
rect 3103 6752 3148 6780
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 4264 6780 4292 6811
rect 4890 6808 4896 6860
rect 4948 6848 4954 6860
rect 5261 6851 5319 6857
rect 5261 6848 5273 6851
rect 4948 6820 5273 6848
rect 4948 6808 4954 6820
rect 5261 6817 5273 6820
rect 5307 6848 5319 6851
rect 6178 6848 6184 6860
rect 5307 6820 6184 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 7006 6808 7012 6860
rect 7064 6848 7070 6860
rect 7469 6851 7527 6857
rect 7469 6848 7481 6851
rect 7064 6820 7481 6848
rect 7064 6808 7070 6820
rect 7469 6817 7481 6820
rect 7515 6848 7527 6851
rect 8202 6848 8208 6860
rect 7515 6820 8208 6848
rect 7515 6817 7527 6820
rect 7469 6811 7527 6817
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 4522 6780 4528 6792
rect 4264 6752 4528 6780
rect 4522 6740 4528 6752
rect 4580 6780 4586 6792
rect 9582 6780 9588 6792
rect 4580 6752 9588 6780
rect 4580 6740 4586 6752
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 9858 6740 9864 6792
rect 9916 6780 9922 6792
rect 10045 6783 10103 6789
rect 10045 6780 10057 6783
rect 9916 6752 10057 6780
rect 9916 6740 9922 6752
rect 10045 6749 10057 6752
rect 10091 6749 10103 6783
rect 10045 6743 10103 6749
rect 3970 6672 3976 6724
rect 4028 6712 4034 6724
rect 4433 6715 4491 6721
rect 4433 6712 4445 6715
rect 4028 6684 4445 6712
rect 4028 6672 4034 6684
rect 4433 6681 4445 6684
rect 4479 6681 4491 6715
rect 4433 6675 4491 6681
rect 4798 6672 4804 6724
rect 4856 6712 4862 6724
rect 5902 6712 5908 6724
rect 4856 6684 5908 6712
rect 4856 6672 4862 6684
rect 5902 6672 5908 6684
rect 5960 6672 5966 6724
rect 5994 6604 6000 6656
rect 6052 6644 6058 6656
rect 6181 6647 6239 6653
rect 6181 6644 6193 6647
rect 6052 6616 6193 6644
rect 6052 6604 6058 6616
rect 6181 6613 6193 6616
rect 6227 6613 6239 6647
rect 8386 6644 8392 6656
rect 8347 6616 8392 6644
rect 6181 6607 6239 6613
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 8536 6616 8769 6644
rect 8536 6604 8542 6616
rect 8757 6613 8769 6616
rect 8803 6644 8815 6647
rect 9490 6644 9496 6656
rect 8803 6616 9496 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 2498 6440 2504 6452
rect 2363 6412 2504 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 2869 6443 2927 6449
rect 2869 6440 2881 6443
rect 2740 6412 2881 6440
rect 2740 6400 2746 6412
rect 2869 6409 2881 6412
rect 2915 6409 2927 6443
rect 3234 6440 3240 6452
rect 3195 6412 3240 6440
rect 2869 6403 2927 6409
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 4522 6440 4528 6452
rect 4483 6412 4528 6440
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 6178 6440 6184 6452
rect 6139 6412 6184 6440
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 9033 6443 9091 6449
rect 9033 6440 9045 6443
rect 8444 6412 9045 6440
rect 8444 6400 8450 6412
rect 9033 6409 9045 6412
rect 9079 6440 9091 6443
rect 9398 6440 9404 6452
rect 9079 6412 9404 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 9858 6372 9864 6384
rect 9819 6344 9864 6372
rect 9858 6332 9864 6344
rect 9916 6332 9922 6384
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 2547 6307 2605 6313
rect 2547 6304 2559 6307
rect 2372 6276 2559 6304
rect 2372 6264 2378 6276
rect 2547 6273 2559 6276
rect 2593 6273 2605 6307
rect 4154 6304 4160 6316
rect 2547 6267 2605 6273
rect 2976 6276 4160 6304
rect 2406 6236 2412 6248
rect 2370 6208 2412 6236
rect 2406 6196 2412 6208
rect 2464 6245 2470 6248
rect 2464 6239 2518 6245
rect 2464 6205 2472 6239
rect 2506 6236 2518 6239
rect 2976 6236 3004 6276
rect 4154 6264 4160 6276
rect 4212 6264 4218 6316
rect 4338 6264 4344 6316
rect 4396 6304 4402 6316
rect 4985 6307 5043 6313
rect 4985 6304 4997 6307
rect 4396 6276 4997 6304
rect 4396 6264 4402 6276
rect 4985 6273 4997 6276
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 6086 6264 6092 6316
rect 6144 6304 6150 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 6144 6276 7481 6304
rect 6144 6264 6150 6276
rect 7469 6273 7481 6276
rect 7515 6304 7527 6307
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 7515 6276 8677 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 9950 6304 9956 6316
rect 8665 6267 8723 6273
rect 8772 6276 9956 6304
rect 2506 6208 3004 6236
rect 2506 6205 2518 6208
rect 2464 6199 2518 6205
rect 2464 6196 2470 6199
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 3292 6208 3433 6236
rect 3292 6196 3298 6208
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3970 6236 3976 6248
rect 3931 6208 3976 6236
rect 3421 6199 3479 6205
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 8772 6236 8800 6276
rect 9950 6264 9956 6276
rect 10008 6304 10014 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 10008 6276 10241 6304
rect 10008 6264 10014 6276
rect 10229 6273 10241 6276
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 8435 6208 8800 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 4154 6128 4160 6180
rect 4212 6168 4218 6180
rect 5306 6171 5364 6177
rect 5306 6168 5318 6171
rect 4212 6140 4257 6168
rect 4908 6140 5318 6168
rect 4212 6128 4218 6140
rect 4908 6112 4936 6140
rect 5306 6137 5318 6140
rect 5352 6168 5364 6171
rect 5442 6168 5448 6180
rect 5352 6140 5448 6168
rect 5352 6137 5364 6140
rect 5306 6131 5364 6137
rect 5442 6128 5448 6140
rect 5500 6168 5506 6180
rect 6549 6171 6607 6177
rect 6549 6168 6561 6171
rect 5500 6140 6561 6168
rect 5500 6128 5506 6140
rect 6549 6137 6561 6140
rect 6595 6168 6607 6171
rect 7285 6171 7343 6177
rect 7285 6168 7297 6171
rect 6595 6140 7297 6168
rect 6595 6137 6607 6140
rect 6549 6131 6607 6137
rect 7285 6137 7297 6140
rect 7331 6168 7343 6171
rect 7466 6168 7472 6180
rect 7331 6140 7472 6168
rect 7331 6137 7343 6140
rect 7285 6131 7343 6137
rect 7466 6128 7472 6140
rect 7524 6168 7530 6180
rect 7790 6171 7848 6177
rect 7790 6168 7802 6171
rect 7524 6140 7802 6168
rect 7524 6128 7530 6140
rect 7790 6137 7802 6140
rect 7836 6137 7848 6171
rect 9306 6168 9312 6180
rect 9267 6140 9312 6168
rect 7790 6131 7848 6137
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 9398 6128 9404 6180
rect 9456 6168 9462 6180
rect 9456 6140 9501 6168
rect 9456 6128 9462 6140
rect 4890 6100 4896 6112
rect 4851 6072 4896 6100
rect 4890 6060 4896 6072
rect 4948 6060 4954 6112
rect 5902 6100 5908 6112
rect 5863 6072 5908 6100
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 10597 6103 10655 6109
rect 10597 6100 10609 6103
rect 9824 6072 10609 6100
rect 9824 6060 9830 6072
rect 10597 6069 10609 6072
rect 10643 6069 10655 6103
rect 10597 6063 10655 6069
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 2406 5896 2412 5908
rect 2367 5868 2412 5896
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 3970 5896 3976 5908
rect 3559 5868 3976 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 7282 5896 7288 5908
rect 7243 5868 7288 5896
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 8202 5896 8208 5908
rect 8163 5868 8208 5896
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 9306 5896 9312 5908
rect 9267 5868 9312 5896
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 9815 5899 9873 5905
rect 9815 5896 9827 5899
rect 9548 5868 9827 5896
rect 9548 5856 9554 5868
rect 9815 5865 9827 5868
rect 9861 5865 9873 5899
rect 9815 5859 9873 5865
rect 5813 5831 5871 5837
rect 5813 5797 5825 5831
rect 5859 5828 5871 5831
rect 5902 5828 5908 5840
rect 5859 5800 5908 5828
rect 5859 5797 5871 5800
rect 5813 5791 5871 5797
rect 5902 5788 5908 5800
rect 5960 5828 5966 5840
rect 6178 5828 6184 5840
rect 5960 5800 6184 5828
rect 5960 5788 5966 5800
rect 6178 5788 6184 5800
rect 6236 5788 6242 5840
rect 4062 5760 4068 5772
rect 4023 5732 4068 5760
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 4338 5720 4344 5772
rect 4396 5760 4402 5772
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 4396 5732 4537 5760
rect 4396 5720 4402 5732
rect 4525 5729 4537 5732
rect 4571 5760 4583 5763
rect 5350 5760 5356 5772
rect 4571 5732 5356 5760
rect 4571 5729 4583 5732
rect 4525 5723 4583 5729
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 7190 5760 7196 5772
rect 7151 5732 7196 5760
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 7650 5760 7656 5772
rect 7611 5732 7656 5760
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 9674 5760 9680 5772
rect 9732 5769 9738 5772
rect 9732 5763 9770 5769
rect 7800 5732 9680 5760
rect 7800 5720 7806 5732
rect 9674 5720 9680 5732
rect 9758 5729 9770 5763
rect 9732 5723 9770 5729
rect 9732 5720 9738 5723
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 5442 5692 5448 5704
rect 4847 5664 5448 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 5718 5692 5724 5704
rect 5679 5664 5724 5692
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 5810 5652 5816 5704
rect 5868 5692 5874 5704
rect 5997 5695 6055 5701
rect 5997 5692 6009 5695
rect 5868 5664 6009 5692
rect 5868 5652 5874 5664
rect 5997 5661 6009 5664
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 5261 5559 5319 5565
rect 5261 5556 5273 5559
rect 4948 5528 5273 5556
rect 4948 5516 4954 5528
rect 5261 5525 5273 5528
rect 5307 5525 5319 5559
rect 5261 5519 5319 5525
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 4617 5355 4675 5361
rect 4617 5352 4629 5355
rect 4120 5324 4629 5352
rect 4120 5312 4126 5324
rect 4617 5321 4629 5324
rect 4663 5321 4675 5355
rect 4617 5315 4675 5321
rect 5077 5355 5135 5361
rect 5077 5321 5089 5355
rect 5123 5352 5135 5355
rect 5626 5352 5632 5364
rect 5123 5324 5632 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 6178 5352 6184 5364
rect 6139 5324 6184 5352
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 7745 5355 7803 5361
rect 7745 5352 7757 5355
rect 7248 5324 7757 5352
rect 7248 5312 7254 5324
rect 7745 5321 7757 5324
rect 7791 5321 7803 5355
rect 9674 5352 9680 5364
rect 9635 5324 9680 5352
rect 7745 5315 7803 5321
rect 9674 5312 9680 5324
rect 9732 5352 9738 5364
rect 13170 5352 13176 5364
rect 9732 5324 13176 5352
rect 9732 5312 9738 5324
rect 13170 5312 13176 5324
rect 13228 5312 13234 5364
rect 3326 5244 3332 5296
rect 3384 5284 3390 5296
rect 3384 5256 5304 5284
rect 3384 5244 3390 5256
rect 5276 5228 5304 5256
rect 5350 5244 5356 5296
rect 5408 5284 5414 5296
rect 6549 5287 6607 5293
rect 6549 5284 6561 5287
rect 5408 5256 6561 5284
rect 5408 5244 5414 5256
rect 6549 5253 6561 5256
rect 6595 5284 6607 5287
rect 7650 5284 7656 5296
rect 6595 5256 7656 5284
rect 6595 5253 6607 5256
rect 6549 5247 6607 5253
rect 7650 5244 7656 5256
rect 7708 5244 7714 5296
rect 9398 5244 9404 5296
rect 9456 5284 9462 5296
rect 9999 5287 10057 5293
rect 9999 5284 10011 5287
rect 9456 5256 10011 5284
rect 9456 5244 9462 5256
rect 9999 5253 10011 5256
rect 10045 5253 10057 5287
rect 9999 5247 10057 5253
rect 4982 5216 4988 5228
rect 3896 5188 4988 5216
rect 3896 5157 3924 5188
rect 4982 5176 4988 5188
rect 5040 5176 5046 5228
rect 5258 5216 5264 5228
rect 5171 5188 5264 5216
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 5718 5216 5724 5228
rect 5679 5188 5724 5216
rect 5718 5176 5724 5188
rect 5776 5176 5782 5228
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 9033 5219 9091 5225
rect 9033 5216 9045 5219
rect 8812 5188 9045 5216
rect 8812 5176 8818 5188
rect 9033 5185 9045 5188
rect 9079 5216 9091 5219
rect 9306 5216 9312 5228
rect 9079 5188 9312 5216
rect 9079 5185 9091 5188
rect 9033 5179 9091 5185
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 3513 5151 3571 5157
rect 3513 5117 3525 5151
rect 3559 5148 3571 5151
rect 3881 5151 3939 5157
rect 3881 5148 3893 5151
rect 3559 5120 3893 5148
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 3881 5117 3893 5120
rect 3927 5117 3939 5151
rect 3881 5111 3939 5117
rect 3970 5108 3976 5160
rect 4028 5148 4034 5160
rect 4065 5151 4123 5157
rect 4065 5148 4077 5151
rect 4028 5120 4077 5148
rect 4028 5108 4034 5120
rect 4065 5117 4077 5120
rect 4111 5117 4123 5151
rect 4065 5111 4123 5117
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6788 5120 6837 5148
rect 6788 5108 6794 5120
rect 6825 5117 6837 5120
rect 6871 5148 6883 5151
rect 7377 5151 7435 5157
rect 7377 5148 7389 5151
rect 6871 5120 7389 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 7377 5117 7389 5120
rect 7423 5117 7435 5151
rect 7377 5111 7435 5117
rect 9928 5151 9986 5157
rect 9928 5117 9940 5151
rect 9974 5148 9986 5151
rect 10042 5148 10048 5160
rect 9974 5120 10048 5148
rect 9974 5117 9986 5120
rect 9928 5111 9986 5117
rect 10042 5108 10048 5120
rect 10100 5148 10106 5160
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 10100 5120 10333 5148
rect 10100 5108 10106 5120
rect 10321 5117 10333 5120
rect 10367 5117 10379 5151
rect 10321 5111 10379 5117
rect 4341 5083 4399 5089
rect 4341 5049 4353 5083
rect 4387 5080 4399 5083
rect 4706 5080 4712 5092
rect 4387 5052 4712 5080
rect 4387 5049 4399 5052
rect 4341 5043 4399 5049
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 5362 5083 5420 5089
rect 5362 5049 5374 5083
rect 5408 5080 5420 5083
rect 5626 5080 5632 5092
rect 5408 5052 5632 5080
rect 5408 5049 5420 5052
rect 5362 5043 5420 5049
rect 5626 5040 5632 5052
rect 5684 5040 5690 5092
rect 8386 5080 8392 5092
rect 8347 5052 8392 5080
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 8481 5083 8539 5089
rect 8481 5049 8493 5083
rect 8527 5049 8539 5083
rect 8481 5043 8539 5049
rect 7006 5012 7012 5024
rect 6967 4984 7012 5012
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 8202 5012 8208 5024
rect 8163 4984 8208 5012
rect 8202 4972 8208 4984
rect 8260 5012 8266 5024
rect 8496 5012 8524 5043
rect 8260 4984 8524 5012
rect 8260 4972 8266 4984
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 3697 4811 3755 4817
rect 3697 4777 3709 4811
rect 3743 4808 3755 4811
rect 3970 4808 3976 4820
rect 3743 4780 3976 4808
rect 3743 4777 3755 4780
rect 3697 4771 3755 4777
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 4338 4808 4344 4820
rect 4299 4780 4344 4808
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 5718 4768 5724 4820
rect 5776 4808 5782 4820
rect 5902 4808 5908 4820
rect 5776 4780 5908 4808
rect 5776 4768 5782 4780
rect 5902 4768 5908 4780
rect 5960 4808 5966 4820
rect 6273 4811 6331 4817
rect 6273 4808 6285 4811
rect 5960 4780 6285 4808
rect 5960 4768 5966 4780
rect 6273 4777 6285 4780
rect 6319 4777 6331 4811
rect 8202 4808 8208 4820
rect 8163 4780 8208 4808
rect 6273 4771 6331 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 2866 4700 2872 4752
rect 2924 4740 2930 4752
rect 4798 4740 4804 4752
rect 2924 4712 4804 4740
rect 2924 4700 2930 4712
rect 4798 4700 4804 4712
rect 4856 4700 4862 4752
rect 4890 4700 4896 4752
rect 4948 4740 4954 4752
rect 5030 4743 5088 4749
rect 5030 4740 5042 4743
rect 4948 4712 5042 4740
rect 4948 4700 4954 4712
rect 5030 4709 5042 4712
rect 5076 4709 5088 4743
rect 5030 4703 5088 4709
rect 5442 4700 5448 4752
rect 5500 4740 5506 4752
rect 7098 4740 7104 4752
rect 5500 4712 7104 4740
rect 5500 4700 5506 4712
rect 7098 4700 7104 4712
rect 7156 4700 7162 4752
rect 7466 4700 7472 4752
rect 7524 4740 7530 4752
rect 7650 4749 7656 4752
rect 7606 4743 7656 4749
rect 7606 4740 7618 4743
rect 7524 4712 7618 4740
rect 7524 4700 7530 4712
rect 7606 4709 7618 4712
rect 7652 4709 7656 4743
rect 7606 4703 7656 4709
rect 7650 4700 7656 4703
rect 7708 4700 7714 4752
rect 8386 4700 8392 4752
rect 8444 4740 8450 4752
rect 8573 4743 8631 4749
rect 8573 4740 8585 4743
rect 8444 4712 8585 4740
rect 8444 4700 8450 4712
rect 8573 4709 8585 4712
rect 8619 4740 8631 4743
rect 9815 4743 9873 4749
rect 9815 4740 9827 4743
rect 8619 4712 9827 4740
rect 8619 4709 8631 4712
rect 8573 4703 8631 4709
rect 9815 4709 9827 4712
rect 9861 4709 9873 4743
rect 9815 4703 9873 4709
rect 3028 4675 3086 4681
rect 3028 4641 3040 4675
rect 3074 4672 3086 4675
rect 3510 4672 3516 4684
rect 3074 4644 3516 4672
rect 3074 4641 3086 4644
rect 3028 4635 3086 4641
rect 3510 4632 3516 4644
rect 3568 4632 3574 4684
rect 4706 4604 4712 4616
rect 4667 4576 4712 4604
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 4816 4604 4844 4700
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 5905 4675 5963 4681
rect 5905 4672 5917 4675
rect 5316 4644 5917 4672
rect 5316 4632 5322 4644
rect 5905 4641 5917 4644
rect 5951 4641 5963 4675
rect 7282 4672 7288 4684
rect 7243 4644 7288 4672
rect 5905 4635 5963 4641
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 9728 4675 9786 4681
rect 9728 4641 9740 4675
rect 9774 4672 9786 4675
rect 9950 4672 9956 4684
rect 9774 4644 9956 4672
rect 9774 4641 9786 4644
rect 9728 4635 9786 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10724 4675 10782 4681
rect 10724 4641 10736 4675
rect 10770 4641 10782 4675
rect 10724 4635 10782 4641
rect 10739 4604 10767 4635
rect 10962 4604 10968 4616
rect 4816 4576 10968 4604
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 3970 4496 3976 4548
rect 4028 4536 4034 4548
rect 5629 4539 5687 4545
rect 5629 4536 5641 4539
rect 4028 4508 5641 4536
rect 4028 4496 4034 4508
rect 5629 4505 5641 4508
rect 5675 4505 5687 4539
rect 5629 4499 5687 4505
rect 2682 4428 2688 4480
rect 2740 4468 2746 4480
rect 3099 4471 3157 4477
rect 3099 4468 3111 4471
rect 2740 4440 3111 4468
rect 2740 4428 2746 4440
rect 3099 4437 3111 4440
rect 3145 4437 3157 4471
rect 3099 4431 3157 4437
rect 8846 4428 8852 4480
rect 8904 4468 8910 4480
rect 8941 4471 8999 4477
rect 8941 4468 8953 4471
rect 8904 4440 8953 4468
rect 8904 4428 8910 4440
rect 8941 4437 8953 4440
rect 8987 4468 8999 4471
rect 10827 4471 10885 4477
rect 10827 4468 10839 4471
rect 8987 4440 10839 4468
rect 8987 4437 8999 4440
rect 8941 4431 8999 4437
rect 10827 4437 10839 4440
rect 10873 4437 10885 4471
rect 10827 4431 10885 4437
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 6181 4267 6239 4273
rect 6181 4264 6193 4267
rect 4764 4236 6193 4264
rect 4764 4224 4770 4236
rect 6181 4233 6193 4236
rect 6227 4233 6239 4267
rect 6181 4227 6239 4233
rect 6641 4267 6699 4273
rect 6641 4233 6653 4267
rect 6687 4264 6699 4267
rect 7282 4264 7288 4276
rect 6687 4236 7288 4264
rect 6687 4233 6699 4236
rect 6641 4227 6699 4233
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 8202 4224 8208 4276
rect 8260 4264 8266 4276
rect 8665 4267 8723 4273
rect 8665 4264 8677 4267
rect 8260 4236 8677 4264
rect 8260 4224 8266 4236
rect 8665 4233 8677 4236
rect 8711 4233 8723 4267
rect 9950 4264 9956 4276
rect 9863 4236 9956 4264
rect 8665 4227 8723 4233
rect 2133 4199 2191 4205
rect 2133 4196 2145 4199
rect 2043 4168 2145 4196
rect 2133 4165 2145 4168
rect 2179 4196 2191 4199
rect 3234 4196 3240 4208
rect 2179 4168 3240 4196
rect 2179 4165 2191 4168
rect 2133 4159 2191 4165
rect 1648 4063 1706 4069
rect 1648 4029 1660 4063
rect 1694 4060 1706 4063
rect 2148 4060 2176 4159
rect 3234 4156 3240 4168
rect 3292 4196 3298 4208
rect 4249 4199 4307 4205
rect 4249 4196 4261 4199
rect 3292 4168 4261 4196
rect 3292 4156 3298 4168
rect 4249 4165 4261 4168
rect 4295 4196 4307 4199
rect 5810 4196 5816 4208
rect 4295 4168 5816 4196
rect 4295 4165 4307 4168
rect 4249 4159 4307 4165
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 2731 4131 2789 4137
rect 2731 4097 2743 4131
rect 2777 4128 2789 4131
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 2777 4100 5273 4128
rect 2777 4097 2789 4100
rect 2731 4091 2789 4097
rect 5261 4097 5273 4100
rect 5307 4128 5319 4131
rect 5626 4128 5632 4140
rect 5307 4100 5632 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 7098 4128 7104 4140
rect 7059 4100 7104 4128
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 1694 4032 2176 4060
rect 2644 4063 2702 4069
rect 1694 4029 1706 4032
rect 1648 4023 1706 4029
rect 2644 4029 2656 4063
rect 2690 4060 2702 4063
rect 2866 4060 2872 4072
rect 2690 4032 2872 4060
rect 2690 4029 2702 4032
rect 2644 4023 2702 4029
rect 2866 4020 2872 4032
rect 2924 4060 2930 4072
rect 3053 4063 3111 4069
rect 3053 4060 3065 4063
rect 2924 4032 3065 4060
rect 2924 4020 2930 4032
rect 3053 4029 3065 4032
rect 3099 4029 3111 4063
rect 3053 4023 3111 4029
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4060 4859 4063
rect 4890 4060 4896 4072
rect 4847 4032 4896 4060
rect 4847 4029 4859 4032
rect 4801 4023 4859 4029
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 2501 3995 2559 4001
rect 2501 3961 2513 3995
rect 2547 3992 2559 3995
rect 3697 3995 3755 4001
rect 3697 3992 3709 3995
rect 2547 3964 3709 3992
rect 2547 3961 2559 3964
rect 2501 3955 2559 3961
rect 3697 3961 3709 3964
rect 3743 3961 3755 3995
rect 3697 3955 3755 3961
rect 3789 3995 3847 4001
rect 3789 3961 3801 3995
rect 3835 3992 3847 3995
rect 3970 3992 3976 4004
rect 3835 3964 3976 3992
rect 3835 3961 3847 3964
rect 3789 3955 3847 3961
rect 106 3884 112 3936
rect 164 3924 170 3936
rect 1719 3927 1777 3933
rect 1719 3924 1731 3927
rect 164 3896 1731 3924
rect 164 3884 170 3896
rect 1719 3893 1731 3896
rect 1765 3893 1777 3927
rect 3510 3924 3516 3936
rect 3471 3896 3516 3924
rect 1719 3887 1777 3893
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 3712 3924 3740 3955
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 5350 3992 5356 4004
rect 5263 3964 5356 3992
rect 5350 3952 5356 3964
rect 5408 3992 5414 4004
rect 5718 3992 5724 4004
rect 5408 3964 5724 3992
rect 5408 3952 5414 3964
rect 5718 3952 5724 3964
rect 5776 3952 5782 4004
rect 5905 3995 5963 4001
rect 5905 3961 5917 3995
rect 5951 3961 5963 3995
rect 5905 3955 5963 3961
rect 7463 3995 7521 4001
rect 7463 3961 7475 3995
rect 7509 3992 7521 3995
rect 7650 3992 7656 4004
rect 7509 3964 7656 3992
rect 7509 3961 7521 3964
rect 7463 3955 7521 3961
rect 5920 3924 5948 3955
rect 7650 3952 7656 3964
rect 7708 3952 7714 4004
rect 8680 3992 8708 4227
rect 9950 4224 9956 4236
rect 10008 4264 10014 4276
rect 10321 4267 10379 4273
rect 10321 4264 10333 4267
rect 10008 4236 10333 4264
rect 10008 4224 10014 4236
rect 10321 4233 10333 4236
rect 10367 4264 10379 4267
rect 10870 4264 10876 4276
rect 10367 4236 10876 4264
rect 10367 4233 10379 4236
rect 10321 4227 10379 4233
rect 8846 4156 8852 4208
rect 8904 4196 8910 4208
rect 9766 4196 9772 4208
rect 8904 4168 8984 4196
rect 8904 4156 8910 4168
rect 8956 4137 8984 4168
rect 9232 4168 9772 4196
rect 9232 4140 9260 4168
rect 9766 4156 9772 4168
rect 9824 4156 9830 4208
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 8919 4100 8953 4128
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 9214 4128 9220 4140
rect 9175 4100 9220 4128
rect 8941 4091 8999 4097
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 10428 4069 10456 4236
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 10962 4224 10968 4276
rect 11020 4264 11026 4276
rect 11020 4236 11065 4264
rect 11020 4224 11026 4236
rect 10413 4063 10471 4069
rect 10413 4029 10425 4063
rect 10459 4029 10471 4063
rect 10413 4023 10471 4029
rect 9033 3995 9091 4001
rect 9033 3992 9045 3995
rect 8680 3964 9045 3992
rect 9033 3961 9045 3964
rect 9079 3961 9091 3995
rect 9033 3955 9091 3961
rect 6086 3924 6092 3936
rect 3712 3896 6092 3924
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8202 3924 8208 3936
rect 8067 3896 8208 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 10597 3927 10655 3933
rect 10597 3893 10609 3927
rect 10643 3924 10655 3927
rect 10686 3924 10692 3936
rect 10643 3896 10692 3924
rect 10643 3893 10655 3896
rect 10597 3887 10655 3893
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 3697 3723 3755 3729
rect 3697 3689 3709 3723
rect 3743 3720 3755 3723
rect 3970 3720 3976 3732
rect 3743 3692 3976 3720
rect 3743 3689 3755 3692
rect 3697 3683 3755 3689
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 5350 3720 5356 3732
rect 5311 3692 5356 3720
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 5626 3720 5632 3732
rect 5587 3692 5632 3720
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 7193 3723 7251 3729
rect 7193 3689 7205 3723
rect 7239 3720 7251 3723
rect 7561 3723 7619 3729
rect 7561 3720 7573 3723
rect 7239 3692 7573 3720
rect 7239 3689 7251 3692
rect 7193 3683 7251 3689
rect 7561 3689 7573 3692
rect 7607 3720 7619 3723
rect 7650 3720 7656 3732
rect 7607 3692 7656 3720
rect 7607 3689 7619 3692
rect 7561 3683 7619 3689
rect 7650 3680 7656 3692
rect 7708 3680 7714 3732
rect 7929 3723 7987 3729
rect 7929 3689 7941 3723
rect 7975 3720 7987 3723
rect 8294 3720 8300 3732
rect 7975 3692 8300 3720
rect 7975 3689 7987 3692
rect 7929 3683 7987 3689
rect 8294 3680 8300 3692
rect 8352 3720 8358 3732
rect 10919 3723 10977 3729
rect 10919 3720 10931 3723
rect 8352 3692 10931 3720
rect 8352 3680 8358 3692
rect 10919 3689 10931 3692
rect 10965 3689 10977 3723
rect 10919 3683 10977 3689
rect 1857 3655 1915 3661
rect 1857 3621 1869 3655
rect 1903 3652 1915 3655
rect 2682 3652 2688 3664
rect 1903 3624 2688 3652
rect 1903 3621 1915 3624
rect 1857 3615 1915 3621
rect 2682 3612 2688 3624
rect 2740 3612 2746 3664
rect 4427 3655 4485 3661
rect 4427 3621 4439 3655
rect 4473 3652 4485 3655
rect 4890 3652 4896 3664
rect 4473 3624 4896 3652
rect 4473 3621 4485 3624
rect 4427 3615 4485 3621
rect 4890 3612 4896 3624
rect 4948 3612 4954 3664
rect 5994 3652 6000 3664
rect 5955 3624 6000 3652
rect 5994 3612 6000 3624
rect 6052 3612 6058 3664
rect 6086 3612 6092 3664
rect 6144 3652 6150 3664
rect 6549 3655 6607 3661
rect 6549 3652 6561 3655
rect 6144 3624 6561 3652
rect 6144 3612 6150 3624
rect 6549 3621 6561 3624
rect 6595 3621 6607 3655
rect 8202 3652 8208 3664
rect 8163 3624 8208 3652
rect 6549 3615 6607 3621
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 8757 3655 8815 3661
rect 8757 3621 8769 3655
rect 8803 3652 8815 3655
rect 9214 3652 9220 3664
rect 8803 3624 9220 3652
rect 8803 3621 8815 3624
rect 8757 3615 8815 3621
rect 9214 3612 9220 3624
rect 9272 3612 9278 3664
rect 2016 3587 2074 3593
rect 2016 3553 2028 3587
rect 2062 3584 2074 3587
rect 2590 3584 2596 3596
rect 2062 3556 2596 3584
rect 2062 3553 2074 3556
rect 2016 3547 2074 3553
rect 2590 3544 2596 3556
rect 2648 3544 2654 3596
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 3200 3556 4077 3584
rect 3200 3544 3206 3556
rect 4065 3553 4077 3556
rect 4111 3584 4123 3587
rect 5350 3584 5356 3596
rect 4111 3556 5356 3584
rect 4111 3553 4123 3556
rect 4065 3547 4123 3553
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 9674 3584 9680 3596
rect 9587 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3584 9738 3596
rect 10226 3584 10232 3596
rect 9732 3556 10232 3584
rect 9732 3544 9738 3556
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 10816 3587 10874 3593
rect 10816 3553 10828 3587
rect 10862 3553 10874 3587
rect 10816 3547 10874 3553
rect 2498 3476 2504 3528
rect 2556 3516 2562 3528
rect 2961 3519 3019 3525
rect 2961 3516 2973 3519
rect 2556 3488 2973 3516
rect 2556 3476 2562 3488
rect 2961 3485 2973 3488
rect 3007 3485 3019 3519
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 2961 3479 3019 3485
rect 4126 3488 5917 3516
rect 2087 3451 2145 3457
rect 2087 3417 2099 3451
rect 2133 3448 2145 3451
rect 4126 3448 4154 3488
rect 5905 3485 5917 3488
rect 5951 3516 5963 3519
rect 6178 3516 6184 3528
rect 5951 3488 6184 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 9398 3516 9404 3528
rect 8159 3488 9404 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 2133 3420 4154 3448
rect 2133 3417 2145 3420
rect 2087 3411 2145 3417
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 10831 3448 10859 3547
rect 11238 3448 11244 3460
rect 6972 3420 11244 3448
rect 6972 3408 6978 3420
rect 11238 3408 11244 3420
rect 11296 3448 11302 3460
rect 11606 3448 11612 3460
rect 11296 3420 11612 3448
rect 11296 3408 11302 3420
rect 11606 3408 11612 3420
rect 11664 3408 11670 3460
rect 2685 3383 2743 3389
rect 2685 3349 2697 3383
rect 2731 3380 2743 3383
rect 2774 3380 2780 3392
rect 2731 3352 2780 3380
rect 2731 3349 2743 3352
rect 2685 3343 2743 3349
rect 2774 3340 2780 3352
rect 2832 3340 2838 3392
rect 3510 3340 3516 3392
rect 3568 3380 3574 3392
rect 4985 3383 5043 3389
rect 4985 3380 4997 3383
rect 3568 3352 4997 3380
rect 3568 3340 3574 3352
rect 4985 3349 4997 3352
rect 5031 3349 5043 3383
rect 4985 3343 5043 3349
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 9861 3383 9919 3389
rect 9861 3380 9873 3383
rect 9364 3352 9873 3380
rect 9364 3340 9370 3352
rect 9861 3349 9873 3352
rect 9907 3349 9919 3383
rect 9861 3343 9919 3349
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 1118 3136 1124 3188
rect 1176 3176 1182 3188
rect 1489 3179 1547 3185
rect 1489 3176 1501 3179
rect 1176 3148 1501 3176
rect 1176 3136 1182 3148
rect 1489 3145 1501 3148
rect 1535 3176 1547 3179
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 1535 3148 2145 3176
rect 1535 3145 1547 3148
rect 1489 3139 1547 3145
rect 2133 3145 2145 3148
rect 2179 3176 2191 3179
rect 2406 3176 2412 3188
rect 2179 3148 2412 3176
rect 2179 3145 2191 3148
rect 2133 3139 2191 3145
rect 2406 3136 2412 3148
rect 2464 3136 2470 3188
rect 2501 3179 2559 3185
rect 2501 3145 2513 3179
rect 2547 3176 2559 3179
rect 2590 3176 2596 3188
rect 2547 3148 2596 3176
rect 2547 3145 2559 3148
rect 2501 3139 2559 3145
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 2958 3136 2964 3188
rect 3016 3176 3022 3188
rect 5350 3176 5356 3188
rect 3016 3148 5212 3176
rect 5311 3148 5356 3176
rect 3016 3136 3022 3148
rect 1719 3111 1777 3117
rect 1719 3077 1731 3111
rect 1765 3108 1777 3111
rect 4982 3108 4988 3120
rect 1765 3080 4988 3108
rect 1765 3077 1777 3080
rect 1719 3071 1777 3077
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 2682 3040 2688 3052
rect 2643 3012 2688 3040
rect 2682 3000 2688 3012
rect 2740 3000 2746 3052
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4212 3012 4257 3040
rect 4212 3000 4218 3012
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2972 3387 2975
rect 5184 2972 5212 3148
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 5905 3179 5963 3185
rect 5905 3145 5917 3179
rect 5951 3176 5963 3179
rect 5994 3176 6000 3188
rect 5951 3148 6000 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6178 3176 6184 3188
rect 6139 3148 6184 3176
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 8021 3179 8079 3185
rect 8021 3145 8033 3179
rect 8067 3176 8079 3179
rect 8202 3176 8208 3188
rect 8067 3148 8208 3176
rect 8067 3145 8079 3148
rect 8021 3139 8079 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9217 3179 9275 3185
rect 9217 3145 9229 3179
rect 9263 3176 9275 3179
rect 9398 3176 9404 3188
rect 9263 3148 9404 3176
rect 9263 3145 9275 3148
rect 9217 3139 9275 3145
rect 9398 3136 9404 3148
rect 9456 3136 9462 3188
rect 9585 3179 9643 3185
rect 9585 3145 9597 3179
rect 9631 3176 9643 3179
rect 9674 3176 9680 3188
rect 9631 3148 9680 3176
rect 9631 3145 9643 3148
rect 9585 3139 9643 3145
rect 9674 3136 9680 3148
rect 9732 3176 9738 3188
rect 10042 3176 10048 3188
rect 9732 3148 10048 3176
rect 9732 3136 9738 3148
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 10226 3176 10232 3188
rect 10187 3148 10232 3176
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 11606 3176 11612 3188
rect 11567 3148 11612 3176
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 5534 3068 5540 3120
rect 5592 3108 5598 3120
rect 8754 3108 8760 3120
rect 5592 3080 8524 3108
rect 8715 3080 8760 3108
rect 5592 3068 5598 3080
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3040 8263 3043
rect 8294 3040 8300 3052
rect 8251 3012 8300 3040
rect 8251 3009 8263 3012
rect 8205 3003 8263 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8496 3040 8524 3080
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 9646 3080 10640 3108
rect 9646 3040 9674 3080
rect 8496 3012 9674 3040
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 3375 2944 5120 2972
rect 5184 2944 6837 2972
rect 3375 2941 3387 2944
rect 3329 2935 3387 2941
rect 2774 2904 2780 2916
rect 2735 2876 2780 2904
rect 2774 2864 2780 2876
rect 2832 2864 2838 2916
rect 4519 2907 4577 2913
rect 4519 2873 4531 2907
rect 4565 2904 4577 2907
rect 4890 2904 4896 2916
rect 4565 2876 4896 2904
rect 4565 2873 4577 2876
rect 4519 2867 4577 2873
rect 3697 2839 3755 2845
rect 3697 2805 3709 2839
rect 3743 2836 3755 2839
rect 3973 2839 4031 2845
rect 3973 2836 3985 2839
rect 3743 2808 3985 2836
rect 3743 2805 3755 2808
rect 3697 2799 3755 2805
rect 3973 2805 3985 2808
rect 4019 2836 4031 2839
rect 4534 2836 4562 2867
rect 4890 2864 4896 2876
rect 4948 2864 4954 2916
rect 5092 2904 5120 2944
rect 6825 2941 6837 2944
rect 6871 2972 6883 2975
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 6871 2944 7389 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 7377 2941 7389 2944
rect 7423 2941 7435 2975
rect 7377 2935 7435 2941
rect 9674 2932 9680 2984
rect 9732 2972 9738 2984
rect 10612 2972 10640 3080
rect 10816 2975 10874 2981
rect 10816 2972 10828 2975
rect 9732 2944 9777 2972
rect 10612 2944 10828 2972
rect 9732 2932 9738 2944
rect 10816 2941 10828 2944
rect 10862 2972 10874 2975
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 10862 2944 11253 2972
rect 10862 2941 10874 2944
rect 10816 2935 10874 2941
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 11241 2935 11299 2941
rect 5902 2904 5908 2916
rect 5092 2876 5908 2904
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 12526 2904 12532 2916
rect 8352 2876 8397 2904
rect 8496 2876 12532 2904
rect 8352 2864 8358 2876
rect 5074 2836 5080 2848
rect 4019 2808 4562 2836
rect 5035 2808 5080 2836
rect 4019 2805 4031 2808
rect 3973 2799 4031 2805
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 7009 2839 7067 2845
rect 7009 2805 7021 2839
rect 7055 2836 7067 2839
rect 8496 2836 8524 2876
rect 12526 2864 12532 2876
rect 12584 2864 12590 2916
rect 9858 2836 9864 2848
rect 7055 2808 8524 2836
rect 9819 2808 9864 2836
rect 7055 2805 7067 2808
rect 7009 2799 7067 2805
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 10410 2796 10416 2848
rect 10468 2836 10474 2848
rect 10919 2839 10977 2845
rect 10919 2836 10931 2839
rect 10468 2808 10931 2836
rect 10468 2796 10474 2808
rect 10919 2805 10931 2808
rect 10965 2805 10977 2839
rect 10919 2799 10977 2805
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 3510 2632 3516 2644
rect 2608 2604 3516 2632
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 2498 2564 2504 2576
rect 2363 2536 2504 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 2498 2524 2504 2536
rect 2556 2524 2562 2576
rect 2608 2573 2636 2604
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4249 2635 4307 2641
rect 4249 2632 4261 2635
rect 4212 2604 4261 2632
rect 4212 2592 4218 2604
rect 4249 2601 4261 2604
rect 4295 2601 4307 2635
rect 4249 2595 4307 2601
rect 5994 2592 6000 2644
rect 6052 2632 6058 2644
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 6052 2604 6653 2632
rect 6052 2592 6058 2604
rect 6641 2601 6653 2604
rect 6687 2601 6699 2635
rect 6641 2595 6699 2601
rect 8113 2635 8171 2641
rect 8113 2601 8125 2635
rect 8159 2632 8171 2635
rect 8202 2632 8208 2644
rect 8159 2604 8208 2632
rect 8159 2601 8171 2604
rect 8113 2595 8171 2601
rect 2593 2567 2651 2573
rect 2593 2533 2605 2567
rect 2639 2533 2651 2567
rect 2593 2527 2651 2533
rect 3145 2567 3203 2573
rect 3145 2533 3157 2567
rect 3191 2564 3203 2567
rect 3234 2564 3240 2576
rect 3191 2536 3240 2564
rect 3191 2533 3203 2536
rect 3145 2527 3203 2533
rect 3234 2524 3240 2536
rect 3292 2524 3298 2576
rect 4801 2567 4859 2573
rect 4801 2564 4813 2567
rect 4126 2536 4813 2564
rect 1464 2499 1522 2505
rect 1464 2465 1476 2499
rect 1510 2496 1522 2499
rect 1510 2468 1992 2496
rect 1510 2465 1522 2468
rect 1464 2459 1522 2465
rect 1964 2369 1992 2468
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 4126 2428 4154 2536
rect 4801 2533 4813 2536
rect 4847 2564 4859 2567
rect 5074 2564 5080 2576
rect 4847 2536 5080 2564
rect 4847 2533 4859 2536
rect 4801 2527 4859 2533
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 5629 2567 5687 2573
rect 5629 2533 5641 2567
rect 5675 2564 5687 2567
rect 6086 2564 6092 2576
rect 5675 2536 6092 2564
rect 5675 2533 5687 2536
rect 5629 2527 5687 2533
rect 6086 2524 6092 2536
rect 6144 2524 6150 2576
rect 6656 2564 6684 2595
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 11609 2635 11667 2641
rect 11609 2601 11621 2635
rect 11655 2632 11667 2635
rect 15562 2632 15568 2644
rect 11655 2604 15568 2632
rect 11655 2601 11667 2604
rect 11609 2595 11667 2601
rect 15562 2592 15568 2604
rect 15620 2592 15626 2644
rect 7101 2567 7159 2573
rect 7101 2564 7113 2567
rect 6656 2536 7113 2564
rect 7101 2533 7113 2536
rect 7147 2533 7159 2567
rect 7101 2527 7159 2533
rect 8662 2524 8668 2576
rect 8720 2564 8726 2576
rect 10873 2567 10931 2573
rect 10873 2564 10885 2567
rect 8720 2536 10885 2564
rect 8720 2524 8726 2536
rect 7926 2456 7932 2508
rect 7984 2496 7990 2508
rect 10336 2505 10364 2536
rect 10873 2533 10885 2536
rect 10919 2533 10931 2567
rect 10873 2527 10931 2533
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 7984 2468 8493 2496
rect 7984 2456 7990 2468
rect 8481 2465 8493 2468
rect 8527 2496 8539 2499
rect 9033 2499 9091 2505
rect 9033 2496 9045 2499
rect 8527 2468 9045 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 9033 2465 9045 2468
rect 9079 2465 9091 2499
rect 9033 2459 9091 2465
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2465 10379 2499
rect 11422 2496 11428 2508
rect 11383 2468 11428 2496
rect 10321 2459 10379 2465
rect 11422 2456 11428 2468
rect 11480 2496 11486 2508
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11480 2468 11989 2496
rect 11480 2456 11486 2468
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 13170 2496 13176 2508
rect 13131 2468 13176 2496
rect 11977 2459 12035 2465
rect 13170 2456 13176 2468
rect 13228 2496 13234 2508
rect 13725 2499 13783 2505
rect 13725 2496 13737 2499
rect 13228 2468 13737 2496
rect 13228 2456 13234 2468
rect 13725 2465 13737 2468
rect 13771 2465 13783 2499
rect 13725 2459 13783 2465
rect 4982 2428 4988 2440
rect 2832 2400 4154 2428
rect 4943 2400 4988 2428
rect 2832 2388 2838 2400
rect 4982 2388 4988 2400
rect 5040 2428 5046 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5040 2400 5917 2428
rect 5040 2388 5046 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2428 6423 2431
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 6411 2400 7021 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 7009 2397 7021 2400
rect 7055 2428 7067 2431
rect 10410 2428 10416 2440
rect 7055 2400 10416 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 1949 2363 2007 2369
rect 1949 2329 1961 2363
rect 1995 2360 2007 2363
rect 6730 2360 6736 2372
rect 1995 2332 6736 2360
rect 1995 2329 2007 2332
rect 1949 2323 2007 2329
rect 6730 2320 6736 2332
rect 6788 2320 6794 2372
rect 7561 2363 7619 2369
rect 7561 2360 7573 2363
rect 6840 2332 7573 2360
rect 1535 2295 1593 2301
rect 1535 2261 1547 2295
rect 1581 2292 1593 2295
rect 3326 2292 3332 2304
rect 1581 2264 3332 2292
rect 1581 2261 1593 2264
rect 1535 2255 1593 2261
rect 3326 2252 3332 2264
rect 3384 2252 3390 2304
rect 5902 2252 5908 2304
rect 5960 2292 5966 2304
rect 6840 2292 6868 2332
rect 7561 2329 7573 2332
rect 7607 2329 7619 2363
rect 7561 2323 7619 2329
rect 10505 2363 10563 2369
rect 10505 2329 10517 2363
rect 10551 2360 10563 2363
rect 11698 2360 11704 2372
rect 10551 2332 11704 2360
rect 10551 2329 10563 2332
rect 10505 2323 10563 2329
rect 11698 2320 11704 2332
rect 11756 2320 11762 2372
rect 13357 2363 13415 2369
rect 13357 2329 13369 2363
rect 13403 2360 13415 2363
rect 14642 2360 14648 2372
rect 13403 2332 14648 2360
rect 13403 2329 13415 2332
rect 13357 2323 13415 2329
rect 14642 2320 14648 2332
rect 14700 2320 14706 2372
rect 5960 2264 6868 2292
rect 5960 2252 5966 2264
rect 8294 2252 8300 2304
rect 8352 2292 8358 2304
rect 8665 2295 8723 2301
rect 8665 2292 8677 2295
rect 8352 2264 8677 2292
rect 8352 2252 8358 2264
rect 8665 2261 8677 2264
rect 8711 2261 8723 2295
rect 8665 2255 8723 2261
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 3418 76 3424 128
rect 3476 116 3482 128
rect 4798 116 4804 128
rect 3476 88 4804 116
rect 3476 76 3482 88
rect 4798 76 4804 88
rect 4856 76 4862 128
rect 7006 76 7012 128
rect 7064 116 7070 128
rect 13722 116 13728 128
rect 7064 88 13728 116
rect 7064 76 7070 88
rect 13722 76 13728 88
rect 13780 76 13786 128
<< via1 >>
rect 1216 39652 1268 39704
rect 3240 39652 3292 39704
rect 1400 39584 1452 39636
rect 2136 39584 2188 39636
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 12440 36660 12492 36712
rect 9956 36524 10008 36576
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 8852 36320 8904 36372
rect 2964 36252 3016 36304
rect 7564 36227 7616 36236
rect 7564 36193 7582 36227
rect 7582 36193 7616 36227
rect 7564 36184 7616 36193
rect 7840 36184 7892 36236
rect 8392 36184 8444 36236
rect 9680 36227 9732 36236
rect 9680 36193 9724 36227
rect 9724 36193 9732 36227
rect 9680 36184 9732 36193
rect 8116 35980 8168 36032
rect 8208 36023 8260 36032
rect 8208 35989 8217 36023
rect 8217 35989 8251 36023
rect 8251 35989 8260 36023
rect 8208 35980 8260 35989
rect 10324 35980 10376 36032
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 13452 35776 13504 35828
rect 7840 35751 7892 35760
rect 7840 35717 7849 35751
rect 7849 35717 7883 35751
rect 7883 35717 7892 35751
rect 7840 35708 7892 35717
rect 11244 35708 11296 35760
rect 8116 35640 8168 35692
rect 8392 35640 8444 35692
rect 9680 35683 9732 35692
rect 9680 35649 9689 35683
rect 9689 35649 9723 35683
rect 9723 35649 9732 35683
rect 9680 35640 9732 35649
rect 10324 35683 10376 35692
rect 10324 35649 10333 35683
rect 10333 35649 10367 35683
rect 10367 35649 10376 35683
rect 10324 35640 10376 35649
rect 4436 35572 4488 35624
rect 8208 35436 8260 35488
rect 8484 35504 8536 35556
rect 10416 35547 10468 35556
rect 10416 35513 10425 35547
rect 10425 35513 10459 35547
rect 10459 35513 10468 35547
rect 10416 35504 10468 35513
rect 10968 35547 11020 35556
rect 10968 35513 10977 35547
rect 10977 35513 11011 35547
rect 11011 35513 11020 35547
rect 10968 35504 11020 35513
rect 9680 35436 9732 35488
rect 10876 35436 10928 35488
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 8024 35232 8076 35284
rect 8116 35232 8168 35284
rect 9956 35232 10008 35284
rect 14648 35232 14700 35284
rect 5816 35164 5868 35216
rect 8208 35207 8260 35216
rect 8208 35173 8217 35207
rect 8217 35173 8251 35207
rect 8251 35173 8260 35207
rect 8208 35164 8260 35173
rect 10600 35207 10652 35216
rect 10600 35173 10609 35207
rect 10609 35173 10643 35207
rect 10643 35173 10652 35207
rect 10600 35164 10652 35173
rect 6736 35096 6788 35148
rect 7012 35096 7064 35148
rect 12164 35096 12216 35148
rect 12992 35139 13044 35148
rect 12992 35105 13001 35139
rect 13001 35105 13035 35139
rect 13035 35105 13044 35139
rect 12992 35096 13044 35105
rect 8116 35071 8168 35080
rect 8116 35037 8125 35071
rect 8125 35037 8159 35071
rect 8159 35037 8168 35071
rect 8116 35028 8168 35037
rect 8300 35028 8352 35080
rect 10508 35071 10560 35080
rect 10508 35037 10517 35071
rect 10517 35037 10551 35071
rect 10551 35037 10560 35071
rect 10508 35028 10560 35037
rect 11428 35028 11480 35080
rect 5816 34960 5868 35012
rect 12624 34960 12676 35012
rect 7656 34935 7708 34944
rect 7656 34901 7665 34935
rect 7665 34901 7699 34935
rect 7699 34901 7708 34935
rect 7656 34892 7708 34901
rect 12532 34892 12584 34944
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 5816 34731 5868 34740
rect 5816 34697 5825 34731
rect 5825 34697 5859 34731
rect 5859 34697 5868 34731
rect 5816 34688 5868 34697
rect 9772 34688 9824 34740
rect 11336 34688 11388 34740
rect 7748 34620 7800 34672
rect 8300 34595 8352 34604
rect 8300 34561 8309 34595
rect 8309 34561 8343 34595
rect 8343 34561 8352 34595
rect 8300 34552 8352 34561
rect 4160 34484 4212 34536
rect 12164 34620 12216 34672
rect 9956 34552 10008 34604
rect 10968 34595 11020 34604
rect 10968 34561 10977 34595
rect 10977 34561 11011 34595
rect 11011 34561 11020 34595
rect 10968 34552 11020 34561
rect 12440 34527 12492 34536
rect 12440 34493 12449 34527
rect 12449 34493 12483 34527
rect 12483 34493 12492 34527
rect 12440 34484 12492 34493
rect 12992 34484 13044 34536
rect 6092 34416 6144 34468
rect 7656 34459 7708 34468
rect 7656 34425 7665 34459
rect 7665 34425 7699 34459
rect 7699 34425 7708 34459
rect 7656 34416 7708 34425
rect 6736 34348 6788 34400
rect 7012 34391 7064 34400
rect 7012 34357 7021 34391
rect 7021 34357 7055 34391
rect 7055 34357 7064 34391
rect 7012 34348 7064 34357
rect 7932 34416 7984 34468
rect 8116 34416 8168 34468
rect 8208 34348 8260 34400
rect 9496 34348 9548 34400
rect 10232 34348 10284 34400
rect 10692 34416 10744 34468
rect 10600 34348 10652 34400
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 8116 34144 8168 34196
rect 9956 34144 10008 34196
rect 15568 34144 15620 34196
rect 6368 34119 6420 34128
rect 6368 34085 6377 34119
rect 6377 34085 6411 34119
rect 6411 34085 6420 34119
rect 6368 34076 6420 34085
rect 7932 34119 7984 34128
rect 7932 34085 7941 34119
rect 7941 34085 7975 34119
rect 7975 34085 7984 34119
rect 7932 34076 7984 34085
rect 8484 34119 8536 34128
rect 8484 34085 8493 34119
rect 8493 34085 8527 34119
rect 8527 34085 8536 34119
rect 8484 34076 8536 34085
rect 5264 34008 5316 34060
rect 10968 34076 11020 34128
rect 12164 34008 12216 34060
rect 12440 34008 12492 34060
rect 13452 34008 13504 34060
rect 7840 33983 7892 33992
rect 7840 33949 7849 33983
rect 7849 33949 7883 33983
rect 7883 33949 7892 33983
rect 7840 33940 7892 33949
rect 9772 33940 9824 33992
rect 11336 33940 11388 33992
rect 6184 33872 6236 33924
rect 8484 33872 8536 33924
rect 11060 33872 11112 33924
rect 7564 33847 7616 33856
rect 7564 33813 7573 33847
rect 7573 33813 7607 33847
rect 7607 33813 7616 33847
rect 7564 33804 7616 33813
rect 10508 33804 10560 33856
rect 12164 33804 12216 33856
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 6092 33600 6144 33652
rect 6368 33600 6420 33652
rect 10232 33643 10284 33652
rect 10232 33609 10241 33643
rect 10241 33609 10275 33643
rect 10275 33609 10284 33643
rect 10232 33600 10284 33609
rect 10968 33643 11020 33652
rect 10968 33609 10977 33643
rect 10977 33609 11011 33643
rect 11011 33609 11020 33643
rect 10968 33600 11020 33609
rect 11520 33600 11572 33652
rect 13452 33643 13504 33652
rect 13452 33609 13461 33643
rect 13461 33609 13495 33643
rect 13495 33609 13504 33643
rect 13452 33600 13504 33609
rect 10416 33532 10468 33584
rect 7564 33507 7616 33516
rect 7564 33473 7573 33507
rect 7573 33473 7607 33507
rect 7607 33473 7616 33507
rect 7564 33464 7616 33473
rect 8024 33464 8076 33516
rect 8300 33464 8352 33516
rect 9772 33464 9824 33516
rect 664 33396 716 33448
rect 5264 33303 5316 33312
rect 5264 33269 5273 33303
rect 5273 33269 5307 33303
rect 5307 33269 5316 33303
rect 5264 33260 5316 33269
rect 9312 33439 9364 33448
rect 6000 33260 6052 33312
rect 9312 33405 9321 33439
rect 9321 33405 9355 33439
rect 9355 33405 9364 33439
rect 9312 33396 9364 33405
rect 12532 33507 12584 33516
rect 12532 33473 12541 33507
rect 12541 33473 12575 33507
rect 12575 33473 12584 33507
rect 12532 33464 12584 33473
rect 12808 33507 12860 33516
rect 12808 33473 12817 33507
rect 12817 33473 12851 33507
rect 12851 33473 12860 33507
rect 12808 33464 12860 33473
rect 7656 33371 7708 33380
rect 7656 33337 7665 33371
rect 7665 33337 7699 33371
rect 7699 33337 7708 33371
rect 7656 33328 7708 33337
rect 9956 33328 10008 33380
rect 10784 33328 10836 33380
rect 12256 33328 12308 33380
rect 7012 33260 7064 33312
rect 8208 33260 8260 33312
rect 9588 33260 9640 33312
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 6184 33099 6236 33108
rect 6184 33065 6193 33099
rect 6193 33065 6227 33099
rect 6227 33065 6236 33099
rect 6184 33056 6236 33065
rect 7104 33099 7156 33108
rect 7104 33065 7113 33099
rect 7113 33065 7147 33099
rect 7147 33065 7156 33099
rect 7104 33056 7156 33065
rect 7656 33099 7708 33108
rect 7656 33065 7665 33099
rect 7665 33065 7699 33099
rect 7699 33065 7708 33099
rect 7656 33056 7708 33065
rect 7932 33099 7984 33108
rect 7932 33065 7941 33099
rect 7941 33065 7975 33099
rect 7975 33065 7984 33099
rect 7932 33056 7984 33065
rect 9956 33056 10008 33108
rect 10416 33056 10468 33108
rect 11520 33056 11572 33108
rect 12532 33099 12584 33108
rect 7840 32988 7892 33040
rect 10968 32988 11020 33040
rect 11704 32988 11756 33040
rect 12532 33065 12541 33099
rect 12541 33065 12575 33099
rect 12575 33065 12584 33099
rect 12532 33056 12584 33065
rect 12808 32988 12860 33040
rect 4068 32920 4120 32972
rect 5724 32963 5776 32972
rect 5724 32929 5768 32963
rect 5768 32929 5776 32963
rect 5724 32920 5776 32929
rect 12992 32963 13044 32972
rect 7380 32852 7432 32904
rect 8300 32852 8352 32904
rect 10416 32852 10468 32904
rect 5264 32784 5316 32836
rect 10784 32784 10836 32836
rect 12992 32929 13001 32963
rect 13001 32929 13035 32963
rect 13035 32929 13044 32963
rect 12992 32920 13044 32929
rect 11520 32895 11572 32904
rect 11520 32861 11529 32895
rect 11529 32861 11563 32895
rect 11563 32861 11572 32895
rect 11520 32852 11572 32861
rect 12440 32784 12492 32836
rect 8760 32716 8812 32768
rect 9312 32759 9364 32768
rect 9312 32725 9321 32759
rect 9321 32725 9355 32759
rect 9355 32725 9364 32759
rect 9312 32716 9364 32725
rect 11336 32759 11388 32768
rect 11336 32725 11345 32759
rect 11345 32725 11379 32759
rect 11379 32725 11388 32759
rect 11336 32716 11388 32725
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 5724 32555 5776 32564
rect 5724 32521 5733 32555
rect 5733 32521 5767 32555
rect 5767 32521 5776 32555
rect 5724 32512 5776 32521
rect 7472 32512 7524 32564
rect 7932 32512 7984 32564
rect 8300 32512 8352 32564
rect 9496 32555 9548 32564
rect 9496 32521 9505 32555
rect 9505 32521 9539 32555
rect 9539 32521 9548 32555
rect 9496 32512 9548 32521
rect 11704 32555 11756 32564
rect 11704 32521 11713 32555
rect 11713 32521 11747 32555
rect 11747 32521 11756 32555
rect 11704 32512 11756 32521
rect 12164 32512 12216 32564
rect 6828 32444 6880 32496
rect 7840 32444 7892 32496
rect 7104 32376 7156 32428
rect 6828 32351 6880 32360
rect 6828 32317 6837 32351
rect 6837 32317 6871 32351
rect 6871 32317 6880 32351
rect 6828 32308 6880 32317
rect 8760 32376 8812 32428
rect 10324 32351 10376 32360
rect 10324 32317 10333 32351
rect 10333 32317 10367 32351
rect 10367 32317 10376 32351
rect 10324 32308 10376 32317
rect 10232 32283 10284 32292
rect 7288 32172 7340 32224
rect 10232 32249 10241 32283
rect 10241 32249 10275 32283
rect 10275 32249 10284 32283
rect 10232 32240 10284 32249
rect 9588 32172 9640 32224
rect 10416 32215 10468 32224
rect 10416 32181 10425 32215
rect 10425 32181 10459 32215
rect 10459 32181 10468 32215
rect 10416 32172 10468 32181
rect 12348 32172 12400 32224
rect 12992 32215 13044 32224
rect 12992 32181 13001 32215
rect 13001 32181 13035 32215
rect 13035 32181 13044 32215
rect 12992 32172 13044 32181
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 9772 32011 9824 32020
rect 9772 31977 9781 32011
rect 9781 31977 9815 32011
rect 9815 31977 9824 32011
rect 9772 31968 9824 31977
rect 11520 31968 11572 32020
rect 6828 31943 6880 31952
rect 6828 31909 6837 31943
rect 6837 31909 6871 31943
rect 6871 31909 6880 31943
rect 6828 31900 6880 31909
rect 5540 31832 5592 31884
rect 6644 31875 6696 31884
rect 6644 31841 6653 31875
rect 6653 31841 6687 31875
rect 6687 31841 6696 31875
rect 6644 31832 6696 31841
rect 7656 31832 7708 31884
rect 8116 31875 8168 31884
rect 8116 31841 8125 31875
rect 8125 31841 8159 31875
rect 8159 31841 8168 31875
rect 8116 31832 8168 31841
rect 8760 31900 8812 31952
rect 9956 31875 10008 31884
rect 9956 31841 9965 31875
rect 9965 31841 9999 31875
rect 9999 31841 10008 31875
rect 9956 31832 10008 31841
rect 10232 31875 10284 31884
rect 10232 31841 10241 31875
rect 10241 31841 10275 31875
rect 10275 31841 10284 31875
rect 10232 31832 10284 31841
rect 11244 31875 11296 31884
rect 11244 31841 11253 31875
rect 11253 31841 11287 31875
rect 11287 31841 11296 31875
rect 11244 31832 11296 31841
rect 11520 31832 11572 31884
rect 15476 31832 15528 31884
rect 10324 31696 10376 31748
rect 7380 31628 7432 31680
rect 8668 31671 8720 31680
rect 8668 31637 8677 31671
rect 8677 31637 8711 31671
rect 8711 31637 8720 31671
rect 8668 31628 8720 31637
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 7380 31331 7432 31340
rect 7380 31297 7389 31331
rect 7389 31297 7423 31331
rect 7423 31297 7432 31331
rect 7380 31288 7432 31297
rect 6920 31263 6972 31272
rect 6920 31229 6929 31263
rect 6929 31229 6963 31263
rect 6963 31229 6972 31263
rect 6920 31220 6972 31229
rect 9312 31331 9364 31340
rect 9312 31297 9321 31331
rect 9321 31297 9355 31331
rect 9355 31297 9364 31331
rect 9312 31288 9364 31297
rect 8668 31263 8720 31272
rect 5540 31084 5592 31136
rect 6644 31127 6696 31136
rect 6644 31093 6653 31127
rect 6653 31093 6687 31127
rect 6687 31093 6696 31127
rect 8668 31229 8677 31263
rect 8677 31229 8711 31263
rect 8711 31229 8720 31263
rect 8668 31220 8720 31229
rect 10232 31424 10284 31476
rect 9956 31356 10008 31408
rect 12072 31356 12124 31408
rect 11060 31288 11112 31340
rect 6644 31084 6696 31093
rect 8116 31084 8168 31136
rect 8668 31084 8720 31136
rect 10968 31152 11020 31204
rect 12164 31152 12216 31204
rect 11244 31084 11296 31136
rect 12440 31084 12492 31136
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 7656 30923 7708 30932
rect 7656 30889 7665 30923
rect 7665 30889 7699 30923
rect 7699 30889 7708 30923
rect 7656 30880 7708 30889
rect 8024 30880 8076 30932
rect 8576 30880 8628 30932
rect 8300 30812 8352 30864
rect 6736 30744 6788 30796
rect 5264 30676 5316 30728
rect 7104 30676 7156 30728
rect 11060 30880 11112 30932
rect 9312 30812 9364 30864
rect 11428 30855 11480 30864
rect 11428 30821 11437 30855
rect 11437 30821 11471 30855
rect 11471 30821 11480 30855
rect 11428 30812 11480 30821
rect 11336 30719 11388 30728
rect 11336 30685 11345 30719
rect 11345 30685 11379 30719
rect 11379 30685 11388 30719
rect 11336 30676 11388 30685
rect 12164 30676 12216 30728
rect 6920 30583 6972 30592
rect 6920 30549 6929 30583
rect 6929 30549 6963 30583
rect 6963 30549 6972 30583
rect 6920 30540 6972 30549
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 8484 30336 8536 30388
rect 11428 30336 11480 30388
rect 7472 30175 7524 30184
rect 7472 30141 7481 30175
rect 7481 30141 7515 30175
rect 7515 30141 7524 30175
rect 7472 30132 7524 30141
rect 12164 30268 12216 30320
rect 11336 30200 11388 30252
rect 9956 30132 10008 30184
rect 6644 29996 6696 30048
rect 7564 30039 7616 30048
rect 7564 30005 7573 30039
rect 7573 30005 7607 30039
rect 7607 30005 7616 30039
rect 7564 29996 7616 30005
rect 8300 30039 8352 30048
rect 8300 30005 8309 30039
rect 8309 30005 8343 30039
rect 8343 30005 8352 30039
rect 8300 29996 8352 30005
rect 9312 30039 9364 30048
rect 9312 30005 9321 30039
rect 9321 30005 9355 30039
rect 9355 30005 9364 30039
rect 9312 29996 9364 30005
rect 10232 30039 10284 30048
rect 10232 30005 10241 30039
rect 10241 30005 10275 30039
rect 10275 30005 10284 30039
rect 10232 29996 10284 30005
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 7472 29835 7524 29844
rect 7472 29801 7481 29835
rect 7481 29801 7515 29835
rect 7515 29801 7524 29835
rect 7472 29792 7524 29801
rect 8024 29792 8076 29844
rect 10968 29835 11020 29844
rect 10968 29801 10977 29835
rect 10977 29801 11011 29835
rect 11011 29801 11020 29835
rect 10968 29792 11020 29801
rect 10232 29724 10284 29776
rect 11980 29767 12032 29776
rect 11980 29733 11989 29767
rect 11989 29733 12023 29767
rect 12023 29733 12032 29767
rect 11980 29724 12032 29733
rect 6644 29656 6696 29708
rect 8024 29699 8076 29708
rect 8024 29665 8033 29699
rect 8033 29665 8067 29699
rect 8067 29665 8076 29699
rect 8024 29656 8076 29665
rect 8668 29656 8720 29708
rect 6736 29588 6788 29640
rect 7196 29631 7248 29640
rect 7196 29597 7205 29631
rect 7205 29597 7239 29631
rect 7239 29597 7248 29631
rect 7196 29588 7248 29597
rect 8852 29588 8904 29640
rect 10600 29588 10652 29640
rect 11888 29631 11940 29640
rect 11888 29597 11897 29631
rect 11897 29597 11931 29631
rect 11931 29597 11940 29631
rect 11888 29588 11940 29597
rect 12164 29631 12216 29640
rect 12164 29597 12173 29631
rect 12173 29597 12207 29631
rect 12207 29597 12216 29631
rect 12164 29588 12216 29597
rect 5632 29452 5684 29504
rect 9956 29495 10008 29504
rect 9956 29461 9965 29495
rect 9965 29461 9999 29495
rect 9999 29461 10008 29495
rect 9956 29452 10008 29461
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 5080 29248 5132 29300
rect 5908 29248 5960 29300
rect 8116 29248 8168 29300
rect 8300 29291 8352 29300
rect 8300 29257 8309 29291
rect 8309 29257 8343 29291
rect 8343 29257 8352 29291
rect 8300 29248 8352 29257
rect 8668 29291 8720 29300
rect 8668 29257 8677 29291
rect 8677 29257 8711 29291
rect 8711 29257 8720 29291
rect 8668 29248 8720 29257
rect 4528 29180 4580 29232
rect 7012 29180 7064 29232
rect 8392 29180 8444 29232
rect 5264 29155 5316 29164
rect 5264 29121 5273 29155
rect 5273 29121 5307 29155
rect 5307 29121 5316 29155
rect 5264 29112 5316 29121
rect 7104 29112 7156 29164
rect 7196 29112 7248 29164
rect 8852 29112 8904 29164
rect 7288 29087 7340 29096
rect 7288 29053 7297 29087
rect 7297 29053 7331 29087
rect 7331 29053 7340 29087
rect 7288 29044 7340 29053
rect 5632 28976 5684 29028
rect 7932 29044 7984 29096
rect 8300 29044 8352 29096
rect 10232 29248 10284 29300
rect 11888 29291 11940 29300
rect 11888 29257 11897 29291
rect 11897 29257 11931 29291
rect 11931 29257 11940 29291
rect 11888 29248 11940 29257
rect 11980 29044 12032 29096
rect 6644 28908 6696 28960
rect 10600 28908 10652 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 7196 28704 7248 28756
rect 7932 28704 7984 28756
rect 9312 28704 9364 28756
rect 9956 28747 10008 28756
rect 9956 28713 9965 28747
rect 9965 28713 9999 28747
rect 9999 28713 10008 28747
rect 9956 28704 10008 28713
rect 8668 28636 8720 28688
rect 4896 28568 4948 28620
rect 6184 28611 6236 28620
rect 6184 28577 6193 28611
rect 6193 28577 6227 28611
rect 6227 28577 6236 28611
rect 6184 28568 6236 28577
rect 6644 28611 6696 28620
rect 6644 28577 6653 28611
rect 6653 28577 6687 28611
rect 6687 28577 6696 28611
rect 6644 28568 6696 28577
rect 6828 28543 6880 28552
rect 6828 28509 6837 28543
rect 6837 28509 6871 28543
rect 6871 28509 6880 28543
rect 6828 28500 6880 28509
rect 7564 28568 7616 28620
rect 9680 28611 9732 28620
rect 9680 28577 9689 28611
rect 9689 28577 9723 28611
rect 9723 28577 9732 28611
rect 9680 28568 9732 28577
rect 10968 28568 11020 28620
rect 11060 28500 11112 28552
rect 8024 28432 8076 28484
rect 8392 28432 8444 28484
rect 4804 28364 4856 28416
rect 5264 28407 5316 28416
rect 5264 28373 5273 28407
rect 5273 28373 5307 28407
rect 5307 28373 5316 28407
rect 5264 28364 5316 28373
rect 5356 28364 5408 28416
rect 6736 28364 6788 28416
rect 9588 28364 9640 28416
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 4436 28203 4488 28212
rect 4436 28169 4445 28203
rect 4445 28169 4479 28203
rect 4479 28169 4488 28203
rect 4436 28160 4488 28169
rect 4896 28203 4948 28212
rect 4896 28169 4905 28203
rect 4905 28169 4939 28203
rect 4939 28169 4948 28203
rect 4896 28160 4948 28169
rect 6644 28160 6696 28212
rect 7564 28160 7616 28212
rect 8668 28160 8720 28212
rect 5632 28092 5684 28144
rect 8300 28092 8352 28144
rect 5356 28024 5408 28076
rect 6828 28067 6880 28076
rect 6828 28033 6837 28067
rect 6837 28033 6871 28067
rect 6871 28033 6880 28067
rect 6828 28024 6880 28033
rect 7472 28024 7524 28076
rect 9680 28024 9732 28076
rect 3516 27956 3568 28008
rect 4436 27956 4488 28008
rect 9588 27999 9640 28008
rect 9588 27965 9597 27999
rect 9597 27965 9631 27999
rect 9631 27965 9640 27999
rect 9588 27956 9640 27965
rect 11060 28203 11112 28212
rect 11060 28169 11069 28203
rect 11069 28169 11103 28203
rect 11103 28169 11112 28203
rect 11060 28160 11112 28169
rect 10600 28024 10652 28076
rect 3056 27888 3108 27940
rect 4896 27888 4948 27940
rect 5264 27888 5316 27940
rect 5908 27888 5960 27940
rect 8576 27888 8628 27940
rect 10968 27888 11020 27940
rect 6000 27820 6052 27872
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 4804 27659 4856 27668
rect 4804 27625 4813 27659
rect 4813 27625 4847 27659
rect 4847 27625 4856 27659
rect 4804 27616 4856 27625
rect 5264 27616 5316 27668
rect 6828 27616 6880 27668
rect 5356 27548 5408 27600
rect 5632 27548 5684 27600
rect 6276 27548 6328 27600
rect 9864 27591 9916 27600
rect 9864 27557 9873 27591
rect 9873 27557 9907 27591
rect 9907 27557 9916 27591
rect 9864 27548 9916 27557
rect 11980 27548 12032 27600
rect 4528 27480 4580 27532
rect 8208 27480 8260 27532
rect 8760 27480 8812 27532
rect 12440 27480 12492 27532
rect 13268 27480 13320 27532
rect 5724 27412 5776 27464
rect 7840 27412 7892 27464
rect 9404 27412 9456 27464
rect 11152 27412 11204 27464
rect 11520 27412 11572 27464
rect 5908 27387 5960 27396
rect 5908 27353 5917 27387
rect 5917 27353 5951 27387
rect 5951 27353 5960 27387
rect 5908 27344 5960 27353
rect 7472 27387 7524 27396
rect 7472 27353 7481 27387
rect 7481 27353 7515 27387
rect 7515 27353 7524 27387
rect 7472 27344 7524 27353
rect 6184 27276 6236 27328
rect 6644 27276 6696 27328
rect 8392 27276 8444 27328
rect 8852 27276 8904 27328
rect 9588 27276 9640 27328
rect 12532 27276 12584 27328
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 5724 27072 5776 27124
rect 6276 27115 6328 27124
rect 6276 27081 6285 27115
rect 6285 27081 6319 27115
rect 6319 27081 6328 27115
rect 6276 27072 6328 27081
rect 7840 27115 7892 27124
rect 7840 27081 7849 27115
rect 7849 27081 7883 27115
rect 7883 27081 7892 27115
rect 7840 27072 7892 27081
rect 13636 27072 13688 27124
rect 4160 27004 4212 27056
rect 4528 27047 4580 27056
rect 4528 27013 4537 27047
rect 4537 27013 4571 27047
rect 4571 27013 4580 27047
rect 4528 27004 4580 27013
rect 7472 27047 7524 27056
rect 4804 26936 4856 26988
rect 7472 27013 7481 27047
rect 7481 27013 7515 27047
rect 7515 27013 7524 27047
rect 7472 27004 7524 27013
rect 11152 27004 11204 27056
rect 6000 26936 6052 26988
rect 7104 26936 7156 26988
rect 9864 26936 9916 26988
rect 3240 26868 3292 26920
rect 4620 26868 4672 26920
rect 6184 26868 6236 26920
rect 4988 26800 5040 26852
rect 5264 26843 5316 26852
rect 5264 26809 5273 26843
rect 5273 26809 5307 26843
rect 5307 26809 5316 26843
rect 5264 26800 5316 26809
rect 3240 26732 3292 26784
rect 4620 26732 4672 26784
rect 8116 26868 8168 26920
rect 11060 26868 11112 26920
rect 12256 26868 12308 26920
rect 12716 26868 12768 26920
rect 9496 26800 9548 26852
rect 9772 26843 9824 26852
rect 9772 26809 9781 26843
rect 9781 26809 9815 26843
rect 9815 26809 9824 26843
rect 9772 26800 9824 26809
rect 11520 26800 11572 26852
rect 8760 26732 8812 26784
rect 11060 26732 11112 26784
rect 11980 26775 12032 26784
rect 11980 26741 11989 26775
rect 11989 26741 12023 26775
rect 12023 26741 12032 26775
rect 11980 26732 12032 26741
rect 12072 26732 12124 26784
rect 13268 26775 13320 26784
rect 13268 26741 13277 26775
rect 13277 26741 13311 26775
rect 13311 26741 13320 26775
rect 13268 26732 13320 26741
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 5632 26571 5684 26580
rect 5632 26537 5641 26571
rect 5641 26537 5675 26571
rect 5675 26537 5684 26571
rect 5632 26528 5684 26537
rect 5724 26528 5776 26580
rect 7104 26571 7156 26580
rect 7104 26537 7113 26571
rect 7113 26537 7147 26571
rect 7147 26537 7156 26571
rect 7104 26528 7156 26537
rect 10048 26528 10100 26580
rect 4160 26460 4212 26512
rect 6184 26460 6236 26512
rect 9864 26503 9916 26512
rect 9864 26469 9873 26503
rect 9873 26469 9907 26503
rect 9907 26469 9916 26503
rect 9864 26460 9916 26469
rect 12624 26460 12676 26512
rect 7840 26435 7892 26444
rect 7840 26401 7849 26435
rect 7849 26401 7883 26435
rect 7883 26401 7892 26435
rect 7840 26392 7892 26401
rect 8300 26435 8352 26444
rect 8300 26401 8309 26435
rect 8309 26401 8343 26435
rect 8343 26401 8352 26435
rect 8300 26392 8352 26401
rect 13084 26435 13136 26444
rect 13084 26401 13093 26435
rect 13093 26401 13127 26435
rect 13127 26401 13136 26435
rect 13084 26392 13136 26401
rect 4804 26324 4856 26376
rect 4988 26324 5040 26376
rect 6460 26324 6512 26376
rect 8392 26367 8444 26376
rect 8392 26333 8401 26367
rect 8401 26333 8435 26367
rect 8435 26333 8444 26367
rect 8392 26324 8444 26333
rect 9956 26324 10008 26376
rect 11060 26324 11112 26376
rect 11704 26324 11756 26376
rect 12072 26324 12124 26376
rect 12256 26324 12308 26376
rect 5356 26256 5408 26308
rect 5908 26256 5960 26308
rect 9404 26256 9456 26308
rect 11244 26256 11296 26308
rect 2872 26188 2924 26240
rect 5540 26188 5592 26240
rect 7196 26188 7248 26240
rect 7656 26188 7708 26240
rect 9496 26231 9548 26240
rect 9496 26197 9505 26231
rect 9505 26197 9539 26231
rect 9539 26197 9548 26231
rect 9496 26188 9548 26197
rect 10692 26231 10744 26240
rect 10692 26197 10701 26231
rect 10701 26197 10735 26231
rect 10735 26197 10744 26231
rect 10692 26188 10744 26197
rect 11152 26231 11204 26240
rect 11152 26197 11161 26231
rect 11161 26197 11195 26231
rect 11195 26197 11204 26231
rect 11152 26188 11204 26197
rect 12624 26188 12676 26240
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 5264 25984 5316 26036
rect 6460 26027 6512 26036
rect 6460 25993 6469 26027
rect 6469 25993 6503 26027
rect 6503 25993 6512 26027
rect 6460 25984 6512 25993
rect 2964 25916 3016 25968
rect 6920 25984 6972 26036
rect 8300 25984 8352 26036
rect 9864 25984 9916 26036
rect 11704 26027 11756 26036
rect 11704 25993 11713 26027
rect 11713 25993 11747 26027
rect 11747 25993 11756 26027
rect 11704 25984 11756 25993
rect 13084 25984 13136 26036
rect 2688 25848 2740 25900
rect 7840 25916 7892 25968
rect 8208 25959 8260 25968
rect 8208 25925 8217 25959
rect 8217 25925 8251 25959
rect 8251 25925 8260 25959
rect 8208 25916 8260 25925
rect 9312 25916 9364 25968
rect 9772 25916 9824 25968
rect 11152 25916 11204 25968
rect 6736 25848 6788 25900
rect 8392 25848 8444 25900
rect 3976 25780 4028 25832
rect 7656 25780 7708 25832
rect 4160 25755 4212 25764
rect 4160 25721 4169 25755
rect 4169 25721 4203 25755
rect 4203 25721 4212 25755
rect 4160 25712 4212 25721
rect 8208 25712 8260 25764
rect 12532 25891 12584 25900
rect 12532 25857 12541 25891
rect 12541 25857 12575 25891
rect 12575 25857 12584 25891
rect 12532 25848 12584 25857
rect 9864 25780 9916 25832
rect 10692 25780 10744 25832
rect 10416 25712 10468 25764
rect 11336 25755 11388 25764
rect 11336 25721 11345 25755
rect 11345 25721 11379 25755
rect 11379 25721 11388 25755
rect 12624 25755 12676 25764
rect 11336 25712 11388 25721
rect 12624 25721 12633 25755
rect 12633 25721 12667 25755
rect 12667 25721 12676 25755
rect 12624 25712 12676 25721
rect 4804 25644 4856 25696
rect 6092 25687 6144 25696
rect 6092 25653 6101 25687
rect 6101 25653 6135 25687
rect 6135 25653 6144 25687
rect 6092 25644 6144 25653
rect 12256 25687 12308 25696
rect 12256 25653 12265 25687
rect 12265 25653 12299 25687
rect 12299 25653 12308 25687
rect 12256 25644 12308 25653
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 4160 25440 4212 25492
rect 5264 25483 5316 25492
rect 5264 25449 5273 25483
rect 5273 25449 5307 25483
rect 5307 25449 5316 25483
rect 5264 25440 5316 25449
rect 6092 25440 6144 25492
rect 8392 25483 8444 25492
rect 8392 25449 8401 25483
rect 8401 25449 8435 25483
rect 8435 25449 8444 25483
rect 8392 25440 8444 25449
rect 8852 25440 8904 25492
rect 9956 25483 10008 25492
rect 9956 25449 9965 25483
rect 9965 25449 9999 25483
rect 9999 25449 10008 25483
rect 9956 25440 10008 25449
rect 10416 25483 10468 25492
rect 10416 25449 10425 25483
rect 10425 25449 10459 25483
rect 10459 25449 10468 25483
rect 10416 25440 10468 25449
rect 11336 25440 11388 25492
rect 12532 25440 12584 25492
rect 6736 25372 6788 25424
rect 8208 25372 8260 25424
rect 11796 25372 11848 25424
rect 2688 25347 2740 25356
rect 2688 25313 2697 25347
rect 2697 25313 2731 25347
rect 2731 25313 2740 25347
rect 2688 25304 2740 25313
rect 2872 25347 2924 25356
rect 2872 25313 2881 25347
rect 2881 25313 2915 25347
rect 2915 25313 2924 25347
rect 2872 25304 2924 25313
rect 9864 25304 9916 25356
rect 10048 25347 10100 25356
rect 10048 25313 10057 25347
rect 10057 25313 10091 25347
rect 10091 25313 10100 25347
rect 10048 25304 10100 25313
rect 11980 25304 12032 25356
rect 13544 25347 13596 25356
rect 13544 25313 13553 25347
rect 13553 25313 13587 25347
rect 13587 25313 13596 25347
rect 13544 25304 13596 25313
rect 4344 25100 4396 25152
rect 8484 25279 8536 25288
rect 5908 25100 5960 25152
rect 8484 25245 8493 25279
rect 8493 25245 8527 25279
rect 8527 25245 8536 25279
rect 8484 25236 8536 25245
rect 12072 25236 12124 25288
rect 9496 25168 9548 25220
rect 7288 25100 7340 25152
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 2688 24896 2740 24948
rect 2872 24939 2924 24948
rect 2872 24905 2881 24939
rect 2881 24905 2915 24939
rect 2915 24905 2924 24939
rect 2872 24896 2924 24905
rect 5264 24896 5316 24948
rect 6736 24896 6788 24948
rect 3976 24760 4028 24812
rect 5908 24803 5960 24812
rect 5908 24769 5917 24803
rect 5917 24769 5951 24803
rect 5951 24769 5960 24803
rect 5908 24760 5960 24769
rect 8484 24896 8536 24948
rect 10232 24896 10284 24948
rect 10416 24939 10468 24948
rect 10416 24905 10425 24939
rect 10425 24905 10459 24939
rect 10459 24905 10468 24939
rect 10416 24896 10468 24905
rect 10692 24896 10744 24948
rect 11796 24939 11848 24948
rect 11796 24905 11805 24939
rect 11805 24905 11839 24939
rect 11839 24905 11848 24939
rect 11796 24896 11848 24905
rect 13544 24939 13596 24948
rect 13544 24905 13553 24939
rect 13553 24905 13587 24939
rect 13587 24905 13596 24939
rect 13544 24896 13596 24905
rect 8852 24803 8904 24812
rect 8852 24769 8861 24803
rect 8861 24769 8895 24803
rect 8895 24769 8904 24803
rect 8852 24760 8904 24769
rect 11244 24760 11296 24812
rect 5632 24735 5684 24744
rect 4160 24624 4212 24676
rect 5632 24701 5641 24735
rect 5641 24701 5675 24735
rect 5675 24701 5684 24735
rect 5632 24692 5684 24701
rect 10508 24735 10560 24744
rect 10508 24701 10517 24735
rect 10517 24701 10551 24735
rect 10551 24701 10560 24735
rect 10508 24692 10560 24701
rect 13084 24760 13136 24812
rect 6644 24624 6696 24676
rect 3424 24599 3476 24608
rect 3424 24565 3433 24599
rect 3433 24565 3467 24599
rect 3467 24565 3476 24599
rect 3424 24556 3476 24565
rect 7288 24667 7340 24676
rect 7288 24633 7297 24667
rect 7297 24633 7331 24667
rect 7331 24633 7340 24667
rect 7288 24624 7340 24633
rect 7656 24624 7708 24676
rect 9312 24624 9364 24676
rect 10416 24624 10468 24676
rect 12900 24735 12952 24744
rect 12900 24701 12909 24735
rect 12909 24701 12943 24735
rect 12943 24701 12952 24735
rect 12900 24692 12952 24701
rect 10692 24624 10744 24676
rect 8116 24556 8168 24608
rect 11428 24599 11480 24608
rect 11428 24565 11437 24599
rect 11437 24565 11471 24599
rect 11471 24565 11480 24599
rect 11428 24556 11480 24565
rect 12532 24599 12584 24608
rect 12532 24565 12541 24599
rect 12541 24565 12575 24599
rect 12575 24565 12584 24599
rect 12532 24556 12584 24565
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 6092 24352 6144 24404
rect 8760 24352 8812 24404
rect 9680 24352 9732 24404
rect 10508 24352 10560 24404
rect 12532 24352 12584 24404
rect 4804 24327 4856 24336
rect 4804 24293 4813 24327
rect 4813 24293 4847 24327
rect 4847 24293 4856 24327
rect 4804 24284 4856 24293
rect 7288 24284 7340 24336
rect 11428 24284 11480 24336
rect 2964 24259 3016 24268
rect 2964 24225 2973 24259
rect 2973 24225 3007 24259
rect 3007 24225 3016 24259
rect 2964 24216 3016 24225
rect 3976 24216 4028 24268
rect 4160 24216 4212 24268
rect 6000 24259 6052 24268
rect 6000 24225 6009 24259
rect 6009 24225 6043 24259
rect 6043 24225 6052 24259
rect 6000 24216 6052 24225
rect 8576 24259 8628 24268
rect 8576 24225 8585 24259
rect 8585 24225 8619 24259
rect 8619 24225 8628 24259
rect 8576 24216 8628 24225
rect 9772 24216 9824 24268
rect 10048 24216 10100 24268
rect 12624 24259 12676 24268
rect 12624 24225 12633 24259
rect 12633 24225 12667 24259
rect 12667 24225 12676 24259
rect 12624 24216 12676 24225
rect 7932 24148 7984 24200
rect 11244 24148 11296 24200
rect 11520 24148 11572 24200
rect 11796 24191 11848 24200
rect 11796 24157 11805 24191
rect 11805 24157 11839 24191
rect 11839 24157 11848 24191
rect 11796 24148 11848 24157
rect 12900 24148 12952 24200
rect 4896 24080 4948 24132
rect 5540 24080 5592 24132
rect 7656 24123 7708 24132
rect 7656 24089 7665 24123
rect 7665 24089 7699 24123
rect 7699 24089 7708 24123
rect 7656 24080 7708 24089
rect 8208 24080 8260 24132
rect 2412 24012 2464 24064
rect 3424 24012 3476 24064
rect 4160 24012 4212 24064
rect 5632 24055 5684 24064
rect 5632 24021 5641 24055
rect 5641 24021 5675 24055
rect 5675 24021 5684 24055
rect 5632 24012 5684 24021
rect 6828 24055 6880 24064
rect 6828 24021 6837 24055
rect 6837 24021 6871 24055
rect 6871 24021 6880 24055
rect 6828 24012 6880 24021
rect 7196 24012 7248 24064
rect 8852 24012 8904 24064
rect 9404 24080 9456 24132
rect 9588 24012 9640 24064
rect 12072 24055 12124 24064
rect 12072 24021 12081 24055
rect 12081 24021 12115 24055
rect 12115 24021 12124 24055
rect 12072 24012 12124 24021
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 3976 23808 4028 23860
rect 8208 23808 8260 23860
rect 8392 23808 8444 23860
rect 8576 23808 8628 23860
rect 11428 23808 11480 23860
rect 2964 23740 3016 23792
rect 4068 23740 4120 23792
rect 6736 23740 6788 23792
rect 4344 23715 4396 23724
rect 4344 23681 4353 23715
rect 4353 23681 4387 23715
rect 4387 23681 4396 23715
rect 4344 23672 4396 23681
rect 6828 23715 6880 23724
rect 6828 23681 6837 23715
rect 6837 23681 6871 23715
rect 6871 23681 6880 23715
rect 6828 23672 6880 23681
rect 3148 23604 3200 23656
rect 3332 23604 3384 23656
rect 4160 23647 4212 23656
rect 4160 23613 4169 23647
rect 4169 23613 4203 23647
rect 4203 23613 4212 23647
rect 4160 23604 4212 23613
rect 2964 23536 3016 23588
rect 3424 23536 3476 23588
rect 4344 23536 4396 23588
rect 4436 23536 4488 23588
rect 5540 23604 5592 23656
rect 5632 23604 5684 23656
rect 6184 23604 6236 23656
rect 7656 23740 7708 23792
rect 8668 23715 8720 23724
rect 8668 23681 8677 23715
rect 8677 23681 8711 23715
rect 8711 23681 8720 23715
rect 8668 23672 8720 23681
rect 8852 23672 8904 23724
rect 10600 23740 10652 23792
rect 12624 23783 12676 23792
rect 12624 23749 12633 23783
rect 12633 23749 12667 23783
rect 12667 23749 12676 23783
rect 12624 23740 12676 23749
rect 12072 23672 12124 23724
rect 12256 23672 12308 23724
rect 12440 23672 12492 23724
rect 10416 23647 10468 23656
rect 5908 23579 5960 23588
rect 5908 23545 5917 23579
rect 5917 23545 5951 23579
rect 5951 23545 5960 23579
rect 5908 23536 5960 23545
rect 6000 23536 6052 23588
rect 6736 23536 6788 23588
rect 6920 23536 6972 23588
rect 3148 23511 3200 23520
rect 3148 23477 3157 23511
rect 3157 23477 3191 23511
rect 3191 23477 3200 23511
rect 3148 23468 3200 23477
rect 4896 23468 4948 23520
rect 8852 23536 8904 23588
rect 10416 23613 10425 23647
rect 10425 23613 10459 23647
rect 10459 23613 10468 23647
rect 10416 23604 10468 23613
rect 9772 23468 9824 23520
rect 10324 23468 10376 23520
rect 11244 23604 11296 23656
rect 11796 23536 11848 23588
rect 12164 23468 12216 23520
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 4344 23307 4396 23316
rect 4344 23273 4353 23307
rect 4353 23273 4387 23307
rect 4387 23273 4396 23307
rect 4344 23264 4396 23273
rect 5908 23264 5960 23316
rect 7288 23307 7340 23316
rect 4988 23239 5040 23248
rect 4988 23205 4997 23239
rect 4997 23205 5031 23239
rect 5031 23205 5040 23239
rect 4988 23196 5040 23205
rect 2872 23128 2924 23180
rect 7288 23273 7297 23307
rect 7297 23273 7331 23307
rect 7331 23273 7340 23307
rect 7288 23264 7340 23273
rect 7932 23307 7984 23316
rect 7932 23273 7941 23307
rect 7941 23273 7975 23307
rect 7975 23273 7984 23307
rect 7932 23264 7984 23273
rect 9496 23264 9548 23316
rect 10324 23264 10376 23316
rect 10692 23264 10744 23316
rect 12348 23264 12400 23316
rect 6920 23196 6972 23248
rect 7840 23196 7892 23248
rect 8852 23196 8904 23248
rect 11520 23196 11572 23248
rect 12164 23196 12216 23248
rect 8116 23171 8168 23180
rect 8116 23137 8125 23171
rect 8125 23137 8159 23171
rect 8159 23137 8168 23171
rect 8116 23128 8168 23137
rect 9680 23171 9732 23180
rect 9680 23137 9689 23171
rect 9689 23137 9723 23171
rect 9723 23137 9732 23171
rect 9680 23128 9732 23137
rect 3516 23060 3568 23112
rect 5356 23060 5408 23112
rect 5540 23103 5592 23112
rect 5540 23069 5549 23103
rect 5549 23069 5583 23103
rect 5583 23069 5592 23103
rect 5540 23060 5592 23069
rect 7196 23060 7248 23112
rect 11428 23060 11480 23112
rect 3148 22967 3200 22976
rect 3148 22933 3157 22967
rect 3157 22933 3191 22967
rect 3191 22933 3200 22967
rect 3148 22924 3200 22933
rect 3332 22924 3384 22976
rect 4344 22924 4396 22976
rect 4804 22924 4856 22976
rect 7012 22924 7064 22976
rect 8484 22924 8536 22976
rect 8852 22924 8904 22976
rect 9588 22924 9640 22976
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 2872 22720 2924 22772
rect 3516 22763 3568 22772
rect 3516 22729 3525 22763
rect 3525 22729 3559 22763
rect 3559 22729 3568 22763
rect 3516 22720 3568 22729
rect 4068 22763 4120 22772
rect 4068 22729 4077 22763
rect 4077 22729 4111 22763
rect 4111 22729 4120 22763
rect 4068 22720 4120 22729
rect 4988 22720 5040 22772
rect 5448 22720 5500 22772
rect 6920 22720 6972 22772
rect 11428 22763 11480 22772
rect 11428 22729 11437 22763
rect 11437 22729 11471 22763
rect 11471 22729 11480 22763
rect 11428 22720 11480 22729
rect 12348 22720 12400 22772
rect 4712 22652 4764 22704
rect 7012 22652 7064 22704
rect 7472 22652 7524 22704
rect 8300 22652 8352 22704
rect 7196 22627 7248 22636
rect 7196 22593 7205 22627
rect 7205 22593 7239 22627
rect 7239 22593 7248 22627
rect 7196 22584 7248 22593
rect 8116 22584 8168 22636
rect 9404 22584 9456 22636
rect 9772 22584 9824 22636
rect 4068 22516 4120 22568
rect 4804 22516 4856 22568
rect 4988 22491 5040 22500
rect 4988 22457 4991 22491
rect 4991 22457 5025 22491
rect 5025 22457 5040 22491
rect 4988 22448 5040 22457
rect 7012 22491 7064 22500
rect 7012 22457 7021 22491
rect 7021 22457 7055 22491
rect 7055 22457 7064 22491
rect 7012 22448 7064 22457
rect 7196 22448 7248 22500
rect 8484 22516 8536 22568
rect 9588 22516 9640 22568
rect 9864 22516 9916 22568
rect 10048 22559 10100 22568
rect 10048 22525 10057 22559
rect 10057 22525 10091 22559
rect 10091 22525 10100 22559
rect 10232 22559 10284 22568
rect 10048 22516 10100 22525
rect 10232 22525 10241 22559
rect 10241 22525 10275 22559
rect 10275 22525 10284 22559
rect 10232 22516 10284 22525
rect 12072 22516 12124 22568
rect 12532 22516 12584 22568
rect 13452 22559 13504 22568
rect 13452 22525 13461 22559
rect 13461 22525 13495 22559
rect 13495 22525 13504 22559
rect 13452 22516 13504 22525
rect 9128 22491 9180 22500
rect 9128 22457 9137 22491
rect 9137 22457 9171 22491
rect 9171 22457 9180 22491
rect 9128 22448 9180 22457
rect 9404 22448 9456 22500
rect 12624 22448 12676 22500
rect 9496 22423 9548 22432
rect 9496 22389 9505 22423
rect 9505 22389 9539 22423
rect 9539 22389 9548 22423
rect 9496 22380 9548 22389
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 10048 22380 10100 22432
rect 11520 22380 11572 22432
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 4344 22219 4396 22228
rect 4344 22185 4353 22219
rect 4353 22185 4387 22219
rect 4387 22185 4396 22219
rect 4344 22176 4396 22185
rect 5448 22219 5500 22228
rect 5448 22185 5457 22219
rect 5457 22185 5491 22219
rect 5491 22185 5500 22219
rect 5448 22176 5500 22185
rect 7472 22176 7524 22228
rect 9128 22176 9180 22228
rect 10416 22219 10468 22228
rect 4988 22108 5040 22160
rect 6184 22108 6236 22160
rect 5908 22040 5960 22092
rect 8484 22040 8536 22092
rect 9772 22040 9824 22092
rect 10416 22185 10425 22219
rect 10425 22185 10459 22219
rect 10459 22185 10468 22219
rect 10416 22176 10468 22185
rect 11520 22176 11572 22228
rect 12532 22151 12584 22160
rect 12532 22117 12541 22151
rect 12541 22117 12575 22151
rect 12575 22117 12584 22151
rect 12532 22108 12584 22117
rect 11520 22040 11572 22092
rect 12072 22083 12124 22092
rect 12072 22049 12081 22083
rect 12081 22049 12115 22083
rect 12115 22049 12124 22083
rect 12072 22040 12124 22049
rect 4528 22015 4580 22024
rect 4528 21981 4537 22015
rect 4537 21981 4571 22015
rect 4571 21981 4580 22015
rect 4528 21972 4580 21981
rect 6828 22015 6880 22024
rect 6828 21981 6837 22015
rect 6837 21981 6871 22015
rect 6871 21981 6880 22015
rect 6828 21972 6880 21981
rect 6920 21972 6972 22024
rect 8760 22015 8812 22024
rect 8760 21981 8769 22015
rect 8769 21981 8803 22015
rect 8803 21981 8812 22015
rect 8760 21972 8812 21981
rect 12164 21904 12216 21956
rect 9864 21879 9916 21888
rect 9864 21845 9873 21879
rect 9873 21845 9907 21879
rect 9907 21845 9916 21879
rect 9864 21836 9916 21845
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 4988 21632 5040 21684
rect 5632 21632 5684 21684
rect 5908 21675 5960 21684
rect 5908 21641 5917 21675
rect 5917 21641 5951 21675
rect 5951 21641 5960 21675
rect 5908 21632 5960 21641
rect 6920 21607 6972 21616
rect 6920 21573 6929 21607
rect 6929 21573 6963 21607
rect 6963 21573 6972 21607
rect 6920 21564 6972 21573
rect 8852 21632 8904 21684
rect 10416 21632 10468 21684
rect 12624 21675 12676 21684
rect 12624 21641 12633 21675
rect 12633 21641 12667 21675
rect 12667 21641 12676 21675
rect 12624 21632 12676 21641
rect 8484 21607 8536 21616
rect 4436 21496 4488 21548
rect 4804 21539 4856 21548
rect 4804 21505 4813 21539
rect 4813 21505 4847 21539
rect 4847 21505 4856 21539
rect 4804 21496 4856 21505
rect 4344 21428 4396 21480
rect 8484 21573 8493 21607
rect 8493 21573 8527 21607
rect 8527 21573 8536 21607
rect 8484 21564 8536 21573
rect 8760 21564 8812 21616
rect 9680 21496 9732 21548
rect 3424 21360 3476 21412
rect 8760 21428 8812 21480
rect 9496 21428 9548 21480
rect 9864 21428 9916 21480
rect 10048 21428 10100 21480
rect 13452 21360 13504 21412
rect 3792 21335 3844 21344
rect 3792 21301 3801 21335
rect 3801 21301 3835 21335
rect 3835 21301 3844 21335
rect 3792 21292 3844 21301
rect 8300 21335 8352 21344
rect 8300 21301 8309 21335
rect 8309 21301 8343 21335
rect 8343 21301 8352 21335
rect 8300 21292 8352 21301
rect 9680 21292 9732 21344
rect 9956 21292 10008 21344
rect 10048 21292 10100 21344
rect 11520 21292 11572 21344
rect 12164 21335 12216 21344
rect 12164 21301 12173 21335
rect 12173 21301 12207 21335
rect 12207 21301 12216 21335
rect 12164 21292 12216 21301
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 3792 21088 3844 21140
rect 4528 21088 4580 21140
rect 6184 21088 6236 21140
rect 8300 21088 8352 21140
rect 10048 21088 10100 21140
rect 10232 21088 10284 21140
rect 11152 21088 11204 21140
rect 12072 21088 12124 21140
rect 4712 21020 4764 21072
rect 5908 21020 5960 21072
rect 6644 21020 6696 21072
rect 7472 21020 7524 21072
rect 8668 21020 8720 21072
rect 8760 21020 8812 21072
rect 9956 21020 10008 21072
rect 4344 20952 4396 21004
rect 7564 20952 7616 21004
rect 7840 20952 7892 21004
rect 9772 20995 9824 21004
rect 9772 20961 9781 20995
rect 9781 20961 9815 20995
rect 9815 20961 9824 20995
rect 9772 20952 9824 20961
rect 9864 20952 9916 21004
rect 11244 20995 11296 21004
rect 11244 20961 11253 20995
rect 11253 20961 11287 20995
rect 11287 20961 11296 20995
rect 11244 20952 11296 20961
rect 11520 20995 11572 21004
rect 11520 20961 11529 20995
rect 11529 20961 11563 20995
rect 11563 20961 11572 20995
rect 11520 20952 11572 20961
rect 3976 20884 4028 20936
rect 6276 20884 6328 20936
rect 8392 20884 8444 20936
rect 4344 20816 4396 20868
rect 7748 20816 7800 20868
rect 8024 20816 8076 20868
rect 9680 20816 9732 20868
rect 12072 20816 12124 20868
rect 6736 20748 6788 20800
rect 9956 20748 10008 20800
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 3516 20544 3568 20596
rect 3976 20544 4028 20596
rect 4528 20408 4580 20460
rect 4068 20272 4120 20324
rect 4712 20544 4764 20596
rect 6276 20587 6328 20596
rect 6276 20553 6285 20587
rect 6285 20553 6319 20587
rect 6319 20553 6328 20587
rect 6276 20544 6328 20553
rect 9772 20587 9824 20596
rect 9772 20553 9781 20587
rect 9781 20553 9815 20587
rect 9815 20553 9824 20587
rect 9772 20544 9824 20553
rect 11244 20544 11296 20596
rect 7472 20519 7524 20528
rect 7472 20485 7481 20519
rect 7481 20485 7515 20519
rect 7515 20485 7524 20519
rect 7472 20476 7524 20485
rect 9496 20476 9548 20528
rect 11060 20476 11112 20528
rect 14740 20476 14792 20528
rect 5540 20408 5592 20460
rect 6000 20408 6052 20460
rect 7840 20451 7892 20460
rect 7840 20417 7849 20451
rect 7849 20417 7883 20451
rect 7883 20417 7892 20451
rect 7840 20408 7892 20417
rect 8484 20408 8536 20460
rect 9404 20408 9456 20460
rect 8300 20383 8352 20392
rect 8300 20349 8309 20383
rect 8309 20349 8343 20383
rect 8343 20349 8352 20383
rect 8760 20383 8812 20392
rect 8300 20340 8352 20349
rect 8760 20349 8769 20383
rect 8769 20349 8803 20383
rect 8803 20349 8812 20383
rect 8760 20340 8812 20349
rect 9956 20383 10008 20392
rect 9956 20349 9965 20383
rect 9965 20349 9999 20383
rect 9999 20349 10008 20383
rect 9956 20340 10008 20349
rect 10140 20340 10192 20392
rect 11152 20340 11204 20392
rect 4804 20315 4856 20324
rect 4804 20281 4813 20315
rect 4813 20281 4847 20315
rect 4847 20281 4856 20315
rect 4804 20272 4856 20281
rect 4896 20315 4948 20324
rect 4896 20281 4905 20315
rect 4905 20281 4939 20315
rect 4939 20281 4948 20315
rect 4896 20272 4948 20281
rect 6736 20272 6788 20324
rect 7012 20315 7064 20324
rect 7012 20281 7021 20315
rect 7021 20281 7055 20315
rect 7055 20281 7064 20315
rect 10692 20315 10744 20324
rect 7012 20272 7064 20281
rect 10692 20281 10701 20315
rect 10701 20281 10735 20315
rect 10735 20281 10744 20315
rect 10692 20272 10744 20281
rect 11520 20272 11572 20324
rect 12256 20272 12308 20324
rect 4252 20247 4304 20256
rect 4252 20213 4261 20247
rect 4261 20213 4295 20247
rect 4295 20213 4304 20247
rect 4252 20204 4304 20213
rect 5080 20204 5132 20256
rect 6644 20247 6696 20256
rect 6644 20213 6653 20247
rect 6653 20213 6687 20247
rect 6687 20213 6696 20247
rect 6644 20204 6696 20213
rect 12072 20204 12124 20256
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 4804 20043 4856 20052
rect 4804 20009 4813 20043
rect 4813 20009 4847 20043
rect 4847 20009 4856 20043
rect 4804 20000 4856 20009
rect 4896 20000 4948 20052
rect 9496 20043 9548 20052
rect 3976 19864 4028 19916
rect 5540 19932 5592 19984
rect 5632 19932 5684 19984
rect 5908 19932 5960 19984
rect 9496 20009 9505 20043
rect 9505 20009 9539 20043
rect 9539 20009 9548 20043
rect 9496 20000 9548 20009
rect 9588 20000 9640 20052
rect 6644 19932 6696 19984
rect 7840 19932 7892 19984
rect 10968 19932 11020 19984
rect 4528 19864 4580 19916
rect 4160 19796 4212 19848
rect 5540 19839 5592 19848
rect 5540 19805 5549 19839
rect 5549 19805 5583 19839
rect 5583 19805 5592 19839
rect 5540 19796 5592 19805
rect 8300 19796 8352 19848
rect 9956 19864 10008 19916
rect 10140 19907 10192 19916
rect 10140 19873 10149 19907
rect 10149 19873 10183 19907
rect 10183 19873 10192 19907
rect 10140 19864 10192 19873
rect 10692 19864 10744 19916
rect 11520 19864 11572 19916
rect 10600 19796 10652 19848
rect 7932 19771 7984 19780
rect 7932 19737 7941 19771
rect 7941 19737 7975 19771
rect 7975 19737 7984 19771
rect 7932 19728 7984 19737
rect 9956 19771 10008 19780
rect 9956 19737 9965 19771
rect 9965 19737 9999 19771
rect 9999 19737 10008 19771
rect 9956 19728 10008 19737
rect 6920 19703 6972 19712
rect 6920 19669 6929 19703
rect 6929 19669 6963 19703
rect 6963 19669 6972 19703
rect 6920 19660 6972 19669
rect 7380 19660 7432 19712
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 3976 19456 4028 19508
rect 4896 19456 4948 19508
rect 7840 19499 7892 19508
rect 7840 19465 7849 19499
rect 7849 19465 7883 19499
rect 7883 19465 7892 19499
rect 7840 19456 7892 19465
rect 10140 19456 10192 19508
rect 11060 19456 11112 19508
rect 11520 19499 11572 19508
rect 11520 19465 11529 19499
rect 11529 19465 11563 19499
rect 11563 19465 11572 19499
rect 11520 19456 11572 19465
rect 3332 19388 3384 19440
rect 6736 19388 6788 19440
rect 4528 19320 4580 19372
rect 2412 19116 2464 19168
rect 3516 19252 3568 19304
rect 4252 19295 4304 19304
rect 4252 19261 4261 19295
rect 4261 19261 4295 19295
rect 4295 19261 4304 19295
rect 4252 19252 4304 19261
rect 5540 19252 5592 19304
rect 5632 19184 5684 19236
rect 7380 19320 7432 19372
rect 7932 19320 7984 19372
rect 11428 19388 11480 19440
rect 12440 19320 12492 19372
rect 9772 19252 9824 19304
rect 4528 19116 4580 19168
rect 5908 19116 5960 19168
rect 6644 19159 6696 19168
rect 6644 19125 6653 19159
rect 6653 19125 6687 19159
rect 6687 19125 6696 19159
rect 7656 19184 7708 19236
rect 9956 19184 10008 19236
rect 6644 19116 6696 19125
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 3332 18912 3384 18964
rect 3516 18912 3568 18964
rect 4252 18955 4304 18964
rect 2780 18887 2832 18896
rect 2780 18853 2789 18887
rect 2789 18853 2823 18887
rect 2823 18853 2832 18887
rect 4252 18921 4261 18955
rect 4261 18921 4295 18955
rect 4295 18921 4304 18955
rect 4252 18912 4304 18921
rect 5540 18912 5592 18964
rect 6184 18912 6236 18964
rect 8300 18955 8352 18964
rect 2780 18844 2832 18853
rect 5172 18844 5224 18896
rect 5724 18844 5776 18896
rect 5908 18887 5960 18896
rect 5908 18853 5911 18887
rect 5911 18853 5945 18887
rect 5945 18853 5960 18887
rect 5908 18844 5960 18853
rect 8300 18921 8309 18955
rect 8309 18921 8343 18955
rect 8343 18921 8352 18955
rect 8300 18912 8352 18921
rect 9588 18912 9640 18964
rect 9956 18912 10008 18964
rect 10600 18912 10652 18964
rect 6920 18844 6972 18896
rect 8024 18844 8076 18896
rect 2044 18776 2096 18828
rect 2964 18776 3016 18828
rect 4712 18776 4764 18828
rect 3332 18708 3384 18760
rect 7196 18776 7248 18828
rect 5724 18708 5776 18760
rect 7380 18751 7432 18760
rect 7380 18717 7389 18751
rect 7389 18717 7423 18751
rect 7423 18717 7432 18751
rect 7380 18708 7432 18717
rect 10140 18776 10192 18828
rect 11428 18776 11480 18828
rect 13084 18776 13136 18828
rect 9772 18751 9824 18760
rect 9772 18717 9781 18751
rect 9781 18717 9815 18751
rect 9815 18717 9824 18751
rect 9772 18708 9824 18717
rect 10416 18751 10468 18760
rect 10416 18717 10425 18751
rect 10425 18717 10459 18751
rect 10459 18717 10468 18751
rect 10416 18708 10468 18717
rect 10692 18708 10744 18760
rect 6736 18640 6788 18692
rect 7932 18683 7984 18692
rect 7932 18649 7941 18683
rect 7941 18649 7975 18683
rect 7975 18649 7984 18683
rect 7932 18640 7984 18649
rect 9680 18640 9732 18692
rect 10232 18640 10284 18692
rect 10784 18640 10836 18692
rect 2596 18572 2648 18624
rect 4988 18615 5040 18624
rect 4988 18581 4997 18615
rect 4997 18581 5031 18615
rect 5031 18581 5040 18615
rect 4988 18572 5040 18581
rect 6828 18615 6880 18624
rect 6828 18581 6837 18615
rect 6837 18581 6871 18615
rect 6871 18581 6880 18615
rect 6828 18572 6880 18581
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 2044 18411 2096 18420
rect 2044 18377 2053 18411
rect 2053 18377 2087 18411
rect 2087 18377 2096 18411
rect 2044 18368 2096 18377
rect 4344 18368 4396 18420
rect 4712 18368 4764 18420
rect 5908 18368 5960 18420
rect 8024 18411 8076 18420
rect 2780 18300 2832 18352
rect 2964 18343 3016 18352
rect 2964 18309 2973 18343
rect 2973 18309 3007 18343
rect 3007 18309 3016 18343
rect 2964 18300 3016 18309
rect 5448 18300 5500 18352
rect 4252 18232 4304 18284
rect 8024 18377 8033 18411
rect 8033 18377 8067 18411
rect 8067 18377 8076 18411
rect 8024 18368 8076 18377
rect 8484 18411 8536 18420
rect 8484 18377 8493 18411
rect 8493 18377 8527 18411
rect 8527 18377 8536 18411
rect 8484 18368 8536 18377
rect 9588 18411 9640 18420
rect 9588 18377 9597 18411
rect 9597 18377 9631 18411
rect 9631 18377 9640 18411
rect 9588 18368 9640 18377
rect 10140 18368 10192 18420
rect 11428 18411 11480 18420
rect 11428 18377 11437 18411
rect 11437 18377 11471 18411
rect 11471 18377 11480 18411
rect 11428 18368 11480 18377
rect 6644 18300 6696 18352
rect 9772 18300 9824 18352
rect 2504 18164 2556 18216
rect 2688 18164 2740 18216
rect 3332 18164 3384 18216
rect 3516 18164 3568 18216
rect 4344 18164 4396 18216
rect 4988 18207 5040 18216
rect 4988 18173 4997 18207
rect 4997 18173 5031 18207
rect 5031 18173 5040 18207
rect 4988 18164 5040 18173
rect 5540 18207 5592 18216
rect 5540 18173 5549 18207
rect 5549 18173 5583 18207
rect 5583 18173 5592 18207
rect 5540 18164 5592 18173
rect 5816 18164 5868 18216
rect 6828 18207 6880 18216
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 5724 18139 5776 18148
rect 5724 18105 5733 18139
rect 5733 18105 5767 18139
rect 5767 18105 5776 18139
rect 5724 18096 5776 18105
rect 7104 18232 7156 18284
rect 8024 18232 8076 18284
rect 9588 18232 9640 18284
rect 9864 18232 9916 18284
rect 11520 18232 11572 18284
rect 8576 18164 8628 18216
rect 10416 18164 10468 18216
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 9312 18139 9364 18148
rect 9312 18105 9321 18139
rect 9321 18105 9355 18139
rect 9355 18105 9364 18139
rect 9312 18096 9364 18105
rect 1400 18028 1452 18080
rect 3332 18028 3384 18080
rect 4712 18028 4764 18080
rect 9864 18028 9916 18080
rect 10784 18071 10836 18080
rect 10784 18037 10793 18071
rect 10793 18037 10827 18071
rect 10827 18037 10836 18071
rect 10784 18028 10836 18037
rect 10968 18028 11020 18080
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 3516 17867 3568 17876
rect 3516 17833 3525 17867
rect 3525 17833 3559 17867
rect 3559 17833 3568 17867
rect 3516 17824 3568 17833
rect 5632 17824 5684 17876
rect 5724 17824 5776 17876
rect 6644 17824 6696 17876
rect 9312 17867 9364 17876
rect 2596 17756 2648 17808
rect 5816 17799 5868 17808
rect 2964 17731 3016 17740
rect 2964 17697 2973 17731
rect 2973 17697 3007 17731
rect 3007 17697 3016 17731
rect 2964 17688 3016 17697
rect 4160 17731 4212 17740
rect 4160 17697 4178 17731
rect 4178 17697 4212 17731
rect 4160 17688 4212 17697
rect 5816 17765 5825 17799
rect 5825 17765 5859 17799
rect 5859 17765 5868 17799
rect 5816 17756 5868 17765
rect 6736 17799 6788 17808
rect 6736 17765 6745 17799
rect 6745 17765 6779 17799
rect 6779 17765 6788 17799
rect 6736 17756 6788 17765
rect 7472 17756 7524 17808
rect 9312 17833 9321 17867
rect 9321 17833 9355 17867
rect 9355 17833 9364 17867
rect 9312 17824 9364 17833
rect 9680 17824 9732 17876
rect 5264 17731 5316 17740
rect 5264 17697 5273 17731
rect 5273 17697 5307 17731
rect 5307 17697 5316 17731
rect 5264 17688 5316 17697
rect 5540 17731 5592 17740
rect 5540 17697 5549 17731
rect 5549 17697 5583 17731
rect 5583 17697 5592 17731
rect 5540 17688 5592 17697
rect 10600 17824 10652 17876
rect 10784 17799 10836 17808
rect 10784 17765 10793 17799
rect 10793 17765 10827 17799
rect 10827 17765 10836 17799
rect 10784 17756 10836 17765
rect 7380 17620 7432 17672
rect 8300 17620 8352 17672
rect 9772 17731 9824 17740
rect 9772 17697 9781 17731
rect 9781 17697 9815 17731
rect 9815 17697 9824 17731
rect 9772 17688 9824 17697
rect 11520 17731 11572 17740
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 12808 17731 12860 17740
rect 12808 17697 12817 17731
rect 12817 17697 12851 17731
rect 12851 17697 12860 17731
rect 12808 17688 12860 17697
rect 13084 17731 13136 17740
rect 13084 17697 13093 17731
rect 13093 17697 13127 17731
rect 13127 17697 13136 17731
rect 13084 17688 13136 17697
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 2504 17595 2556 17604
rect 2504 17561 2513 17595
rect 2513 17561 2547 17595
rect 2547 17561 2556 17595
rect 2504 17552 2556 17561
rect 6828 17552 6880 17604
rect 8852 17552 8904 17604
rect 12900 17595 12952 17604
rect 12900 17561 12909 17595
rect 12909 17561 12943 17595
rect 12943 17561 12952 17595
rect 12900 17552 12952 17561
rect 4712 17484 4764 17536
rect 8484 17527 8536 17536
rect 8484 17493 8493 17527
rect 8493 17493 8527 17527
rect 8527 17493 8536 17527
rect 8484 17484 8536 17493
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 5264 17323 5316 17332
rect 3148 17212 3200 17264
rect 3884 17212 3936 17264
rect 5264 17289 5273 17323
rect 5273 17289 5307 17323
rect 5307 17289 5316 17323
rect 5264 17280 5316 17289
rect 5540 17280 5592 17332
rect 8300 17323 8352 17332
rect 8300 17289 8309 17323
rect 8309 17289 8343 17323
rect 8343 17289 8352 17323
rect 8300 17280 8352 17289
rect 9772 17280 9824 17332
rect 11520 17280 11572 17332
rect 12808 17280 12860 17332
rect 2964 17144 3016 17196
rect 4068 17076 4120 17128
rect 4712 17119 4764 17128
rect 4712 17085 4721 17119
rect 4721 17085 4755 17119
rect 4755 17085 4764 17119
rect 4712 17076 4764 17085
rect 6184 17076 6236 17128
rect 4988 17051 5040 17060
rect 4988 17017 4997 17051
rect 4997 17017 5031 17051
rect 5031 17017 5040 17051
rect 4988 17008 5040 17017
rect 7196 17119 7248 17128
rect 7196 17085 7205 17119
rect 7205 17085 7239 17119
rect 7239 17085 7248 17119
rect 7196 17076 7248 17085
rect 13084 17212 13136 17264
rect 8576 17144 8628 17196
rect 8208 17076 8260 17128
rect 8944 17119 8996 17128
rect 8944 17085 8953 17119
rect 8953 17085 8987 17119
rect 8987 17085 8996 17119
rect 8944 17076 8996 17085
rect 9312 17119 9364 17128
rect 9312 17085 9321 17119
rect 9321 17085 9355 17119
rect 9355 17085 9364 17119
rect 9312 17076 9364 17085
rect 11520 17144 11572 17196
rect 11980 17144 12032 17196
rect 10600 17119 10652 17128
rect 10600 17085 10609 17119
rect 10609 17085 10643 17119
rect 10643 17085 10652 17119
rect 10600 17076 10652 17085
rect 10784 17076 10836 17128
rect 11244 17076 11296 17128
rect 7564 17008 7616 17060
rect 8300 17008 8352 17060
rect 4160 16983 4212 16992
rect 4160 16949 4169 16983
rect 4169 16949 4203 16983
rect 4203 16949 4212 16983
rect 11520 17008 11572 17060
rect 12900 17051 12952 17060
rect 12900 17017 12909 17051
rect 12909 17017 12943 17051
rect 12943 17017 12952 17051
rect 12900 17008 12952 17017
rect 14740 17008 14792 17060
rect 9772 16983 9824 16992
rect 4160 16940 4212 16949
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 11060 16983 11112 16992
rect 11060 16949 11069 16983
rect 11069 16949 11103 16983
rect 11103 16949 11112 16983
rect 11060 16940 11112 16949
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 3884 16736 3936 16788
rect 4068 16736 4120 16788
rect 4988 16736 5040 16788
rect 6736 16736 6788 16788
rect 6828 16736 6880 16788
rect 9312 16736 9364 16788
rect 10784 16779 10836 16788
rect 10784 16745 10793 16779
rect 10793 16745 10827 16779
rect 10827 16745 10836 16779
rect 10784 16736 10836 16745
rect 11336 16736 11388 16788
rect 8944 16668 8996 16720
rect 3424 16600 3476 16652
rect 4252 16643 4304 16652
rect 4252 16609 4261 16643
rect 4261 16609 4295 16643
rect 4295 16609 4304 16643
rect 4252 16600 4304 16609
rect 4712 16643 4764 16652
rect 4160 16532 4212 16584
rect 4712 16609 4721 16643
rect 4721 16609 4755 16643
rect 4755 16609 4764 16643
rect 4712 16600 4764 16609
rect 6644 16643 6696 16652
rect 6644 16609 6653 16643
rect 6653 16609 6687 16643
rect 6687 16609 6696 16643
rect 6644 16600 6696 16609
rect 7196 16600 7248 16652
rect 7564 16643 7616 16652
rect 7564 16609 7573 16643
rect 7573 16609 7607 16643
rect 7607 16609 7616 16643
rect 7564 16600 7616 16609
rect 7656 16643 7708 16652
rect 7656 16609 7665 16643
rect 7665 16609 7699 16643
rect 7699 16609 7708 16643
rect 7656 16600 7708 16609
rect 8208 16600 8260 16652
rect 10324 16668 10376 16720
rect 10968 16668 11020 16720
rect 12808 16668 12860 16720
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 10692 16600 10744 16652
rect 12348 16600 12400 16652
rect 13544 16643 13596 16652
rect 13544 16609 13553 16643
rect 13553 16609 13587 16643
rect 13587 16609 13596 16643
rect 13544 16600 13596 16609
rect 4804 16575 4856 16584
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 10140 16575 10192 16584
rect 10140 16541 10149 16575
rect 10149 16541 10183 16575
rect 10183 16541 10192 16575
rect 10140 16532 10192 16541
rect 10600 16532 10652 16584
rect 11244 16532 11296 16584
rect 12716 16532 12768 16584
rect 7196 16507 7248 16516
rect 7196 16473 7205 16507
rect 7205 16473 7239 16507
rect 7239 16473 7248 16507
rect 7196 16464 7248 16473
rect 10048 16464 10100 16516
rect 12900 16464 12952 16516
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 3516 16192 3568 16244
rect 4528 16235 4580 16244
rect 4528 16201 4537 16235
rect 4537 16201 4571 16235
rect 4571 16201 4580 16235
rect 4528 16192 4580 16201
rect 6644 16192 6696 16244
rect 7656 16192 7708 16244
rect 10048 16235 10100 16244
rect 10048 16201 10057 16235
rect 10057 16201 10091 16235
rect 10091 16201 10100 16235
rect 10048 16192 10100 16201
rect 4252 16124 4304 16176
rect 4988 16056 5040 16108
rect 5080 15988 5132 16040
rect 8760 16056 8812 16108
rect 7380 16031 7432 16040
rect 7380 15997 7389 16031
rect 7389 15997 7423 16031
rect 7423 15997 7432 16031
rect 7380 15988 7432 15997
rect 8852 16031 8904 16040
rect 8852 15997 8861 16031
rect 8861 15997 8895 16031
rect 8895 15997 8904 16031
rect 8852 15988 8904 15997
rect 9312 16031 9364 16040
rect 9312 15997 9321 16031
rect 9321 15997 9355 16031
rect 9355 15997 9364 16031
rect 9312 15988 9364 15997
rect 12164 16124 12216 16176
rect 11152 16056 11204 16108
rect 4528 15920 4580 15972
rect 10968 15963 11020 15972
rect 10968 15929 10977 15963
rect 10977 15929 11011 15963
rect 11011 15929 11020 15963
rect 10968 15920 11020 15929
rect 11980 15920 12032 15972
rect 13544 15963 13596 15972
rect 13544 15929 13553 15963
rect 13553 15929 13587 15963
rect 13587 15929 13596 15963
rect 13544 15920 13596 15929
rect 4252 15852 4304 15904
rect 5540 15895 5592 15904
rect 5540 15861 5549 15895
rect 5549 15861 5583 15895
rect 5583 15861 5592 15895
rect 5540 15852 5592 15861
rect 7288 15852 7340 15904
rect 9588 15895 9640 15904
rect 9588 15861 9597 15895
rect 9597 15861 9631 15895
rect 9631 15861 9640 15895
rect 9588 15852 9640 15861
rect 12348 15852 12400 15904
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 5080 15648 5132 15700
rect 4528 15580 4580 15632
rect 4988 15580 5040 15632
rect 5540 15580 5592 15632
rect 6552 15623 6604 15632
rect 6552 15589 6561 15623
rect 6561 15589 6595 15623
rect 6595 15589 6604 15623
rect 6552 15580 6604 15589
rect 7564 15648 7616 15700
rect 7196 15580 7248 15632
rect 4804 15512 4856 15564
rect 8852 15580 8904 15632
rect 8208 15555 8260 15564
rect 8208 15521 8217 15555
rect 8217 15521 8251 15555
rect 8251 15521 8260 15555
rect 9404 15648 9456 15700
rect 9956 15648 10008 15700
rect 11152 15691 11204 15700
rect 11152 15657 11161 15691
rect 11161 15657 11195 15691
rect 11195 15657 11204 15691
rect 11152 15648 11204 15657
rect 11796 15623 11848 15632
rect 8208 15512 8260 15521
rect 9772 15512 9824 15564
rect 9956 15512 10008 15564
rect 11796 15589 11805 15623
rect 11805 15589 11839 15623
rect 11839 15589 11848 15623
rect 11796 15580 11848 15589
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 4160 15308 4212 15360
rect 5540 15351 5592 15360
rect 5540 15317 5549 15351
rect 5549 15317 5583 15351
rect 5583 15317 5592 15351
rect 5540 15308 5592 15317
rect 5632 15308 5684 15360
rect 7656 15444 7708 15496
rect 8300 15444 8352 15496
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 7380 15308 7432 15360
rect 8576 15308 8628 15360
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 4804 15104 4856 15156
rect 6552 15147 6604 15156
rect 6552 15113 6561 15147
rect 6561 15113 6595 15147
rect 6595 15113 6604 15147
rect 6552 15104 6604 15113
rect 7656 15104 7708 15156
rect 9404 15147 9456 15156
rect 9404 15113 9413 15147
rect 9413 15113 9447 15147
rect 9447 15113 9456 15147
rect 9404 15104 9456 15113
rect 10324 15147 10376 15156
rect 10324 15113 10333 15147
rect 10333 15113 10367 15147
rect 10367 15113 10376 15147
rect 10324 15104 10376 15113
rect 10968 15104 11020 15156
rect 11796 15147 11848 15156
rect 11796 15113 11805 15147
rect 11805 15113 11839 15147
rect 11839 15113 11848 15147
rect 11796 15104 11848 15113
rect 4436 15036 4488 15088
rect 4988 15036 5040 15088
rect 2688 14943 2740 14952
rect 2688 14909 2697 14943
rect 2697 14909 2731 14943
rect 2731 14909 2740 14943
rect 2688 14900 2740 14909
rect 4160 14968 4212 15020
rect 8484 15036 8536 15088
rect 7196 15011 7248 15020
rect 7196 14977 7205 15011
rect 7205 14977 7239 15011
rect 7239 14977 7248 15011
rect 7196 14968 7248 14977
rect 8208 14900 8260 14952
rect 8576 14900 8628 14952
rect 11796 14900 11848 14952
rect 4436 14832 4488 14884
rect 5540 14832 5592 14884
rect 6920 14875 6972 14884
rect 6920 14841 6929 14875
rect 6929 14841 6963 14875
rect 6963 14841 6972 14875
rect 6920 14832 6972 14841
rect 4896 14807 4948 14816
rect 4896 14773 4905 14807
rect 4905 14773 4939 14807
rect 4939 14773 4948 14807
rect 4896 14764 4948 14773
rect 6736 14764 6788 14816
rect 11704 14832 11756 14884
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 8484 14807 8536 14816
rect 8484 14773 8493 14807
rect 8493 14773 8527 14807
rect 8527 14773 8536 14807
rect 8484 14764 8536 14773
rect 9864 14807 9916 14816
rect 9864 14773 9873 14807
rect 9873 14773 9907 14807
rect 9907 14773 9916 14807
rect 9864 14764 9916 14773
rect 10600 14764 10652 14816
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 2688 14560 2740 14612
rect 5908 14560 5960 14612
rect 6920 14560 6972 14612
rect 8852 14603 8904 14612
rect 8852 14569 8861 14603
rect 8861 14569 8895 14603
rect 8895 14569 8904 14603
rect 8852 14560 8904 14569
rect 9772 14560 9824 14612
rect 4712 14535 4764 14544
rect 4712 14501 4721 14535
rect 4721 14501 4755 14535
rect 4755 14501 4764 14535
rect 4712 14492 4764 14501
rect 4896 14492 4948 14544
rect 4988 14492 5040 14544
rect 6736 14535 6788 14544
rect 6736 14501 6745 14535
rect 6745 14501 6779 14535
rect 6779 14501 6788 14535
rect 6736 14492 6788 14501
rect 7104 14492 7156 14544
rect 9864 14492 9916 14544
rect 2964 14356 3016 14408
rect 4620 14399 4672 14408
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 5080 14399 5132 14408
rect 5080 14365 5089 14399
rect 5089 14365 5123 14399
rect 5123 14365 5132 14399
rect 5080 14356 5132 14365
rect 7748 14424 7800 14476
rect 8484 14424 8536 14476
rect 9588 14424 9640 14476
rect 11336 14424 11388 14476
rect 6368 14356 6420 14408
rect 11060 14356 11112 14408
rect 4436 14288 4488 14340
rect 7380 14288 7432 14340
rect 11336 14288 11388 14340
rect 13268 14288 13320 14340
rect 4252 14220 4304 14272
rect 4804 14220 4856 14272
rect 5264 14220 5316 14272
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 8576 14263 8628 14272
rect 8576 14229 8585 14263
rect 8585 14229 8619 14263
rect 8619 14229 8628 14263
rect 8576 14220 8628 14229
rect 10692 14220 10744 14272
rect 10968 14220 11020 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 4620 14059 4672 14068
rect 4620 14025 4629 14059
rect 4629 14025 4663 14059
rect 4663 14025 4672 14059
rect 4620 14016 4672 14025
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 7104 14059 7156 14068
rect 7104 14025 7113 14059
rect 7113 14025 7147 14059
rect 7147 14025 7156 14059
rect 7104 14016 7156 14025
rect 9496 14016 9548 14068
rect 9864 14016 9916 14068
rect 10968 14059 11020 14068
rect 10968 14025 10977 14059
rect 10977 14025 11011 14059
rect 11011 14025 11020 14059
rect 10968 14016 11020 14025
rect 11060 14016 11112 14068
rect 11520 14016 11572 14068
rect 10140 13948 10192 14000
rect 2688 13812 2740 13864
rect 3608 13855 3660 13864
rect 3608 13821 3617 13855
rect 3617 13821 3651 13855
rect 3651 13821 3660 13855
rect 3608 13812 3660 13821
rect 4436 13880 4488 13932
rect 7288 13923 7340 13932
rect 7288 13889 7297 13923
rect 7297 13889 7331 13923
rect 7331 13889 7340 13923
rect 7288 13880 7340 13889
rect 9496 13880 9548 13932
rect 5080 13812 5132 13864
rect 5264 13787 5316 13796
rect 5264 13753 5273 13787
rect 5273 13753 5307 13787
rect 5307 13753 5316 13787
rect 5264 13744 5316 13753
rect 5356 13787 5408 13796
rect 5356 13753 5365 13787
rect 5365 13753 5399 13787
rect 5399 13753 5408 13787
rect 5356 13744 5408 13753
rect 5816 13676 5868 13728
rect 7104 13744 7156 13796
rect 8116 13744 8168 13796
rect 9312 13744 9364 13796
rect 10600 13787 10652 13796
rect 8392 13676 8444 13728
rect 10600 13753 10609 13787
rect 10609 13753 10643 13787
rect 10643 13753 10652 13787
rect 10600 13744 10652 13753
rect 10692 13676 10744 13728
rect 11428 13719 11480 13728
rect 11428 13685 11437 13719
rect 11437 13685 11471 13719
rect 11471 13685 11480 13719
rect 11428 13676 11480 13685
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 3608 13515 3660 13524
rect 3608 13481 3617 13515
rect 3617 13481 3651 13515
rect 3651 13481 3660 13515
rect 3608 13472 3660 13481
rect 4620 13515 4672 13524
rect 4620 13481 4629 13515
rect 4629 13481 4663 13515
rect 4663 13481 4672 13515
rect 4620 13472 4672 13481
rect 7104 13472 7156 13524
rect 7748 13515 7800 13524
rect 7748 13481 7757 13515
rect 7757 13481 7791 13515
rect 7791 13481 7800 13515
rect 7748 13472 7800 13481
rect 5264 13404 5316 13456
rect 8208 13447 8260 13456
rect 3332 13336 3384 13388
rect 4252 13336 4304 13388
rect 4988 13336 5040 13388
rect 8208 13413 8217 13447
rect 8217 13413 8251 13447
rect 8251 13413 8260 13447
rect 8208 13404 8260 13413
rect 10048 13447 10100 13456
rect 10048 13413 10057 13447
rect 10057 13413 10091 13447
rect 10091 13413 10100 13447
rect 10048 13404 10100 13413
rect 10600 13447 10652 13456
rect 10600 13413 10609 13447
rect 10609 13413 10643 13447
rect 10643 13413 10652 13447
rect 10600 13404 10652 13413
rect 11428 13379 11480 13388
rect 11428 13345 11437 13379
rect 11437 13345 11471 13379
rect 11471 13345 11480 13379
rect 11428 13336 11480 13345
rect 6828 13311 6880 13320
rect 6828 13277 6837 13311
rect 6837 13277 6871 13311
rect 6871 13277 6880 13311
rect 6828 13268 6880 13277
rect 8852 13268 8904 13320
rect 9496 13268 9548 13320
rect 8024 13200 8076 13252
rect 4712 13132 4764 13184
rect 4896 13175 4948 13184
rect 4896 13141 4905 13175
rect 4905 13141 4939 13175
rect 4939 13141 4948 13175
rect 4896 13132 4948 13141
rect 6000 13175 6052 13184
rect 6000 13141 6009 13175
rect 6009 13141 6043 13175
rect 6043 13141 6052 13175
rect 6000 13132 6052 13141
rect 8760 13132 8812 13184
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 5080 12928 5132 12980
rect 4252 12860 4304 12912
rect 5172 12860 5224 12912
rect 4896 12792 4948 12844
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 4160 12767 4212 12776
rect 4160 12733 4169 12767
rect 4169 12733 4203 12767
rect 4203 12733 4212 12767
rect 4160 12724 4212 12733
rect 4528 12724 4580 12776
rect 4988 12767 5040 12776
rect 4988 12733 4997 12767
rect 4997 12733 5031 12767
rect 5031 12733 5040 12767
rect 4988 12724 5040 12733
rect 7104 12928 7156 12980
rect 8208 12928 8260 12980
rect 8392 12971 8444 12980
rect 8392 12937 8401 12971
rect 8401 12937 8435 12971
rect 8435 12937 8444 12971
rect 8392 12928 8444 12937
rect 11428 12971 11480 12980
rect 11428 12937 11437 12971
rect 11437 12937 11471 12971
rect 11471 12937 11480 12971
rect 11428 12928 11480 12937
rect 8024 12792 8076 12844
rect 10048 12792 10100 12844
rect 7840 12724 7892 12776
rect 10692 12767 10744 12776
rect 10692 12733 10701 12767
rect 10701 12733 10735 12767
rect 10735 12733 10744 12767
rect 10692 12724 10744 12733
rect 4068 12656 4120 12708
rect 4712 12656 4764 12708
rect 5356 12699 5408 12708
rect 5356 12665 5365 12699
rect 5365 12665 5399 12699
rect 5399 12665 5408 12699
rect 5356 12656 5408 12665
rect 6000 12656 6052 12708
rect 8668 12699 8720 12708
rect 8668 12665 8677 12699
rect 8677 12665 8711 12699
rect 8711 12665 8720 12699
rect 8668 12656 8720 12665
rect 3332 12588 3384 12640
rect 7104 12588 7156 12640
rect 7748 12631 7800 12640
rect 7748 12597 7757 12631
rect 7757 12597 7791 12631
rect 7791 12597 7800 12631
rect 7748 12588 7800 12597
rect 8392 12588 8444 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 4160 12384 4212 12436
rect 4712 12427 4764 12436
rect 4712 12393 4721 12427
rect 4721 12393 4755 12427
rect 4755 12393 4764 12427
rect 4712 12384 4764 12393
rect 6000 12427 6052 12436
rect 6000 12393 6009 12427
rect 6009 12393 6043 12427
rect 6043 12393 6052 12427
rect 6000 12384 6052 12393
rect 7656 12427 7708 12436
rect 7656 12393 7665 12427
rect 7665 12393 7699 12427
rect 7699 12393 7708 12427
rect 7656 12384 7708 12393
rect 10692 12427 10744 12436
rect 10692 12393 10701 12427
rect 10701 12393 10735 12427
rect 10735 12393 10744 12427
rect 10692 12384 10744 12393
rect 112 12316 164 12368
rect 5080 12359 5132 12368
rect 5080 12325 5089 12359
rect 5089 12325 5123 12359
rect 5123 12325 5132 12359
rect 5080 12316 5132 12325
rect 7012 12316 7064 12368
rect 7748 12316 7800 12368
rect 8208 12359 8260 12368
rect 8208 12325 8217 12359
rect 8217 12325 8251 12359
rect 8251 12325 8260 12359
rect 8208 12316 8260 12325
rect 8852 12316 8904 12368
rect 9496 12359 9548 12368
rect 9496 12325 9505 12359
rect 9505 12325 9539 12359
rect 9539 12325 9548 12359
rect 9496 12316 9548 12325
rect 2964 12248 3016 12300
rect 9956 12291 10008 12300
rect 9956 12257 9965 12291
rect 9965 12257 9999 12291
rect 9999 12257 10008 12291
rect 9956 12248 10008 12257
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 11428 12248 11480 12300
rect 4988 12223 5040 12232
rect 4988 12189 4997 12223
rect 4997 12189 5031 12223
rect 5031 12189 5040 12223
rect 4988 12180 5040 12189
rect 5632 12223 5684 12232
rect 5632 12189 5641 12223
rect 5641 12189 5675 12223
rect 5675 12189 5684 12223
rect 5632 12180 5684 12189
rect 6828 12180 6880 12232
rect 8576 12180 8628 12232
rect 8024 12112 8076 12164
rect 8760 12112 8812 12164
rect 6644 12044 6696 12096
rect 10324 12044 10376 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 5080 11840 5132 11892
rect 6828 11840 6880 11892
rect 7012 11883 7064 11892
rect 7012 11849 7021 11883
rect 7021 11849 7055 11883
rect 7055 11849 7064 11883
rect 7012 11840 7064 11849
rect 7104 11840 7156 11892
rect 8208 11840 8260 11892
rect 3516 11679 3568 11688
rect 3516 11645 3525 11679
rect 3525 11645 3559 11679
rect 3559 11645 3568 11679
rect 3516 11636 3568 11645
rect 4160 11636 4212 11688
rect 4252 11611 4304 11620
rect 4252 11577 4261 11611
rect 4261 11577 4295 11611
rect 4295 11577 4304 11611
rect 4252 11568 4304 11577
rect 4344 11568 4396 11620
rect 7656 11747 7708 11756
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 5816 11611 5868 11620
rect 5080 11500 5132 11552
rect 5816 11577 5825 11611
rect 5825 11577 5859 11611
rect 5859 11577 5868 11611
rect 5816 11568 5868 11577
rect 7104 11568 7156 11620
rect 8944 11772 8996 11824
rect 10416 11772 10468 11824
rect 11244 11636 11296 11688
rect 9496 11568 9548 11620
rect 9956 11568 10008 11620
rect 11428 11636 11480 11688
rect 8668 11500 8720 11552
rect 10140 11500 10192 11552
rect 11336 11500 11388 11552
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 2872 11160 2924 11212
rect 4160 11296 4212 11348
rect 4528 11296 4580 11348
rect 5080 11296 5132 11348
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 9496 11339 9548 11348
rect 9496 11305 9505 11339
rect 9505 11305 9539 11339
rect 9539 11305 9548 11339
rect 9496 11296 9548 11305
rect 7104 11228 7156 11280
rect 8116 11228 8168 11280
rect 10232 11228 10284 11280
rect 10416 11271 10468 11280
rect 10416 11237 10425 11271
rect 10425 11237 10459 11271
rect 10459 11237 10468 11271
rect 10416 11228 10468 11237
rect 11612 11228 11664 11280
rect 6644 11160 6696 11212
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 10600 11092 10652 11144
rect 11980 11092 12032 11144
rect 8760 11024 8812 11076
rect 4160 10956 4212 11008
rect 4988 10956 5040 11008
rect 7932 10956 7984 11008
rect 8116 10956 8168 11008
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 2412 10795 2464 10804
rect 2412 10761 2421 10795
rect 2421 10761 2455 10795
rect 2455 10761 2464 10795
rect 2412 10752 2464 10761
rect 2872 10795 2924 10804
rect 2872 10761 2881 10795
rect 2881 10761 2915 10795
rect 2915 10761 2924 10795
rect 2872 10752 2924 10761
rect 4160 10752 4212 10804
rect 4252 10752 4304 10804
rect 6644 10752 6696 10804
rect 7012 10752 7064 10804
rect 7104 10752 7156 10804
rect 10232 10795 10284 10804
rect 10232 10761 10241 10795
rect 10241 10761 10275 10795
rect 10275 10761 10284 10795
rect 10232 10752 10284 10761
rect 10600 10795 10652 10804
rect 10600 10761 10609 10795
rect 10609 10761 10643 10795
rect 10643 10761 10652 10795
rect 10600 10752 10652 10761
rect 11612 10795 11664 10804
rect 11612 10761 11621 10795
rect 11621 10761 11655 10795
rect 11655 10761 11664 10795
rect 11612 10752 11664 10761
rect 9404 10684 9456 10736
rect 3148 10616 3200 10668
rect 7288 10616 7340 10668
rect 10416 10616 10468 10668
rect 4436 10591 4488 10600
rect 4436 10557 4445 10591
rect 4445 10557 4479 10591
rect 4479 10557 4488 10591
rect 4436 10548 4488 10557
rect 7564 10548 7616 10600
rect 10876 10591 10928 10600
rect 10876 10557 10894 10591
rect 10894 10557 10928 10591
rect 10876 10548 10928 10557
rect 4528 10480 4580 10532
rect 7104 10480 7156 10532
rect 9312 10523 9364 10532
rect 9312 10489 9321 10523
rect 9321 10489 9355 10523
rect 9355 10489 9364 10523
rect 9312 10480 9364 10489
rect 9404 10523 9456 10532
rect 9404 10489 9413 10523
rect 9413 10489 9447 10523
rect 9447 10489 9456 10523
rect 9404 10480 9456 10489
rect 4068 10412 4120 10464
rect 5356 10455 5408 10464
rect 5356 10421 5365 10455
rect 5365 10421 5399 10455
rect 5399 10421 5408 10455
rect 5356 10412 5408 10421
rect 11980 10455 12032 10464
rect 11980 10421 11989 10455
rect 11989 10421 12023 10455
rect 12023 10421 12032 10455
rect 11980 10412 12032 10421
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 4344 10208 4396 10260
rect 4436 10208 4488 10260
rect 7104 10208 7156 10260
rect 7472 10251 7524 10260
rect 7472 10217 7481 10251
rect 7481 10217 7515 10251
rect 7515 10217 7524 10251
rect 7472 10208 7524 10217
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 5356 10140 5408 10192
rect 8116 10140 8168 10192
rect 8760 10183 8812 10192
rect 8760 10149 8769 10183
rect 8769 10149 8803 10183
rect 8803 10149 8812 10183
rect 8760 10140 8812 10149
rect 4712 10072 4764 10124
rect 9680 10072 9732 10124
rect 10048 10072 10100 10124
rect 3976 10004 4028 10056
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 7932 10004 7984 10056
rect 2596 9936 2648 9988
rect 8024 9936 8076 9988
rect 2964 9868 3016 9920
rect 4528 9868 4580 9920
rect 7564 9868 7616 9920
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 3976 9707 4028 9716
rect 3976 9673 3985 9707
rect 3985 9673 4019 9707
rect 4019 9673 4028 9707
rect 3976 9664 4028 9673
rect 4712 9707 4764 9716
rect 4712 9673 4721 9707
rect 4721 9673 4755 9707
rect 4755 9673 4764 9707
rect 4712 9664 4764 9673
rect 6092 9664 6144 9716
rect 8116 9707 8168 9716
rect 8116 9673 8125 9707
rect 8125 9673 8159 9707
rect 8159 9673 8168 9707
rect 8116 9664 8168 9673
rect 11980 9664 12032 9716
rect 2688 9596 2740 9648
rect 5816 9639 5868 9648
rect 2412 9528 2464 9580
rect 3240 9528 3292 9580
rect 5448 9528 5500 9580
rect 5816 9605 5825 9639
rect 5825 9605 5859 9639
rect 5859 9605 5868 9639
rect 5816 9596 5868 9605
rect 7932 9596 7984 9648
rect 7380 9528 7432 9580
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 5080 9460 5132 9512
rect 5356 9435 5408 9444
rect 5356 9401 5365 9435
rect 5365 9401 5399 9435
rect 5399 9401 5408 9435
rect 5356 9392 5408 9401
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 5080 9367 5132 9376
rect 5080 9333 5089 9367
rect 5089 9333 5123 9367
rect 5123 9333 5132 9367
rect 5080 9324 5132 9333
rect 5448 9324 5500 9376
rect 7104 9460 7156 9512
rect 8668 9528 8720 9580
rect 8484 9503 8536 9512
rect 8484 9469 8502 9503
rect 8502 9469 8536 9503
rect 8484 9460 8536 9469
rect 7196 9392 7248 9444
rect 7104 9324 7156 9376
rect 8668 9324 8720 9376
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 5356 9120 5408 9172
rect 7380 9120 7432 9172
rect 8576 9120 8628 9172
rect 4068 9052 4120 9104
rect 6184 9052 6236 9104
rect 7288 9095 7340 9104
rect 3516 8984 3568 9036
rect 4436 9027 4488 9036
rect 4436 8993 4445 9027
rect 4445 8993 4479 9027
rect 4479 8993 4488 9027
rect 4436 8984 4488 8993
rect 4712 9027 4764 9036
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 4712 8984 4764 8993
rect 7288 9061 7297 9095
rect 7297 9061 7331 9095
rect 7331 9061 7340 9095
rect 7288 9052 7340 9061
rect 7564 9052 7616 9104
rect 9680 9052 9732 9104
rect 7104 9027 7156 9036
rect 7104 8993 7113 9027
rect 7113 8993 7147 9027
rect 7147 8993 7156 9027
rect 7104 8984 7156 8993
rect 8300 8984 8352 9036
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 8852 8848 8904 8900
rect 5356 8823 5408 8832
rect 5356 8789 5365 8823
rect 5365 8789 5399 8823
rect 5399 8789 5408 8823
rect 5356 8780 5408 8789
rect 8208 8780 8260 8832
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 4896 8576 4948 8628
rect 6184 8619 6236 8628
rect 664 8508 716 8560
rect 4620 8508 4672 8560
rect 6184 8585 6193 8619
rect 6193 8585 6227 8619
rect 6227 8585 6236 8619
rect 6184 8576 6236 8585
rect 8300 8576 8352 8628
rect 4252 8372 4304 8424
rect 4712 8372 4764 8424
rect 5356 8372 5408 8424
rect 4344 8347 4396 8356
rect 4344 8313 4353 8347
rect 4353 8313 4387 8347
rect 4387 8313 4396 8347
rect 4344 8304 4396 8313
rect 4620 8304 4672 8356
rect 5264 8304 5316 8356
rect 3976 8236 4028 8288
rect 4160 8236 4212 8288
rect 4436 8236 4488 8288
rect 9956 8508 10008 8560
rect 8208 8440 8260 8492
rect 7012 8304 7064 8356
rect 7472 8372 7524 8424
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 8852 8372 8904 8424
rect 6644 8236 6696 8288
rect 8208 8236 8260 8288
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 3976 8032 4028 8084
rect 4252 8075 4304 8084
rect 4252 8041 4261 8075
rect 4261 8041 4295 8075
rect 4295 8041 4304 8075
rect 4252 8032 4304 8041
rect 4804 8075 4856 8084
rect 4804 8041 4813 8075
rect 4813 8041 4847 8075
rect 4847 8041 4856 8075
rect 4804 8032 4856 8041
rect 3056 7964 3108 8016
rect 7564 8032 7616 8084
rect 7656 8032 7708 8084
rect 4988 7896 5040 7948
rect 6092 7964 6144 8016
rect 6644 8007 6696 8016
rect 6644 7973 6653 8007
rect 6653 7973 6687 8007
rect 6687 7973 6696 8007
rect 6644 7964 6696 7973
rect 8208 8007 8260 8016
rect 8208 7973 8217 8007
rect 8217 7973 8251 8007
rect 8251 7973 8260 8007
rect 8208 7964 8260 7973
rect 8852 7964 8904 8016
rect 5356 7939 5408 7948
rect 5356 7905 5365 7939
rect 5365 7905 5399 7939
rect 5399 7905 5408 7939
rect 5356 7896 5408 7905
rect 9956 7939 10008 7948
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 4436 7828 4488 7880
rect 6092 7828 6144 7880
rect 6828 7828 6880 7880
rect 8484 7828 8536 7880
rect 9312 7828 9364 7880
rect 4160 7760 4212 7812
rect 9864 7760 9916 7812
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 6644 7488 6696 7540
rect 8208 7488 8260 7540
rect 6828 7420 6880 7472
rect 4068 7352 4120 7404
rect 4804 7352 4856 7404
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 3976 7284 4028 7336
rect 4528 7284 4580 7336
rect 4896 7216 4948 7268
rect 5448 7216 5500 7268
rect 9956 7488 10008 7540
rect 8944 7420 8996 7472
rect 9680 7420 9732 7472
rect 9496 7395 9548 7404
rect 9496 7361 9505 7395
rect 9505 7361 9539 7395
rect 9539 7361 9548 7395
rect 9496 7352 9548 7361
rect 9496 7216 9548 7268
rect 9772 7216 9824 7268
rect 4436 7148 4488 7200
rect 5632 7191 5684 7200
rect 5632 7157 5641 7191
rect 5641 7157 5675 7191
rect 5675 7157 5684 7191
rect 5632 7148 5684 7157
rect 7472 7191 7524 7200
rect 7472 7157 7481 7191
rect 7481 7157 7515 7191
rect 7515 7157 7524 7191
rect 7472 7148 7524 7157
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 4344 6944 4396 6996
rect 9496 6987 9548 6996
rect 9496 6953 9505 6987
rect 9505 6953 9539 6987
rect 9539 6953 9548 6987
rect 9496 6944 9548 6953
rect 2688 6876 2740 6928
rect 4988 6919 5040 6928
rect 4988 6885 4997 6919
rect 4997 6885 5031 6919
rect 5031 6885 5040 6919
rect 4988 6876 5040 6885
rect 5448 6876 5500 6928
rect 7564 6876 7616 6928
rect 9956 6876 10008 6928
rect 2504 6808 2556 6860
rect 3976 6808 4028 6860
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 4896 6808 4948 6860
rect 6184 6808 6236 6860
rect 7012 6808 7064 6860
rect 8208 6808 8260 6860
rect 4528 6740 4580 6792
rect 9588 6740 9640 6792
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 9864 6740 9916 6792
rect 3976 6672 4028 6724
rect 4804 6672 4856 6724
rect 5908 6672 5960 6724
rect 6000 6604 6052 6656
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 8484 6604 8536 6656
rect 9496 6604 9548 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 2504 6400 2556 6452
rect 2688 6400 2740 6452
rect 3240 6443 3292 6452
rect 3240 6409 3249 6443
rect 3249 6409 3283 6443
rect 3283 6409 3292 6443
rect 3240 6400 3292 6409
rect 4528 6443 4580 6452
rect 4528 6409 4537 6443
rect 4537 6409 4571 6443
rect 4571 6409 4580 6443
rect 4528 6400 4580 6409
rect 6184 6443 6236 6452
rect 6184 6409 6193 6443
rect 6193 6409 6227 6443
rect 6227 6409 6236 6443
rect 6184 6400 6236 6409
rect 8392 6400 8444 6452
rect 9404 6400 9456 6452
rect 9864 6375 9916 6384
rect 9864 6341 9873 6375
rect 9873 6341 9907 6375
rect 9907 6341 9916 6375
rect 9864 6332 9916 6341
rect 2320 6264 2372 6316
rect 2412 6196 2464 6248
rect 4160 6264 4212 6316
rect 4344 6264 4396 6316
rect 6092 6264 6144 6316
rect 3240 6196 3292 6248
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 9956 6264 10008 6316
rect 4160 6171 4212 6180
rect 4160 6137 4169 6171
rect 4169 6137 4203 6171
rect 4203 6137 4212 6171
rect 4160 6128 4212 6137
rect 5448 6128 5500 6180
rect 7472 6128 7524 6180
rect 9312 6171 9364 6180
rect 9312 6137 9321 6171
rect 9321 6137 9355 6171
rect 9355 6137 9364 6171
rect 9312 6128 9364 6137
rect 9404 6171 9456 6180
rect 9404 6137 9413 6171
rect 9413 6137 9447 6171
rect 9447 6137 9456 6171
rect 9404 6128 9456 6137
rect 4896 6103 4948 6112
rect 4896 6069 4905 6103
rect 4905 6069 4939 6103
rect 4939 6069 4948 6103
rect 4896 6060 4948 6069
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 9772 6060 9824 6112
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 2412 5899 2464 5908
rect 2412 5865 2421 5899
rect 2421 5865 2455 5899
rect 2455 5865 2464 5899
rect 2412 5856 2464 5865
rect 3976 5856 4028 5908
rect 7288 5899 7340 5908
rect 7288 5865 7297 5899
rect 7297 5865 7331 5899
rect 7331 5865 7340 5899
rect 7288 5856 7340 5865
rect 8208 5899 8260 5908
rect 8208 5865 8217 5899
rect 8217 5865 8251 5899
rect 8251 5865 8260 5899
rect 8208 5856 8260 5865
rect 9312 5899 9364 5908
rect 9312 5865 9321 5899
rect 9321 5865 9355 5899
rect 9355 5865 9364 5899
rect 9312 5856 9364 5865
rect 9496 5856 9548 5908
rect 5908 5788 5960 5840
rect 6184 5788 6236 5840
rect 4068 5763 4120 5772
rect 4068 5729 4077 5763
rect 4077 5729 4111 5763
rect 4111 5729 4120 5763
rect 4068 5720 4120 5729
rect 4344 5720 4396 5772
rect 5356 5720 5408 5772
rect 7196 5763 7248 5772
rect 7196 5729 7205 5763
rect 7205 5729 7239 5763
rect 7239 5729 7248 5763
rect 7196 5720 7248 5729
rect 7656 5763 7708 5772
rect 7656 5729 7665 5763
rect 7665 5729 7699 5763
rect 7699 5729 7708 5763
rect 7656 5720 7708 5729
rect 7748 5720 7800 5772
rect 9680 5763 9732 5772
rect 9680 5729 9724 5763
rect 9724 5729 9732 5763
rect 9680 5720 9732 5729
rect 5448 5652 5500 5704
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 5816 5652 5868 5704
rect 4896 5516 4948 5568
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 4068 5312 4120 5364
rect 5632 5312 5684 5364
rect 6184 5355 6236 5364
rect 6184 5321 6193 5355
rect 6193 5321 6227 5355
rect 6227 5321 6236 5355
rect 6184 5312 6236 5321
rect 7196 5312 7248 5364
rect 9680 5355 9732 5364
rect 9680 5321 9689 5355
rect 9689 5321 9723 5355
rect 9723 5321 9732 5355
rect 9680 5312 9732 5321
rect 13176 5312 13228 5364
rect 3332 5244 3384 5296
rect 5356 5244 5408 5296
rect 7656 5244 7708 5296
rect 9404 5244 9456 5296
rect 4988 5176 5040 5228
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 5724 5219 5776 5228
rect 5724 5185 5733 5219
rect 5733 5185 5767 5219
rect 5767 5185 5776 5219
rect 5724 5176 5776 5185
rect 8760 5176 8812 5228
rect 9312 5176 9364 5228
rect 3976 5108 4028 5160
rect 6736 5108 6788 5160
rect 10048 5108 10100 5160
rect 4712 5040 4764 5092
rect 5632 5040 5684 5092
rect 8392 5083 8444 5092
rect 8392 5049 8401 5083
rect 8401 5049 8435 5083
rect 8435 5049 8444 5083
rect 8392 5040 8444 5049
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 8208 5015 8260 5024
rect 8208 4981 8217 5015
rect 8217 4981 8251 5015
rect 8251 4981 8260 5015
rect 8208 4972 8260 4981
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 3976 4768 4028 4820
rect 4344 4811 4396 4820
rect 4344 4777 4353 4811
rect 4353 4777 4387 4811
rect 4387 4777 4396 4811
rect 4344 4768 4396 4777
rect 5724 4768 5776 4820
rect 5908 4768 5960 4820
rect 8208 4811 8260 4820
rect 8208 4777 8217 4811
rect 8217 4777 8251 4811
rect 8251 4777 8260 4811
rect 8208 4768 8260 4777
rect 2872 4700 2924 4752
rect 4804 4700 4856 4752
rect 4896 4700 4948 4752
rect 5448 4700 5500 4752
rect 7104 4743 7156 4752
rect 7104 4709 7113 4743
rect 7113 4709 7147 4743
rect 7147 4709 7156 4743
rect 7104 4700 7156 4709
rect 7472 4700 7524 4752
rect 7656 4700 7708 4752
rect 8392 4700 8444 4752
rect 3516 4632 3568 4684
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 5264 4632 5316 4684
rect 7288 4675 7340 4684
rect 7288 4641 7297 4675
rect 7297 4641 7331 4675
rect 7331 4641 7340 4675
rect 7288 4632 7340 4641
rect 9956 4632 10008 4684
rect 10968 4564 11020 4616
rect 3976 4496 4028 4548
rect 2688 4428 2740 4480
rect 8852 4428 8904 4480
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 4712 4224 4764 4276
rect 7288 4224 7340 4276
rect 8208 4224 8260 4276
rect 9956 4267 10008 4276
rect 3240 4156 3292 4208
rect 5816 4156 5868 4208
rect 5632 4088 5684 4140
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 2872 4020 2924 4072
rect 4896 4020 4948 4072
rect 112 3884 164 3936
rect 3516 3927 3568 3936
rect 3516 3893 3525 3927
rect 3525 3893 3559 3927
rect 3559 3893 3568 3927
rect 3516 3884 3568 3893
rect 3976 3952 4028 4004
rect 5356 3995 5408 4004
rect 5356 3961 5365 3995
rect 5365 3961 5399 3995
rect 5399 3961 5408 3995
rect 5356 3952 5408 3961
rect 5724 3952 5776 4004
rect 7656 3952 7708 4004
rect 9956 4233 9965 4267
rect 9965 4233 9999 4267
rect 9999 4233 10008 4267
rect 9956 4224 10008 4233
rect 8852 4156 8904 4208
rect 9772 4156 9824 4208
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 10876 4224 10928 4276
rect 10968 4267 11020 4276
rect 10968 4233 10977 4267
rect 10977 4233 11011 4267
rect 11011 4233 11020 4267
rect 10968 4224 11020 4233
rect 6092 3884 6144 3936
rect 8208 3884 8260 3936
rect 10692 3884 10744 3936
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 3976 3680 4028 3732
rect 5356 3723 5408 3732
rect 5356 3689 5365 3723
rect 5365 3689 5399 3723
rect 5399 3689 5408 3723
rect 5356 3680 5408 3689
rect 5632 3723 5684 3732
rect 5632 3689 5641 3723
rect 5641 3689 5675 3723
rect 5675 3689 5684 3723
rect 5632 3680 5684 3689
rect 7656 3680 7708 3732
rect 8300 3680 8352 3732
rect 2688 3612 2740 3664
rect 4896 3612 4948 3664
rect 6000 3655 6052 3664
rect 6000 3621 6009 3655
rect 6009 3621 6043 3655
rect 6043 3621 6052 3655
rect 6000 3612 6052 3621
rect 6092 3612 6144 3664
rect 8208 3655 8260 3664
rect 8208 3621 8217 3655
rect 8217 3621 8251 3655
rect 8251 3621 8260 3655
rect 8208 3612 8260 3621
rect 9220 3612 9272 3664
rect 2596 3544 2648 3596
rect 3148 3544 3200 3596
rect 5356 3544 5408 3596
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 10232 3544 10284 3596
rect 2504 3476 2556 3528
rect 6184 3476 6236 3528
rect 9404 3476 9456 3528
rect 6920 3408 6972 3460
rect 11244 3408 11296 3460
rect 11612 3408 11664 3460
rect 2780 3340 2832 3392
rect 3516 3340 3568 3392
rect 9312 3340 9364 3392
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 1124 3136 1176 3188
rect 2412 3136 2464 3188
rect 2596 3136 2648 3188
rect 2964 3136 3016 3188
rect 5356 3179 5408 3188
rect 4988 3068 5040 3120
rect 2688 3043 2740 3052
rect 2688 3009 2697 3043
rect 2697 3009 2731 3043
rect 2731 3009 2740 3043
rect 2688 3000 2740 3009
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 5356 3145 5365 3179
rect 5365 3145 5399 3179
rect 5399 3145 5408 3179
rect 5356 3136 5408 3145
rect 6000 3136 6052 3188
rect 6184 3179 6236 3188
rect 6184 3145 6193 3179
rect 6193 3145 6227 3179
rect 6227 3145 6236 3179
rect 6184 3136 6236 3145
rect 8208 3136 8260 3188
rect 9404 3136 9456 3188
rect 9680 3136 9732 3188
rect 10048 3136 10100 3188
rect 10232 3179 10284 3188
rect 10232 3145 10241 3179
rect 10241 3145 10275 3179
rect 10275 3145 10284 3179
rect 10232 3136 10284 3145
rect 11612 3179 11664 3188
rect 11612 3145 11621 3179
rect 11621 3145 11655 3179
rect 11655 3145 11664 3179
rect 11612 3136 11664 3145
rect 5540 3068 5592 3120
rect 8760 3111 8812 3120
rect 8300 3000 8352 3052
rect 8760 3077 8769 3111
rect 8769 3077 8803 3111
rect 8803 3077 8812 3111
rect 8760 3068 8812 3077
rect 2780 2907 2832 2916
rect 2780 2873 2789 2907
rect 2789 2873 2823 2907
rect 2823 2873 2832 2907
rect 2780 2864 2832 2873
rect 4896 2864 4948 2916
rect 9680 2975 9732 2984
rect 9680 2941 9689 2975
rect 9689 2941 9723 2975
rect 9723 2941 9732 2975
rect 9680 2932 9732 2941
rect 5908 2864 5960 2916
rect 8300 2907 8352 2916
rect 8300 2873 8309 2907
rect 8309 2873 8343 2907
rect 8343 2873 8352 2907
rect 8300 2864 8352 2873
rect 5080 2839 5132 2848
rect 5080 2805 5089 2839
rect 5089 2805 5123 2839
rect 5123 2805 5132 2839
rect 5080 2796 5132 2805
rect 12532 2864 12584 2916
rect 9864 2839 9916 2848
rect 9864 2805 9873 2839
rect 9873 2805 9907 2839
rect 9907 2805 9916 2839
rect 9864 2796 9916 2805
rect 10416 2796 10468 2848
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 3516 2635 3568 2644
rect 2504 2567 2556 2576
rect 2504 2533 2513 2567
rect 2513 2533 2547 2567
rect 2547 2533 2556 2567
rect 2504 2524 2556 2533
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 4160 2592 4212 2644
rect 6000 2592 6052 2644
rect 3240 2524 3292 2576
rect 2780 2388 2832 2440
rect 5080 2567 5132 2576
rect 5080 2533 5089 2567
rect 5089 2533 5123 2567
rect 5123 2533 5132 2567
rect 5080 2524 5132 2533
rect 6092 2524 6144 2576
rect 8208 2592 8260 2644
rect 15568 2592 15620 2644
rect 8668 2524 8720 2576
rect 7932 2456 7984 2508
rect 11428 2499 11480 2508
rect 11428 2465 11437 2499
rect 11437 2465 11471 2499
rect 11471 2465 11480 2499
rect 11428 2456 11480 2465
rect 13176 2499 13228 2508
rect 13176 2465 13185 2499
rect 13185 2465 13219 2499
rect 13219 2465 13228 2499
rect 13176 2456 13228 2465
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 10416 2388 10468 2440
rect 6736 2320 6788 2372
rect 3332 2252 3384 2304
rect 5908 2252 5960 2304
rect 11704 2320 11756 2372
rect 14648 2320 14700 2372
rect 8300 2252 8352 2304
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 3424 76 3476 128
rect 4804 76 4856 128
rect 7012 76 7064 128
rect 13728 76 13780 128
<< metal2 >>
rect 386 39658 442 40000
rect 1214 39704 1270 40000
rect 386 39630 704 39658
rect 386 39520 442 39630
rect 676 33454 704 39630
rect 1214 39652 1216 39704
rect 1268 39652 1270 39704
rect 1214 39520 1270 39652
rect 1400 39636 1452 39642
rect 1400 39578 1452 39584
rect 2134 39636 2190 40000
rect 3054 39658 3110 40000
rect 2134 39584 2136 39636
rect 2188 39584 2190 39636
rect 664 33448 716 33454
rect 664 33390 716 33396
rect 1412 18086 1440 39578
rect 2134 39520 2190 39584
rect 2976 39630 3110 39658
rect 3240 39704 3292 39710
rect 3240 39646 3292 39652
rect 3882 39658 3938 40000
rect 4802 39658 4858 40000
rect 5722 39658 5778 40000
rect 6550 39658 6606 40000
rect 7470 39658 7526 40000
rect 8390 39658 8446 40000
rect 9218 39658 9274 40000
rect 10138 39658 10194 40000
rect 2976 36310 3004 39630
rect 3054 39520 3110 39630
rect 2964 36304 3016 36310
rect 2964 36246 3016 36252
rect 3056 27940 3108 27946
rect 3056 27882 3108 27888
rect 2872 26240 2924 26246
rect 2872 26182 2924 26188
rect 2688 25900 2740 25906
rect 2688 25842 2740 25848
rect 2700 25362 2728 25842
rect 2884 25362 2912 26182
rect 2964 25968 3016 25974
rect 2964 25910 3016 25916
rect 2688 25356 2740 25362
rect 2688 25298 2740 25304
rect 2872 25356 2924 25362
rect 2872 25298 2924 25304
rect 2700 24954 2728 25298
rect 2884 24954 2912 25298
rect 2688 24948 2740 24954
rect 2688 24890 2740 24896
rect 2872 24948 2924 24954
rect 2872 24890 2924 24896
rect 2412 24064 2464 24070
rect 2412 24006 2464 24012
rect 2424 19174 2452 24006
rect 2884 23186 2912 24890
rect 2976 24274 3004 25910
rect 2964 24268 3016 24274
rect 2964 24210 3016 24216
rect 2976 23798 3004 24210
rect 2964 23792 3016 23798
rect 2964 23734 3016 23740
rect 2964 23588 3016 23594
rect 2964 23530 3016 23536
rect 2872 23180 2924 23186
rect 2872 23122 2924 23128
rect 2884 22778 2912 23122
rect 2872 22772 2924 22778
rect 2872 22714 2924 22720
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 2056 18426 2084 18770
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 110 12472 166 12481
rect 110 12407 166 12416
rect 124 12374 152 12407
rect 112 12368 164 12374
rect 112 12310 164 12316
rect 2424 11218 2452 19110
rect 2780 18896 2832 18902
rect 2780 18838 2832 18844
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2516 17610 2544 18158
rect 2608 17814 2636 18566
rect 2792 18358 2820 18838
rect 2976 18834 3004 23530
rect 2964 18828 3016 18834
rect 2964 18770 3016 18776
rect 2976 18358 3004 18770
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2964 18352 3016 18358
rect 2964 18294 3016 18300
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2596 17808 2648 17814
rect 2596 17750 2648 17756
rect 2504 17604 2556 17610
rect 2504 17546 2556 17552
rect 2700 14958 2728 18158
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2976 17202 3004 17682
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2700 14618 2728 14894
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2700 13870 2728 14554
rect 2976 14414 3004 15438
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2424 10810 2452 11154
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2424 9586 2452 10746
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 664 8560 716 8566
rect 664 8502 716 8508
rect 112 3936 164 3942
rect 112 3878 164 3884
rect 124 2553 152 3878
rect 110 2544 166 2553
rect 110 2479 166 2488
rect 386 82 442 480
rect 676 82 704 8502
rect 2318 6896 2374 6905
rect 2318 6831 2374 6840
rect 2504 6860 2556 6866
rect 2332 6322 2360 6831
rect 2504 6802 2556 6808
rect 2516 6458 2544 6802
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2424 5914 2452 6190
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2608 3754 2636 9930
rect 2700 9654 2728 13806
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 2976 11898 3004 12242
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2884 10810 2912 11154
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2964 9920 3016 9926
rect 3068 9908 3096 27882
rect 3252 26926 3280 39646
rect 3882 39630 4108 39658
rect 3882 39520 3938 39630
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 4080 32978 4108 39630
rect 4802 39630 4936 39658
rect 4802 39520 4858 39630
rect 4436 35624 4488 35630
rect 4436 35566 4488 35572
rect 4160 34536 4212 34542
rect 4160 34478 4212 34484
rect 4068 32972 4120 32978
rect 4068 32914 4120 32920
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3516 28008 3568 28014
rect 3516 27950 3568 27956
rect 3240 26920 3292 26926
rect 3240 26862 3292 26868
rect 3240 26784 3292 26790
rect 3240 26726 3292 26732
rect 3148 23656 3200 23662
rect 3146 23624 3148 23633
rect 3200 23624 3202 23633
rect 3146 23559 3202 23568
rect 3160 23526 3188 23559
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 3148 22976 3200 22982
rect 3148 22918 3200 22924
rect 3160 17270 3188 22918
rect 3148 17264 3200 17270
rect 3148 17206 3200 17212
rect 3252 13814 3280 26726
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3436 24070 3464 24550
rect 3424 24064 3476 24070
rect 3424 24006 3476 24012
rect 3332 23656 3384 23662
rect 3332 23598 3384 23604
rect 3344 22982 3372 23598
rect 3424 23588 3476 23594
rect 3528 23576 3556 27950
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 4172 27062 4200 34478
rect 4448 28218 4476 35566
rect 4528 29232 4580 29238
rect 4528 29174 4580 29180
rect 4436 28212 4488 28218
rect 4436 28154 4488 28160
rect 4448 28014 4476 28154
rect 4436 28008 4488 28014
rect 4436 27950 4488 27956
rect 4540 27538 4568 29174
rect 4908 28626 4936 39630
rect 5722 39630 5948 39658
rect 5722 39520 5778 39630
rect 5814 37224 5870 37233
rect 5814 37159 5870 37168
rect 5828 35222 5856 37159
rect 5816 35216 5868 35222
rect 5816 35158 5868 35164
rect 5816 35012 5868 35018
rect 5816 34954 5868 34960
rect 5828 34746 5856 34954
rect 5816 34740 5868 34746
rect 5816 34682 5868 34688
rect 5264 34060 5316 34066
rect 5264 34002 5316 34008
rect 5276 33318 5304 34002
rect 5264 33312 5316 33318
rect 5264 33254 5316 33260
rect 5276 32842 5304 33254
rect 5724 32972 5776 32978
rect 5724 32914 5776 32920
rect 5264 32836 5316 32842
rect 5264 32778 5316 32784
rect 5736 32570 5764 32914
rect 5724 32564 5776 32570
rect 5724 32506 5776 32512
rect 5540 31884 5592 31890
rect 5540 31826 5592 31832
rect 5552 31142 5580 31826
rect 5540 31136 5592 31142
rect 5540 31078 5592 31084
rect 5264 30728 5316 30734
rect 5264 30670 5316 30676
rect 5080 29300 5132 29306
rect 5080 29242 5132 29248
rect 4896 28620 4948 28626
rect 4896 28562 4948 28568
rect 4804 28416 4856 28422
rect 4804 28358 4856 28364
rect 4816 27674 4844 28358
rect 4908 28218 4936 28562
rect 4896 28212 4948 28218
rect 4896 28154 4948 28160
rect 4908 27946 4936 28154
rect 4896 27940 4948 27946
rect 4896 27882 4948 27888
rect 4804 27668 4856 27674
rect 4804 27610 4856 27616
rect 4528 27532 4580 27538
rect 4528 27474 4580 27480
rect 4540 27062 4568 27474
rect 4160 27056 4212 27062
rect 4160 26998 4212 27004
rect 4528 27056 4580 27062
rect 4528 26998 4580 27004
rect 4816 26994 4844 27610
rect 4804 26988 4856 26994
rect 4804 26930 4856 26936
rect 4620 26920 4672 26926
rect 4620 26862 4672 26868
rect 4632 26790 4660 26862
rect 4988 26852 5040 26858
rect 4988 26794 5040 26800
rect 4620 26784 4672 26790
rect 4620 26726 4672 26732
rect 4160 26512 4212 26518
rect 4160 26454 4212 26460
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3976 25832 4028 25838
rect 3976 25774 4028 25780
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3988 24818 4016 25774
rect 4172 25770 4200 26454
rect 4160 25764 4212 25770
rect 4160 25706 4212 25712
rect 4172 25498 4200 25706
rect 4160 25492 4212 25498
rect 4160 25434 4212 25440
rect 4344 25152 4396 25158
rect 4344 25094 4396 25100
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 4160 24676 4212 24682
rect 4160 24618 4212 24624
rect 4172 24274 4200 24618
rect 3976 24268 4028 24274
rect 3976 24210 4028 24216
rect 4160 24268 4212 24274
rect 4160 24210 4212 24216
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3988 23866 4016 24210
rect 4172 24070 4200 24210
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 3976 23860 4028 23866
rect 3976 23802 4028 23808
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 3476 23548 3556 23576
rect 3424 23530 3476 23536
rect 3516 23112 3568 23118
rect 3516 23054 3568 23060
rect 3332 22976 3384 22982
rect 3332 22918 3384 22924
rect 3528 22778 3556 23054
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 4080 22778 4108 23734
rect 4172 23662 4200 24006
rect 4356 23730 4384 25094
rect 4344 23724 4396 23730
rect 4344 23666 4396 23672
rect 4160 23656 4212 23662
rect 4160 23598 4212 23604
rect 4344 23588 4396 23594
rect 4344 23530 4396 23536
rect 4436 23588 4488 23594
rect 4436 23530 4488 23536
rect 4356 23322 4384 23530
rect 4344 23316 4396 23322
rect 4344 23258 4396 23264
rect 4356 22982 4384 23258
rect 4344 22976 4396 22982
rect 4344 22918 4396 22924
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 4080 22574 4108 22714
rect 4068 22568 4120 22574
rect 4068 22510 4120 22516
rect 4356 22234 4384 22918
rect 4344 22228 4396 22234
rect 4344 22170 4396 22176
rect 4158 21992 4214 22001
rect 4158 21927 4214 21936
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3424 21412 3476 21418
rect 3424 21354 3476 21360
rect 3332 19440 3384 19446
rect 3332 19382 3384 19388
rect 3344 18970 3372 19382
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3344 18222 3372 18702
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3160 13786 3280 13814
rect 3344 13814 3372 18022
rect 3436 16658 3464 21354
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 3804 21146 3832 21286
rect 3792 21140 3844 21146
rect 3792 21082 3844 21088
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3988 20602 4016 20878
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 3528 19394 3556 20538
rect 4068 20324 4120 20330
rect 4068 20266 4120 20272
rect 3976 19916 4028 19922
rect 3976 19858 4028 19864
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3988 19514 4016 19858
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 3974 19408 4030 19417
rect 3528 19366 3648 19394
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3528 18970 3556 19246
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3620 18612 3648 19366
rect 3974 19343 4030 19352
rect 3528 18584 3648 18612
rect 3528 18222 3556 18584
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3528 17882 3556 18158
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 3514 16960 3570 16969
rect 3514 16895 3570 16904
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3528 16250 3556 16895
rect 3896 16794 3924 17206
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3608 13864 3660 13870
rect 3344 13786 3464 13814
rect 3608 13806 3660 13812
rect 3160 13376 3188 13786
rect 3332 13388 3384 13394
rect 3160 13348 3332 13376
rect 3332 13330 3384 13336
rect 3344 12646 3372 13330
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10674 3188 11086
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3016 9880 3096 9908
rect 2964 9862 3016 9868
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2700 6934 2728 9590
rect 2976 9382 3004 9862
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2700 6458 2728 6870
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2872 4752 2924 4758
rect 2872 4694 2924 4700
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2424 3726 2636 3754
rect 2424 3194 2452 3726
rect 2700 3670 2728 4422
rect 2884 4078 2912 4694
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 1124 3188 1176 3194
rect 1124 3130 1176 3136
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 386 54 704 82
rect 1136 82 1164 3130
rect 2516 2582 2544 3470
rect 2608 3194 2636 3538
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2608 3097 2636 3130
rect 2594 3088 2650 3097
rect 2700 3058 2728 3606
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2594 3023 2650 3032
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2792 2922 2820 3334
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2504 2576 2556 2582
rect 2504 2518 2556 2524
rect 2792 2446 2820 2858
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 1214 82 1270 480
rect 1136 54 1270 82
rect 386 0 442 54
rect 1214 0 1270 54
rect 2134 82 2190 480
rect 2884 82 2912 4014
rect 2976 3194 3004 9318
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 3068 1306 3096 7958
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3160 3602 3188 6734
rect 3252 6458 3280 9522
rect 3344 7426 3372 12582
rect 3436 7562 3464 13786
rect 3620 13530 3648 13806
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3514 11792 3570 11801
rect 3514 11727 3570 11736
rect 3528 11694 3556 11727
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3528 9042 3556 11630
rect 3988 11393 4016 19343
rect 4080 17134 4108 20266
rect 4172 19854 4200 21927
rect 4356 21486 4384 22170
rect 4448 21554 4476 23530
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4436 21548 4488 21554
rect 4436 21490 4488 21496
rect 4344 21480 4396 21486
rect 4344 21422 4396 21428
rect 4356 21010 4384 21422
rect 4540 21146 4568 21966
rect 4528 21140 4580 21146
rect 4528 21082 4580 21088
rect 4344 21004 4396 21010
rect 4344 20946 4396 20952
rect 4344 20868 4396 20874
rect 4344 20810 4396 20816
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 4264 19417 4292 20198
rect 4250 19408 4306 19417
rect 4250 19343 4306 19352
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 4264 18970 4292 19246
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4264 18290 4292 18906
rect 4356 18426 4384 20810
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 4540 19922 4568 20402
rect 4528 19916 4580 19922
rect 4528 19858 4580 19864
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 4540 19174 4568 19314
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4172 16998 4200 17682
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4080 12714 4108 16730
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 4172 15366 4200 16526
rect 4264 16182 4292 16594
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 4264 15910 4292 16118
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4172 15026 4200 15302
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4172 12782 4200 14962
rect 4264 14278 4292 15846
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 4264 12918 4292 13330
rect 4252 12912 4304 12918
rect 4252 12854 4304 12860
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 3974 11384 4030 11393
rect 3974 11319 4030 11328
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 4080 10690 4108 12650
rect 4172 12442 4200 12718
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4172 11694 4200 12378
rect 4356 11778 4384 18158
rect 4540 16250 4568 19110
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4540 15978 4568 16186
rect 4528 15972 4580 15978
rect 4528 15914 4580 15920
rect 4540 15638 4568 15914
rect 4528 15632 4580 15638
rect 4528 15574 4580 15580
rect 4436 15088 4488 15094
rect 4436 15030 4488 15036
rect 4632 15042 4660 26726
rect 5000 26382 5028 26794
rect 4804 26376 4856 26382
rect 4804 26318 4856 26324
rect 4988 26376 5040 26382
rect 4988 26318 5040 26324
rect 4816 25702 4844 26318
rect 4804 25696 4856 25702
rect 4804 25638 4856 25644
rect 4816 24342 4844 25638
rect 4804 24336 4856 24342
rect 4804 24278 4856 24284
rect 4896 24132 4948 24138
rect 4896 24074 4948 24080
rect 4908 23526 4936 24074
rect 4896 23520 4948 23526
rect 4896 23462 4948 23468
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 4712 22704 4764 22710
rect 4712 22646 4764 22652
rect 4724 21078 4752 22646
rect 4816 22574 4844 22918
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 4816 21554 4844 22510
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4712 21072 4764 21078
rect 4712 21014 4764 21020
rect 4724 20602 4752 21014
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 4908 20448 4936 23462
rect 4988 23248 5040 23254
rect 4988 23190 5040 23196
rect 5000 22778 5028 23190
rect 4988 22772 5040 22778
rect 4988 22714 5040 22720
rect 4988 22500 5040 22506
rect 4988 22442 5040 22448
rect 5000 22166 5028 22442
rect 4988 22160 5040 22166
rect 4988 22102 5040 22108
rect 5000 21690 5028 22102
rect 4988 21684 5040 21690
rect 4988 21626 5040 21632
rect 4908 20420 5028 20448
rect 4804 20324 4856 20330
rect 4804 20266 4856 20272
rect 4896 20324 4948 20330
rect 4896 20266 4948 20272
rect 4816 20058 4844 20266
rect 4908 20058 4936 20266
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4908 19514 4936 19994
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4724 18426 4752 18770
rect 5000 18630 5028 20420
rect 5092 20262 5120 29242
rect 5276 29170 5304 30670
rect 5264 29164 5316 29170
rect 5264 29106 5316 29112
rect 5264 28416 5316 28422
rect 5264 28358 5316 28364
rect 5356 28416 5408 28422
rect 5356 28358 5408 28364
rect 5276 27946 5304 28358
rect 5368 28082 5396 28358
rect 5356 28076 5408 28082
rect 5356 28018 5408 28024
rect 5264 27940 5316 27946
rect 5264 27882 5316 27888
rect 5276 27674 5304 27882
rect 5264 27668 5316 27674
rect 5264 27610 5316 27616
rect 5276 26858 5304 27610
rect 5368 27606 5396 28018
rect 5356 27600 5408 27606
rect 5356 27542 5408 27548
rect 5264 26852 5316 26858
rect 5264 26794 5316 26800
rect 5276 26042 5304 26794
rect 5356 26308 5408 26314
rect 5356 26250 5408 26256
rect 5264 26036 5316 26042
rect 5264 25978 5316 25984
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 5276 24954 5304 25434
rect 5264 24948 5316 24954
rect 5264 24890 5316 24896
rect 5368 23118 5396 26250
rect 5552 26246 5580 31078
rect 5632 29504 5684 29510
rect 5632 29446 5684 29452
rect 5644 29034 5672 29446
rect 5920 29306 5948 39630
rect 6550 39630 6868 39658
rect 6550 39520 6606 39630
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6736 35148 6788 35154
rect 6736 35090 6788 35096
rect 6092 34468 6144 34474
rect 6092 34410 6144 34416
rect 6104 33658 6132 34410
rect 6748 34406 6776 35090
rect 6736 34400 6788 34406
rect 6736 34342 6788 34348
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6368 34128 6420 34134
rect 6368 34070 6420 34076
rect 6184 33924 6236 33930
rect 6184 33866 6236 33872
rect 6092 33652 6144 33658
rect 6092 33594 6144 33600
rect 6000 33312 6052 33318
rect 6000 33254 6052 33260
rect 5908 29300 5960 29306
rect 5908 29242 5960 29248
rect 5632 29028 5684 29034
rect 5632 28970 5684 28976
rect 5644 28150 5672 28970
rect 5632 28144 5684 28150
rect 5632 28086 5684 28092
rect 6012 28064 6040 33254
rect 6196 33114 6224 33866
rect 6380 33658 6408 34070
rect 6368 33652 6420 33658
rect 6368 33594 6420 33600
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6184 33108 6236 33114
rect 6184 33050 6236 33056
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6644 31884 6696 31890
rect 6644 31826 6696 31832
rect 6656 31142 6684 31826
rect 6644 31136 6696 31142
rect 6644 31078 6696 31084
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6656 30054 6684 31078
rect 6748 30802 6776 34342
rect 6840 32502 6868 39630
rect 7470 39630 7604 39658
rect 7470 39520 7526 39630
rect 7576 36242 7604 39630
rect 8036 39630 8446 39658
rect 7564 36236 7616 36242
rect 7564 36178 7616 36184
rect 7840 36236 7892 36242
rect 7840 36178 7892 36184
rect 7852 35766 7880 36178
rect 7840 35760 7892 35766
rect 7840 35702 7892 35708
rect 8036 35290 8064 39630
rect 8390 39520 8446 39630
rect 8864 39630 9274 39658
rect 8864 36378 8892 39630
rect 9218 39520 9274 39630
rect 9784 39630 10194 39658
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8852 36372 8904 36378
rect 8852 36314 8904 36320
rect 8392 36236 8444 36242
rect 8392 36178 8444 36184
rect 9680 36236 9732 36242
rect 9680 36178 9732 36184
rect 8116 36032 8168 36038
rect 8116 35974 8168 35980
rect 8208 36032 8260 36038
rect 8208 35974 8260 35980
rect 8128 35698 8156 35974
rect 8116 35692 8168 35698
rect 8116 35634 8168 35640
rect 8128 35290 8156 35634
rect 8220 35494 8248 35974
rect 8404 35698 8432 36178
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 9692 35698 9720 36178
rect 8392 35692 8444 35698
rect 8392 35634 8444 35640
rect 9680 35692 9732 35698
rect 9680 35634 9732 35640
rect 8208 35488 8260 35494
rect 8208 35430 8260 35436
rect 8024 35284 8076 35290
rect 8024 35226 8076 35232
rect 8116 35284 8168 35290
rect 8116 35226 8168 35232
rect 8220 35222 8248 35430
rect 8208 35216 8260 35222
rect 8208 35158 8260 35164
rect 7012 35148 7064 35154
rect 7012 35090 7064 35096
rect 7024 34406 7052 35090
rect 8116 35080 8168 35086
rect 8116 35022 8168 35028
rect 7656 34944 7708 34950
rect 7656 34886 7708 34892
rect 7668 34474 7696 34886
rect 7748 34672 7800 34678
rect 7748 34614 7800 34620
rect 7656 34468 7708 34474
rect 7656 34410 7708 34416
rect 7012 34400 7064 34406
rect 7012 34342 7064 34348
rect 7024 33318 7052 34342
rect 7564 33856 7616 33862
rect 7564 33798 7616 33804
rect 7576 33522 7604 33798
rect 7564 33516 7616 33522
rect 7564 33458 7616 33464
rect 7656 33380 7708 33386
rect 7656 33322 7708 33328
rect 7012 33312 7064 33318
rect 7012 33254 7064 33260
rect 7668 33114 7696 33322
rect 7104 33108 7156 33114
rect 7104 33050 7156 33056
rect 7656 33108 7708 33114
rect 7656 33050 7708 33056
rect 6828 32496 6880 32502
rect 6828 32438 6880 32444
rect 7116 32434 7144 33050
rect 7380 32904 7432 32910
rect 7380 32846 7432 32852
rect 7104 32428 7156 32434
rect 7104 32370 7156 32376
rect 6828 32360 6880 32366
rect 6828 32302 6880 32308
rect 6840 31958 6868 32302
rect 7288 32224 7340 32230
rect 7288 32166 7340 32172
rect 6828 31952 6880 31958
rect 6828 31894 6880 31900
rect 6920 31272 6972 31278
rect 6920 31214 6972 31220
rect 6736 30796 6788 30802
rect 6736 30738 6788 30744
rect 6932 30598 6960 31214
rect 7104 30728 7156 30734
rect 7104 30670 7156 30676
rect 6920 30592 6972 30598
rect 6920 30534 6972 30540
rect 6644 30048 6696 30054
rect 6644 29990 6696 29996
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6656 29714 6684 29990
rect 6644 29708 6696 29714
rect 6644 29650 6696 29656
rect 6656 28966 6684 29650
rect 6736 29640 6788 29646
rect 6736 29582 6788 29588
rect 6644 28960 6696 28966
rect 6644 28902 6696 28908
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6656 28626 6684 28902
rect 6184 28620 6236 28626
rect 6184 28562 6236 28568
rect 6644 28620 6696 28626
rect 6644 28562 6696 28568
rect 5828 28036 6040 28064
rect 5632 27600 5684 27606
rect 5632 27542 5684 27548
rect 5644 26586 5672 27542
rect 5724 27464 5776 27470
rect 5724 27406 5776 27412
rect 5736 27130 5764 27406
rect 5724 27124 5776 27130
rect 5724 27066 5776 27072
rect 5736 26586 5764 27066
rect 5828 27033 5856 28036
rect 5908 27940 5960 27946
rect 5908 27882 5960 27888
rect 5920 27402 5948 27882
rect 6000 27872 6052 27878
rect 6000 27814 6052 27820
rect 5908 27396 5960 27402
rect 5908 27338 5960 27344
rect 5814 27024 5870 27033
rect 5814 26959 5870 26968
rect 5632 26580 5684 26586
rect 5632 26522 5684 26528
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 5540 26240 5592 26246
rect 5540 26182 5592 26188
rect 5632 24744 5684 24750
rect 5632 24686 5684 24692
rect 5540 24132 5592 24138
rect 5540 24074 5592 24080
rect 5552 23662 5580 24074
rect 5644 24070 5672 24686
rect 5632 24064 5684 24070
rect 5632 24006 5684 24012
rect 5644 23662 5672 24006
rect 5540 23656 5592 23662
rect 5540 23598 5592 23604
rect 5632 23656 5684 23662
rect 5632 23598 5684 23604
rect 5828 23474 5856 26959
rect 5920 26314 5948 27338
rect 6012 26994 6040 27814
rect 6196 27334 6224 28562
rect 6656 28218 6684 28562
rect 6748 28422 6776 29582
rect 6828 28552 6880 28558
rect 6828 28494 6880 28500
rect 6736 28416 6788 28422
rect 6736 28358 6788 28364
rect 6644 28212 6696 28218
rect 6644 28154 6696 28160
rect 6840 28082 6868 28494
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6840 27674 6868 28018
rect 6828 27668 6880 27674
rect 6828 27610 6880 27616
rect 6276 27600 6328 27606
rect 6276 27542 6328 27548
rect 6184 27328 6236 27334
rect 6184 27270 6236 27276
rect 6288 27130 6316 27542
rect 6644 27328 6696 27334
rect 6644 27270 6696 27276
rect 6276 27124 6328 27130
rect 6276 27066 6328 27072
rect 6000 26988 6052 26994
rect 6000 26930 6052 26936
rect 6184 26920 6236 26926
rect 6184 26862 6236 26868
rect 6196 26518 6224 26862
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6184 26512 6236 26518
rect 6104 26472 6184 26500
rect 5908 26308 5960 26314
rect 5908 26250 5960 26256
rect 6104 25702 6132 26472
rect 6184 26454 6236 26460
rect 6460 26376 6512 26382
rect 6460 26318 6512 26324
rect 6472 26042 6500 26318
rect 6460 26036 6512 26042
rect 6460 25978 6512 25984
rect 6092 25696 6144 25702
rect 6092 25638 6144 25644
rect 6104 25498 6132 25638
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6092 25492 6144 25498
rect 6092 25434 6144 25440
rect 5908 25152 5960 25158
rect 5908 25094 5960 25100
rect 5920 24818 5948 25094
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 6656 24682 6684 27270
rect 6734 26888 6790 26897
rect 6734 26823 6790 26832
rect 6748 25906 6776 26823
rect 6932 26042 6960 30534
rect 7012 29232 7064 29238
rect 7012 29174 7064 29180
rect 6920 26036 6972 26042
rect 6920 25978 6972 25984
rect 6736 25900 6788 25906
rect 6736 25842 6788 25848
rect 6736 25424 6788 25430
rect 6736 25366 6788 25372
rect 6748 24954 6776 25366
rect 6736 24948 6788 24954
rect 6736 24890 6788 24896
rect 6644 24676 6696 24682
rect 6644 24618 6696 24624
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6092 24404 6144 24410
rect 6092 24346 6144 24352
rect 6000 24268 6052 24274
rect 6000 24210 6052 24216
rect 6012 23594 6040 24210
rect 5908 23588 5960 23594
rect 5908 23530 5960 23536
rect 6000 23588 6052 23594
rect 6000 23530 6052 23536
rect 5736 23446 5856 23474
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5460 22234 5488 22714
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5552 20466 5580 23054
rect 5632 21684 5684 21690
rect 5632 21626 5684 21632
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 5552 19990 5580 20402
rect 5644 19990 5672 21626
rect 5540 19984 5592 19990
rect 5540 19926 5592 19932
rect 5632 19984 5684 19990
rect 5632 19926 5684 19932
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5552 19310 5580 19790
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5632 19236 5684 19242
rect 5632 19178 5684 19184
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5172 18896 5224 18902
rect 5172 18838 5224 18844
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 4724 18086 4752 18362
rect 5000 18222 5028 18566
rect 4988 18216 5040 18222
rect 4988 18158 5040 18164
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4724 17134 4752 17478
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4724 16658 4752 17070
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 5000 16794 5028 17002
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4816 15570 4844 16526
rect 5000 16114 5028 16730
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 5092 15706 5120 15982
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4816 15162 4844 15506
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 5000 15094 5028 15574
rect 4988 15088 5040 15094
rect 4448 14890 4476 15030
rect 4632 15014 4844 15042
rect 4988 15030 5040 15036
rect 4436 14884 4488 14890
rect 4436 14826 4488 14832
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4436 14340 4488 14346
rect 4436 14282 4488 14288
rect 4448 13938 4476 14282
rect 4632 14074 4660 14350
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4724 13814 4752 14486
rect 4816 14396 4844 15014
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4908 14550 4936 14758
rect 5000 14550 5028 15030
rect 4896 14544 4948 14550
rect 4896 14486 4948 14492
rect 4988 14544 5040 14550
rect 4988 14486 5040 14492
rect 5092 14414 5120 15642
rect 5080 14408 5132 14414
rect 4816 14368 4936 14396
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4632 13786 4752 13814
rect 4632 13530 4660 13786
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4434 11792 4490 11801
rect 4356 11750 4434 11778
rect 4434 11727 4490 11736
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4172 11354 4200 11630
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4264 11150 4292 11562
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4172 10810 4200 10950
rect 4264 10810 4292 11086
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4080 10662 4200 10690
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3988 9722 4016 9998
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 3974 9616 4030 9625
rect 4080 9602 4108 10406
rect 4030 9574 4108 9602
rect 3974 9551 4030 9560
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3988 8294 4016 9551
rect 4172 9500 4200 10662
rect 4356 10266 4384 11562
rect 4540 11354 4568 12718
rect 4724 12714 4752 13126
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4724 12442 4752 12650
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4448 10266 4476 10542
rect 4540 10538 4568 11290
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4540 9926 4568 10474
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4080 9472 4200 9500
rect 4080 9110 4108 9472
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3436 7534 3556 7562
rect 3344 7398 3464 7426
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3252 6254 3280 6394
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3332 5296 3384 5302
rect 3332 5238 3384 5244
rect 3240 4208 3292 4214
rect 3240 4150 3292 4156
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3252 2582 3280 4150
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 3344 2310 3372 5238
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 2134 54 2912 82
rect 2976 1278 3096 1306
rect 2976 82 3004 1278
rect 3054 82 3110 480
rect 3436 134 3464 7398
rect 3528 4690 3556 7534
rect 3988 7342 4016 8026
rect 4080 7410 4108 9046
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4172 7970 4200 8230
rect 4264 8090 4292 8366
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4172 7942 4292 7970
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3988 6866 4016 7278
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3988 6730 4016 6802
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3988 6254 4016 6666
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3988 5914 4016 6190
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3988 5166 4016 5850
rect 4080 5778 4108 7346
rect 4172 6322 4200 7754
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4080 5370 4108 5714
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3988 4826 4016 5102
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3528 3942 3556 4626
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3988 4010 4016 4490
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3528 3641 3556 3878
rect 3988 3738 4016 3946
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3514 3632 3570 3641
rect 3514 3567 3570 3576
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 2650 3556 3334
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 4172 3058 4200 6122
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4172 2650 4200 2994
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 2976 54 3110 82
rect 3424 128 3476 134
rect 3424 70 3476 76
rect 3882 82 3938 480
rect 4264 82 4292 7942
rect 4356 7002 4384 8298
rect 4448 8294 4476 8978
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4448 7206 4476 7822
rect 4540 7342 4568 9862
rect 4724 9722 4752 10066
rect 4712 9716 4764 9722
rect 4632 9676 4712 9704
rect 4632 8566 4660 9676
rect 4712 9658 4764 9664
rect 4816 9674 4844 14214
rect 4908 13297 4936 14368
rect 5080 14350 5132 14356
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 4894 13288 4950 13297
rect 4894 13223 4950 13232
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4908 12850 4936 13126
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 5000 12782 5028 13330
rect 5092 12986 5120 13806
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5184 12918 5212 18838
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5276 17338 5304 17682
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5276 13802 5304 14214
rect 5460 13814 5488 18294
rect 5552 18222 5580 18906
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5552 17746 5580 18158
rect 5644 17882 5672 19178
rect 5736 18902 5764 23446
rect 5920 23322 5948 23530
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 5908 22092 5960 22098
rect 5908 22034 5960 22040
rect 5920 21690 5948 22034
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 5920 21078 5948 21626
rect 5908 21072 5960 21078
rect 5908 21014 5960 21020
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 5908 19984 5960 19990
rect 5908 19926 5960 19932
rect 5920 19174 5948 19926
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5920 18902 5948 19110
rect 5724 18896 5776 18902
rect 5724 18838 5776 18844
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5736 18154 5764 18702
rect 5920 18426 5948 18838
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5816 18216 5868 18222
rect 5816 18158 5868 18164
rect 5724 18148 5776 18154
rect 5724 18090 5776 18096
rect 5736 17882 5764 18090
rect 5632 17876 5684 17882
rect 5632 17818 5684 17824
rect 5724 17876 5776 17882
rect 5724 17818 5776 17824
rect 5828 17814 5856 18158
rect 5816 17808 5868 17814
rect 5816 17750 5868 17756
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5552 17338 5580 17682
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5552 15638 5580 15846
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5552 14890 5580 15302
rect 5540 14884 5592 14890
rect 5540 14826 5592 14832
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 5356 13796 5408 13802
rect 5460 13786 5580 13814
rect 5356 13738 5408 13744
rect 5276 13462 5304 13738
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5262 13288 5318 13297
rect 5262 13223 5318 13232
rect 5172 12912 5224 12918
rect 5172 12854 5224 12860
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 5080 12368 5132 12374
rect 5080 12310 5132 12316
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 5000 11014 5028 12174
rect 5092 11898 5120 12310
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5092 11558 5120 11834
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 11354 5120 11494
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 4816 9646 4936 9674
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4724 8430 4752 8978
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4356 6322 4384 6938
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4344 5772 4396 5778
rect 4448 5760 4476 7142
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 6458 4568 6734
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4396 5732 4476 5760
rect 4344 5714 4396 5720
rect 4356 4826 4384 5714
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4632 4049 4660 8298
rect 4816 8090 4844 8910
rect 4908 8634 4936 9646
rect 5080 9512 5132 9518
rect 5078 9480 5080 9489
rect 5132 9480 5134 9489
rect 5078 9415 5134 9424
rect 5092 9382 5120 9415
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5276 8362 5304 13223
rect 5368 12714 5396 13738
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 10198 5396 10406
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5368 9450 5396 10134
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5368 9178 5396 9386
rect 5460 9382 5488 9522
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 8430 5396 8774
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4816 7410 4844 8026
rect 5368 7954 5396 8366
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4896 7268 4948 7274
rect 4896 7210 4948 7216
rect 4908 6866 4936 7210
rect 5000 6934 5028 7890
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5460 6934 5488 7210
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4724 4622 4752 5034
rect 4816 4758 4844 6666
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4908 5574 4936 6054
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4908 4758 4936 5510
rect 5000 5234 5028 6870
rect 5460 6186 5488 6870
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5368 5302 5396 5714
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5356 5296 5408 5302
rect 5356 5238 5408 5244
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4724 4282 4752 4558
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4908 4078 4936 4694
rect 5276 4690 5304 5170
rect 5460 4758 5488 5646
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 4896 4072 4948 4078
rect 4618 4040 4674 4049
rect 4896 4014 4948 4020
rect 4618 3975 4674 3984
rect 4632 3097 4660 3975
rect 4908 3670 4936 4014
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5368 3738 5396 3946
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 4618 3088 4674 3097
rect 4618 3023 4674 3032
rect 4908 2922 4936 3606
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5368 3194 5396 3538
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5552 3126 5580 13786
rect 5644 12850 5672 15302
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 5816 13728 5868 13734
rect 5920 13716 5948 14554
rect 5868 13688 5948 13716
rect 5816 13670 5868 13676
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5644 12238 5672 12786
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5644 10062 5672 12174
rect 5828 11626 5856 13670
rect 6012 13274 6040 20402
rect 5920 13246 6040 13274
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5828 9654 5856 11562
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5644 5370 5672 7142
rect 5920 6730 5948 13246
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 6012 12714 6040 13126
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 6012 12442 6040 12650
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 6104 9722 6132 24346
rect 6748 23798 6776 24890
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 6736 23792 6788 23798
rect 6736 23734 6788 23740
rect 6840 23730 6868 24006
rect 6828 23724 6880 23730
rect 6828 23666 6880 23672
rect 6184 23656 6236 23662
rect 6184 23598 6236 23604
rect 6196 22166 6224 23598
rect 6736 23588 6788 23594
rect 6736 23530 6788 23536
rect 6748 23497 6776 23530
rect 6734 23488 6790 23497
rect 6289 23420 6585 23440
rect 6734 23423 6790 23432
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6184 22160 6236 22166
rect 6184 22102 6236 22108
rect 6196 21146 6224 22102
rect 6840 22030 6868 23666
rect 6920 23588 6972 23594
rect 6920 23530 6972 23536
rect 6932 23254 6960 23530
rect 7024 23474 7052 29174
rect 7116 29170 7144 30670
rect 7196 29640 7248 29646
rect 7196 29582 7248 29588
rect 7208 29170 7236 29582
rect 7104 29164 7156 29170
rect 7104 29106 7156 29112
rect 7196 29164 7248 29170
rect 7196 29106 7248 29112
rect 7208 28762 7236 29106
rect 7300 29102 7328 32166
rect 7392 31686 7420 32846
rect 7472 32564 7524 32570
rect 7472 32506 7524 32512
rect 7380 31680 7432 31686
rect 7380 31622 7432 31628
rect 7392 31346 7420 31622
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7484 30376 7512 32506
rect 7656 31884 7708 31890
rect 7656 31826 7708 31832
rect 7668 30938 7696 31826
rect 7656 30932 7708 30938
rect 7656 30874 7708 30880
rect 7392 30348 7512 30376
rect 7288 29096 7340 29102
rect 7288 29038 7340 29044
rect 7196 28756 7248 28762
rect 7196 28698 7248 28704
rect 7104 26988 7156 26994
rect 7104 26930 7156 26936
rect 7116 26586 7144 26930
rect 7104 26580 7156 26586
rect 7104 26522 7156 26528
rect 7196 26240 7248 26246
rect 7196 26182 7248 26188
rect 7208 24070 7236 26182
rect 7288 25152 7340 25158
rect 7288 25094 7340 25100
rect 7300 24682 7328 25094
rect 7288 24676 7340 24682
rect 7288 24618 7340 24624
rect 7288 24336 7340 24342
rect 7288 24278 7340 24284
rect 7196 24064 7248 24070
rect 7196 24006 7248 24012
rect 7024 23446 7144 23474
rect 6920 23248 6972 23254
rect 6920 23190 6972 23196
rect 6932 22778 6960 23190
rect 7012 22976 7064 22982
rect 7012 22918 7064 22924
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 7024 22710 7052 22918
rect 7012 22704 7064 22710
rect 7012 22646 7064 22652
rect 7024 22506 7052 22646
rect 7012 22500 7064 22506
rect 7012 22442 7064 22448
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6932 21622 6960 21966
rect 6920 21616 6972 21622
rect 6920 21558 6972 21564
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6184 21140 6236 21146
rect 6184 21082 6236 21088
rect 6196 18970 6224 21082
rect 6644 21072 6696 21078
rect 6644 21014 6696 21020
rect 6276 20936 6328 20942
rect 6276 20878 6328 20884
rect 6288 20602 6316 20878
rect 6276 20596 6328 20602
rect 6276 20538 6328 20544
rect 6656 20262 6684 21014
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6748 20330 6776 20742
rect 6736 20324 6788 20330
rect 7012 20324 7064 20330
rect 6736 20266 6788 20272
rect 6932 20284 7012 20312
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6656 19990 6684 20198
rect 6644 19984 6696 19990
rect 6644 19926 6696 19932
rect 6748 19446 6776 20266
rect 6932 19718 6960 20284
rect 7012 20266 7064 20272
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 6656 18358 6684 19110
rect 6932 18902 6960 19654
rect 6920 18896 6972 18902
rect 6920 18838 6972 18844
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6656 17882 6684 18294
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6748 17814 6776 18634
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6840 18222 6868 18566
rect 7116 18290 7144 23446
rect 7300 23322 7328 24278
rect 7392 23769 7420 30348
rect 7472 30184 7524 30190
rect 7472 30126 7524 30132
rect 7484 29850 7512 30126
rect 7564 30048 7616 30054
rect 7564 29990 7616 29996
rect 7472 29844 7524 29850
rect 7472 29786 7524 29792
rect 7484 28082 7512 29786
rect 7576 28626 7604 29990
rect 7564 28620 7616 28626
rect 7564 28562 7616 28568
rect 7576 28218 7604 28562
rect 7564 28212 7616 28218
rect 7564 28154 7616 28160
rect 7472 28076 7524 28082
rect 7472 28018 7524 28024
rect 7472 27396 7524 27402
rect 7472 27338 7524 27344
rect 7484 27062 7512 27338
rect 7472 27056 7524 27062
rect 7472 26998 7524 27004
rect 7378 23760 7434 23769
rect 7378 23695 7434 23704
rect 7288 23316 7340 23322
rect 7288 23258 7340 23264
rect 7196 23112 7248 23118
rect 7196 23054 7248 23060
rect 7208 22642 7236 23054
rect 7484 22710 7512 26998
rect 7656 26240 7708 26246
rect 7656 26182 7708 26188
rect 7668 25838 7696 26182
rect 7656 25832 7708 25838
rect 7656 25774 7708 25780
rect 7668 24682 7696 25774
rect 7656 24676 7708 24682
rect 7656 24618 7708 24624
rect 7668 24138 7696 24618
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 7668 23798 7696 24074
rect 7656 23792 7708 23798
rect 7656 23734 7708 23740
rect 7760 23474 7788 34614
rect 8128 34474 8156 35022
rect 7932 34468 7984 34474
rect 7932 34410 7984 34416
rect 8116 34468 8168 34474
rect 8116 34410 8168 34416
rect 7944 34134 7972 34410
rect 8128 34202 8156 34410
rect 8220 34406 8248 35158
rect 8300 35080 8352 35086
rect 8300 35022 8352 35028
rect 8312 34610 8340 35022
rect 8300 34604 8352 34610
rect 8300 34546 8352 34552
rect 8208 34400 8260 34406
rect 8208 34342 8260 34348
rect 8116 34196 8168 34202
rect 8116 34138 8168 34144
rect 7932 34128 7984 34134
rect 7932 34070 7984 34076
rect 7840 33992 7892 33998
rect 7840 33934 7892 33940
rect 7852 33046 7880 33934
rect 7944 33114 7972 34070
rect 8312 33522 8340 34546
rect 8024 33516 8076 33522
rect 8024 33458 8076 33464
rect 8300 33516 8352 33522
rect 8300 33458 8352 33464
rect 7932 33108 7984 33114
rect 7932 33050 7984 33056
rect 7840 33040 7892 33046
rect 7840 32982 7892 32988
rect 7944 32570 7972 33050
rect 7932 32564 7984 32570
rect 7932 32506 7984 32512
rect 7840 32496 7892 32502
rect 7840 32438 7892 32444
rect 7852 28370 7880 32438
rect 8036 30938 8064 33458
rect 8208 33312 8260 33318
rect 8208 33254 8260 33260
rect 8116 31884 8168 31890
rect 8116 31826 8168 31832
rect 8128 31142 8156 31826
rect 8116 31136 8168 31142
rect 8116 31078 8168 31084
rect 8024 30932 8076 30938
rect 8024 30874 8076 30880
rect 8036 29850 8064 30874
rect 8024 29844 8076 29850
rect 8024 29786 8076 29792
rect 8024 29708 8076 29714
rect 8024 29650 8076 29656
rect 7932 29096 7984 29102
rect 7932 29038 7984 29044
rect 7944 28762 7972 29038
rect 7932 28756 7984 28762
rect 7932 28698 7984 28704
rect 8036 28490 8064 29650
rect 8116 29300 8168 29306
rect 8116 29242 8168 29248
rect 8024 28484 8076 28490
rect 8024 28426 8076 28432
rect 7852 28342 8064 28370
rect 7840 27464 7892 27470
rect 7840 27406 7892 27412
rect 7852 27130 7880 27406
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 7840 26444 7892 26450
rect 7840 26386 7892 26392
rect 7852 25974 7880 26386
rect 7840 25968 7892 25974
rect 7840 25910 7892 25916
rect 7576 23446 7788 23474
rect 7472 22704 7524 22710
rect 7472 22646 7524 22652
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 7196 22500 7248 22506
rect 7196 22442 7248 22448
rect 7208 18834 7236 22442
rect 7484 22234 7512 22646
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7472 21072 7524 21078
rect 7472 21014 7524 21020
rect 7484 20534 7512 21014
rect 7576 21010 7604 23446
rect 7852 23254 7880 25910
rect 7932 24200 7984 24206
rect 7932 24142 7984 24148
rect 7944 23322 7972 24142
rect 7932 23316 7984 23322
rect 7932 23258 7984 23264
rect 7840 23248 7892 23254
rect 7840 23190 7892 23196
rect 7564 21004 7616 21010
rect 7564 20946 7616 20952
rect 7840 21004 7892 21010
rect 7840 20946 7892 20952
rect 7748 20868 7800 20874
rect 7748 20810 7800 20816
rect 7472 20528 7524 20534
rect 7472 20470 7524 20476
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7392 19378 7420 19654
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7104 18284 7156 18290
rect 7104 18226 7156 18232
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 6196 14929 6224 17070
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6748 16794 6776 17750
rect 7392 17678 7420 18702
rect 7484 17814 7512 20470
rect 7656 19236 7708 19242
rect 7656 19178 7708 19184
rect 7472 17808 7524 17814
rect 7472 17750 7524 17756
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 6828 17604 6880 17610
rect 6828 17546 6880 17552
rect 6840 16794 6868 17546
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 7208 16658 7236 17070
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7576 16658 7604 17002
rect 7668 16658 7696 19178
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 6656 16250 6684 16594
rect 7208 16522 7236 16594
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 7196 15632 7248 15638
rect 7196 15574 7248 15580
rect 6564 15162 6592 15574
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 7208 15026 7236 15574
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 6182 14920 6238 14929
rect 6182 14855 6238 14864
rect 6920 14884 6972 14890
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6196 9194 6224 14855
rect 6920 14826 6972 14832
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6748 14550 6776 14758
rect 6932 14618 6960 14826
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6380 14074 6408 14350
rect 7116 14074 7144 14486
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7116 13802 7144 14010
rect 7300 13938 7328 15846
rect 7392 15366 7420 15982
rect 7576 15706 7604 16594
rect 7668 16250 7696 16594
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7668 15502 7696 16186
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7392 14346 7420 15302
rect 7668 15162 7696 15438
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7760 15042 7788 20810
rect 7852 20466 7880 20946
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7840 19984 7892 19990
rect 7840 19926 7892 19932
rect 7852 19514 7880 19926
rect 7944 19786 7972 23258
rect 8036 20874 8064 28342
rect 8128 26926 8156 29242
rect 8220 27538 8248 33254
rect 8300 32904 8352 32910
rect 8300 32846 8352 32852
rect 8312 32570 8340 32846
rect 8300 32564 8352 32570
rect 8300 32506 8352 32512
rect 8300 30864 8352 30870
rect 8300 30806 8352 30812
rect 8312 30054 8340 30806
rect 8300 30048 8352 30054
rect 8300 29990 8352 29996
rect 8312 29306 8340 29990
rect 8300 29300 8352 29306
rect 8300 29242 8352 29248
rect 8404 29238 8432 35634
rect 8484 35556 8536 35562
rect 8484 35498 8536 35504
rect 8496 34134 8524 35498
rect 9692 35494 9720 35634
rect 9680 35488 9732 35494
rect 9680 35430 9732 35436
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 9784 34746 9812 39630
rect 10138 39520 10194 39630
rect 11058 39658 11114 40000
rect 11886 39658 11942 40000
rect 12806 39658 12862 40000
rect 13726 39658 13782 40000
rect 11058 39630 11376 39658
rect 11058 39520 11114 39630
rect 9956 36576 10008 36582
rect 9956 36518 10008 36524
rect 9968 35290 9996 36518
rect 10324 36032 10376 36038
rect 10324 35974 10376 35980
rect 10336 35698 10364 35974
rect 11244 35760 11296 35766
rect 11244 35702 11296 35708
rect 10324 35692 10376 35698
rect 10324 35634 10376 35640
rect 10416 35556 10468 35562
rect 10416 35498 10468 35504
rect 10968 35556 11020 35562
rect 10968 35498 11020 35504
rect 9956 35284 10008 35290
rect 9956 35226 10008 35232
rect 9772 34740 9824 34746
rect 9772 34682 9824 34688
rect 9968 34610 9996 35226
rect 9956 34604 10008 34610
rect 9956 34546 10008 34552
rect 9496 34400 9548 34406
rect 9496 34342 9548 34348
rect 10232 34400 10284 34406
rect 10232 34342 10284 34348
rect 8484 34128 8536 34134
rect 8484 34070 8536 34076
rect 8496 33930 8524 34070
rect 8484 33924 8536 33930
rect 8484 33866 8536 33872
rect 8496 33134 8524 33866
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 9312 33448 9364 33454
rect 9312 33390 9364 33396
rect 8496 33106 8616 33134
rect 8482 31920 8538 31929
rect 8482 31855 8538 31864
rect 8496 30394 8524 31855
rect 8588 30938 8616 33106
rect 9324 32774 9352 33390
rect 8760 32768 8812 32774
rect 8760 32710 8812 32716
rect 9312 32768 9364 32774
rect 9312 32710 9364 32716
rect 8772 32434 8800 32710
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8760 32428 8812 32434
rect 8760 32370 8812 32376
rect 8772 31958 8800 32370
rect 8760 31952 8812 31958
rect 8760 31894 8812 31900
rect 8668 31680 8720 31686
rect 8668 31622 8720 31628
rect 8680 31278 8708 31622
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 9324 31346 9352 32710
rect 9508 32570 9536 34342
rect 9956 34196 10008 34202
rect 9956 34138 10008 34144
rect 9772 33992 9824 33998
rect 9772 33934 9824 33940
rect 9784 33522 9812 33934
rect 9772 33516 9824 33522
rect 9772 33458 9824 33464
rect 9588 33312 9640 33318
rect 9588 33254 9640 33260
rect 9496 32564 9548 32570
rect 9496 32506 9548 32512
rect 9600 32230 9628 33254
rect 9588 32224 9640 32230
rect 9588 32166 9640 32172
rect 9784 32026 9812 33458
rect 9968 33386 9996 34138
rect 10244 33658 10272 34342
rect 10232 33652 10284 33658
rect 10232 33594 10284 33600
rect 10428 33590 10456 35498
rect 10876 35488 10928 35494
rect 10876 35430 10928 35436
rect 10600 35216 10652 35222
rect 10600 35158 10652 35164
rect 10508 35080 10560 35086
rect 10508 35022 10560 35028
rect 10520 33862 10548 35022
rect 10612 34406 10640 35158
rect 10692 34468 10744 34474
rect 10692 34410 10744 34416
rect 10600 34400 10652 34406
rect 10600 34342 10652 34348
rect 10508 33856 10560 33862
rect 10508 33798 10560 33804
rect 10416 33584 10468 33590
rect 10416 33526 10468 33532
rect 9956 33380 10008 33386
rect 9956 33322 10008 33328
rect 9968 33114 9996 33322
rect 10428 33114 10456 33526
rect 9956 33108 10008 33114
rect 9956 33050 10008 33056
rect 10416 33108 10468 33114
rect 10416 33050 10468 33056
rect 9968 32985 9996 33050
rect 10416 32904 10468 32910
rect 10416 32846 10468 32852
rect 10324 32360 10376 32366
rect 10324 32302 10376 32308
rect 10232 32292 10284 32298
rect 10232 32234 10284 32240
rect 9772 32020 9824 32026
rect 9772 31962 9824 31968
rect 10244 31890 10272 32234
rect 9956 31884 10008 31890
rect 9956 31826 10008 31832
rect 10232 31884 10284 31890
rect 10232 31826 10284 31832
rect 9968 31414 9996 31826
rect 10244 31482 10272 31826
rect 10336 31754 10364 32302
rect 10428 32230 10456 32846
rect 10416 32224 10468 32230
rect 10416 32166 10468 32172
rect 10324 31748 10376 31754
rect 10324 31690 10376 31696
rect 10232 31476 10284 31482
rect 10232 31418 10284 31424
rect 9956 31408 10008 31414
rect 9956 31350 10008 31356
rect 9312 31340 9364 31346
rect 9312 31282 9364 31288
rect 8668 31272 8720 31278
rect 8668 31214 8720 31220
rect 8668 31136 8720 31142
rect 8668 31078 8720 31084
rect 8576 30932 8628 30938
rect 8576 30874 8628 30880
rect 8484 30388 8536 30394
rect 8484 30330 8536 30336
rect 8680 29714 8708 31078
rect 9312 30864 9364 30870
rect 9312 30806 9364 30812
rect 10230 30832 10286 30841
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 9324 30054 9352 30806
rect 10230 30767 10286 30776
rect 9956 30184 10008 30190
rect 9956 30126 10008 30132
rect 9312 30048 9364 30054
rect 9312 29990 9364 29996
rect 8668 29708 8720 29714
rect 8668 29650 8720 29656
rect 8680 29306 8708 29650
rect 8852 29640 8904 29646
rect 8852 29582 8904 29588
rect 8668 29300 8720 29306
rect 8668 29242 8720 29248
rect 8392 29232 8444 29238
rect 8392 29174 8444 29180
rect 8300 29096 8352 29102
rect 8300 29038 8352 29044
rect 8312 28150 8340 29038
rect 8680 28694 8708 29242
rect 8864 29170 8892 29582
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8852 29164 8904 29170
rect 8852 29106 8904 29112
rect 9324 28762 9352 29990
rect 9968 29510 9996 30126
rect 10244 30054 10272 30767
rect 10232 30048 10284 30054
rect 10232 29990 10284 29996
rect 10244 29782 10272 29990
rect 10232 29776 10284 29782
rect 10232 29718 10284 29724
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 9968 28762 9996 29446
rect 10244 29306 10272 29718
rect 10600 29640 10652 29646
rect 10600 29582 10652 29588
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 10612 28966 10640 29582
rect 10600 28960 10652 28966
rect 10704 28948 10732 34410
rect 10784 33380 10836 33386
rect 10784 33322 10836 33328
rect 10796 32842 10824 33322
rect 10784 32836 10836 32842
rect 10784 32778 10836 32784
rect 10704 28920 10824 28948
rect 10600 28902 10652 28908
rect 9312 28756 9364 28762
rect 9312 28698 9364 28704
rect 9956 28756 10008 28762
rect 9956 28698 10008 28704
rect 8668 28688 8720 28694
rect 8668 28630 8720 28636
rect 8392 28484 8444 28490
rect 8392 28426 8444 28432
rect 8300 28144 8352 28150
rect 8300 28086 8352 28092
rect 8208 27532 8260 27538
rect 8208 27474 8260 27480
rect 8116 26920 8168 26926
rect 8116 26862 8168 26868
rect 8312 26568 8340 28086
rect 8404 27334 8432 28426
rect 8680 28218 8708 28630
rect 9680 28620 9732 28626
rect 9680 28562 9732 28568
rect 9588 28416 9640 28422
rect 9588 28358 9640 28364
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8668 28212 8720 28218
rect 8668 28154 8720 28160
rect 9600 28014 9628 28358
rect 9692 28082 9720 28562
rect 10612 28082 10640 28902
rect 9680 28076 9732 28082
rect 9680 28018 9732 28024
rect 10600 28076 10652 28082
rect 10600 28018 10652 28024
rect 9588 28008 9640 28014
rect 9588 27950 9640 27956
rect 8576 27940 8628 27946
rect 8576 27882 8628 27888
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8220 26540 8340 26568
rect 8220 25974 8248 26540
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 8312 26042 8340 26386
rect 8392 26376 8444 26382
rect 8392 26318 8444 26324
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 8208 25968 8260 25974
rect 8208 25910 8260 25916
rect 8220 25770 8248 25910
rect 8208 25764 8260 25770
rect 8208 25706 8260 25712
rect 8220 25430 8248 25706
rect 8208 25424 8260 25430
rect 8208 25366 8260 25372
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 8128 23186 8156 24550
rect 8208 24132 8260 24138
rect 8208 24074 8260 24080
rect 8220 23866 8248 24074
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8206 23760 8262 23769
rect 8206 23695 8262 23704
rect 8116 23180 8168 23186
rect 8116 23122 8168 23128
rect 8128 22642 8156 23122
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 8024 20868 8076 20874
rect 8024 20810 8076 20816
rect 7932 19780 7984 19786
rect 7932 19722 7984 19728
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7944 19378 7972 19722
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 7944 18698 7972 19314
rect 8024 18896 8076 18902
rect 8024 18838 8076 18844
rect 7932 18692 7984 18698
rect 7932 18634 7984 18640
rect 8036 18426 8064 18838
rect 8220 18612 8248 23695
rect 8312 22710 8340 25978
rect 8404 25906 8432 26318
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 8404 25498 8432 25842
rect 8392 25492 8444 25498
rect 8392 25434 8444 25440
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8496 24954 8524 25230
rect 8484 24948 8536 24954
rect 8484 24890 8536 24896
rect 8588 24834 8616 27882
rect 8760 27532 8812 27538
rect 8760 27474 8812 27480
rect 8772 26790 8800 27474
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 8852 27328 8904 27334
rect 8852 27270 8904 27276
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 8496 24806 8616 24834
rect 8392 23860 8444 23866
rect 8392 23802 8444 23808
rect 8300 22704 8352 22710
rect 8300 22646 8352 22652
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8312 21146 8340 21286
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 8312 20398 8340 21082
rect 8404 20942 8432 23802
rect 8496 23474 8524 24806
rect 8772 24410 8800 26726
rect 8864 25498 8892 27270
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 9416 26314 9444 27406
rect 9600 27334 9628 27950
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 9496 26852 9548 26858
rect 9496 26794 9548 26800
rect 9404 26308 9456 26314
rect 9404 26250 9456 26256
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 9312 25968 9364 25974
rect 9312 25910 9364 25916
rect 8852 25492 8904 25498
rect 8852 25434 8904 25440
rect 8864 24818 8892 25434
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 8852 24812 8904 24818
rect 8852 24754 8904 24760
rect 9324 24682 9352 25910
rect 9312 24676 9364 24682
rect 9312 24618 9364 24624
rect 8760 24404 8812 24410
rect 8760 24346 8812 24352
rect 8576 24268 8628 24274
rect 8576 24210 8628 24216
rect 8588 23866 8616 24210
rect 9416 24138 9444 26250
rect 9508 26246 9536 26794
rect 9496 26240 9548 26246
rect 9496 26182 9548 26188
rect 9508 25226 9536 26182
rect 9496 25220 9548 25226
rect 9496 25162 9548 25168
rect 9404 24132 9456 24138
rect 9404 24074 9456 24080
rect 9600 24070 9628 27270
rect 9692 24410 9720 28018
rect 9864 27600 9916 27606
rect 9864 27542 9916 27548
rect 9876 26994 9904 27542
rect 9864 26988 9916 26994
rect 9864 26930 9916 26936
rect 9772 26852 9824 26858
rect 9772 26794 9824 26800
rect 9784 25974 9812 26794
rect 9876 26518 9904 26930
rect 10048 26580 10100 26586
rect 10048 26522 10100 26528
rect 9864 26512 9916 26518
rect 9864 26454 9916 26460
rect 9876 26042 9904 26454
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 9772 25968 9824 25974
rect 9772 25910 9824 25916
rect 9864 25832 9916 25838
rect 9864 25774 9916 25780
rect 9876 25362 9904 25774
rect 9968 25498 9996 26318
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 10060 25362 10088 26522
rect 10692 26240 10744 26246
rect 10692 26182 10744 26188
rect 10704 25838 10732 26182
rect 10692 25832 10744 25838
rect 10692 25774 10744 25780
rect 10416 25764 10468 25770
rect 10416 25706 10468 25712
rect 10428 25498 10456 25706
rect 10416 25492 10468 25498
rect 10416 25434 10468 25440
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 10048 25356 10100 25362
rect 10048 25298 10100 25304
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 8852 24064 8904 24070
rect 8852 24006 8904 24012
rect 9588 24064 9640 24070
rect 9588 24006 9640 24012
rect 8576 23860 8628 23866
rect 8576 23802 8628 23808
rect 8864 23730 8892 24006
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 8668 23724 8720 23730
rect 8668 23666 8720 23672
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 8496 23446 8616 23474
rect 8484 22976 8536 22982
rect 8484 22918 8536 22924
rect 8496 22574 8524 22918
rect 8484 22568 8536 22574
rect 8484 22510 8536 22516
rect 8484 22092 8536 22098
rect 8484 22034 8536 22040
rect 8496 21622 8524 22034
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8312 18970 8340 19790
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8220 18584 8432 18612
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 7576 15014 7788 15042
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 7116 13530 7144 13738
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6840 12238 6868 13262
rect 7116 12986 7144 13466
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7116 12646 7144 12922
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6656 11218 6684 12038
rect 6840 11898 6868 12174
rect 7024 11898 7052 12310
rect 7116 11898 7144 12582
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7116 11626 7144 11834
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 7116 11286 7144 11562
rect 7104 11280 7156 11286
rect 6734 11248 6790 11257
rect 6644 11212 6696 11218
rect 7104 11222 7156 11228
rect 6734 11183 6790 11192
rect 6644 11154 6696 11160
rect 6656 10810 6684 11154
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6104 9166 6224 9194
rect 6104 8022 6132 9166
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6196 8634 6224 9046
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6656 8022 6684 8230
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5920 5846 5948 6054
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5644 5098 5672 5306
rect 5736 5234 5764 5646
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5644 4264 5672 5034
rect 5736 4826 5764 5170
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5644 4236 5764 4264
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5644 3738 5672 4082
rect 5736 4010 5764 4236
rect 5828 4214 5856 5646
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 5000 2446 5028 3062
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5092 2582 5120 2790
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 2134 0 2190 54
rect 3054 0 3110 54
rect 3882 54 4292 82
rect 4802 128 4858 480
rect 4802 76 4804 128
rect 4856 76 4858 128
rect 3882 0 3938 54
rect 4802 0 4858 76
rect 5552 82 5580 3062
rect 5920 2922 5948 4762
rect 6012 3670 6040 6598
rect 6104 6322 6132 7822
rect 6656 7546 6684 7958
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6196 6458 6224 6802
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 6196 5370 6224 5782
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6748 5166 6776 11183
rect 7116 10810 7144 11222
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6840 7886 6868 9998
rect 7024 8514 7052 10746
rect 7116 10538 7144 10746
rect 7300 10674 7328 11086
rect 7576 10690 7604 15014
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7760 13530 7788 14418
rect 8036 13814 8064 18226
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8312 17338 8340 17614
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8220 16658 8248 17070
rect 8312 17066 8340 17274
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8220 15570 8248 16594
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8208 14952 8260 14958
rect 8206 14920 8208 14929
rect 8260 14920 8262 14929
rect 8206 14855 8262 14864
rect 8220 14822 8248 14855
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8036 13802 8156 13814
rect 8036 13796 8168 13802
rect 8036 13786 8116 13796
rect 8116 13738 8168 13744
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 8036 12850 8064 13194
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7668 11762 7696 12378
rect 7760 12374 7788 12582
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7288 10668 7340 10674
rect 7576 10662 7788 10690
rect 7288 10610 7340 10616
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 7116 10266 7144 10474
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7116 9382 7144 9454
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7116 9042 7144 9318
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7024 8486 7144 8514
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6840 7478 6868 7822
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 7024 6866 7052 8298
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7116 5250 7144 8486
rect 7208 5778 7236 9386
rect 7300 9110 7328 10610
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7392 9178 7420 9522
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7484 8430 7512 10202
rect 7576 9926 7604 10542
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7576 9586 7604 9862
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7484 7206 7512 8366
rect 7576 8090 7604 9046
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7668 7410 7696 8026
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7484 6916 7512 7142
rect 7564 6928 7616 6934
rect 7484 6888 7564 6916
rect 7484 6186 7512 6888
rect 7564 6870 7616 6876
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7208 5370 7236 5714
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7116 5222 7236 5250
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6104 3670 6132 3878
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 6012 3194 6040 3606
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 5920 2310 5948 2858
rect 6012 2650 6040 3130
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6104 2582 6132 3606
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6196 3194 6224 3470
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6092 2576 6144 2582
rect 6092 2518 6144 2524
rect 6748 2378 6776 5102
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 5722 82 5778 480
rect 5552 54 5778 82
rect 5722 0 5778 54
rect 6550 82 6606 480
rect 6932 82 6960 3402
rect 7024 134 7052 4966
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 7116 4146 7144 4694
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 6550 54 6960 82
rect 7012 128 7064 134
rect 7012 70 7064 76
rect 7208 82 7236 5222
rect 7300 4690 7328 5850
rect 7484 4758 7512 6122
rect 7760 5778 7788 10662
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7668 5302 7696 5714
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7300 4282 7328 4626
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7668 4010 7696 4694
rect 7852 4154 7880 12718
rect 8036 12170 8064 12786
rect 8024 12164 8076 12170
rect 8024 12106 8076 12112
rect 8128 12050 8156 13738
rect 8220 13462 8248 14214
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8220 12986 8248 13398
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8036 12022 8156 12050
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7944 10062 7972 10950
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7944 9654 7972 9998
rect 8036 9994 8064 12022
rect 8220 11898 8248 12310
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 8128 11014 8156 11222
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8128 10198 8156 10950
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 8128 9722 8156 10134
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 8312 9042 8340 15438
rect 8404 13814 8432 18584
rect 8496 18426 8524 20402
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8496 18034 8524 18362
rect 8588 18222 8616 23446
rect 8680 21078 8708 23666
rect 8852 23588 8904 23594
rect 8852 23530 8904 23536
rect 8864 23254 8892 23530
rect 9692 23497 9720 24346
rect 10060 24274 10088 25298
rect 10428 24954 10456 25434
rect 10232 24948 10284 24954
rect 10232 24890 10284 24896
rect 10416 24948 10468 24954
rect 10416 24890 10468 24896
rect 10692 24948 10744 24954
rect 10692 24890 10744 24896
rect 9772 24268 9824 24274
rect 9772 24210 9824 24216
rect 10048 24268 10100 24274
rect 10048 24210 10100 24216
rect 9784 23526 9812 24210
rect 9772 23520 9824 23526
rect 9678 23488 9734 23497
rect 9508 23446 9678 23474
rect 9508 23322 9536 23446
rect 9772 23462 9824 23468
rect 9678 23423 9734 23432
rect 9496 23316 9548 23322
rect 9496 23258 9548 23264
rect 8852 23248 8904 23254
rect 8852 23190 8904 23196
rect 8864 22982 8892 23190
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 8852 22976 8904 22982
rect 8852 22918 8904 22924
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9416 22506 9444 22578
rect 9600 22574 9628 22918
rect 9588 22568 9640 22574
rect 9588 22510 9640 22516
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 9404 22500 9456 22506
rect 9404 22442 9456 22448
rect 9140 22234 9168 22442
rect 9496 22432 9548 22438
rect 9496 22374 9548 22380
rect 9128 22228 9180 22234
rect 9128 22170 9180 22176
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 8772 21622 8800 21966
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 8760 21616 8812 21622
rect 8760 21558 8812 21564
rect 8760 21480 8812 21486
rect 8864 21468 8892 21626
rect 9508 21486 9536 22374
rect 9496 21480 9548 21486
rect 8812 21440 8892 21468
rect 9416 21440 9496 21468
rect 8760 21422 8812 21428
rect 8772 21078 8800 21422
rect 8668 21072 8720 21078
rect 8668 21014 8720 21020
rect 8760 21072 8812 21078
rect 8760 21014 8812 21020
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 9416 20466 9444 21440
rect 9496 21422 9548 21428
rect 9496 20528 9548 20534
rect 9496 20470 9548 20476
rect 9404 20460 9456 20466
rect 9404 20402 9456 20408
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8496 18006 8616 18034
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8496 15094 8524 17478
rect 8588 17202 8616 18006
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8772 16114 8800 20334
rect 9508 20058 9536 20470
rect 9600 20058 9628 22510
rect 9692 21554 9720 23122
rect 9784 22642 9812 23462
rect 10244 23202 10272 24890
rect 10508 24744 10560 24750
rect 10508 24686 10560 24692
rect 10416 24676 10468 24682
rect 10416 24618 10468 24624
rect 10428 23662 10456 24618
rect 10520 24410 10548 24686
rect 10704 24682 10732 24890
rect 10692 24676 10744 24682
rect 10692 24618 10744 24624
rect 10508 24404 10560 24410
rect 10508 24346 10560 24352
rect 10600 23792 10652 23798
rect 10600 23734 10652 23740
rect 10416 23656 10468 23662
rect 10416 23598 10468 23604
rect 10324 23520 10376 23526
rect 10324 23462 10376 23468
rect 10336 23322 10364 23462
rect 10612 23338 10640 23734
rect 10690 23624 10746 23633
rect 10690 23559 10746 23568
rect 10324 23316 10376 23322
rect 10324 23258 10376 23264
rect 10520 23310 10640 23338
rect 10704 23322 10732 23559
rect 10692 23316 10744 23322
rect 10244 23174 10456 23202
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9864 22568 9916 22574
rect 9864 22510 9916 22516
rect 10048 22568 10100 22574
rect 10048 22510 10100 22516
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9784 22098 9812 22374
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9680 21344 9732 21350
rect 9784 21332 9812 22034
rect 9876 21894 9904 22510
rect 10060 22438 10088 22510
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9876 21486 9904 21830
rect 9864 21480 9916 21486
rect 10048 21480 10100 21486
rect 9864 21422 9916 21428
rect 9968 21440 10048 21468
rect 9732 21304 9812 21332
rect 9680 21286 9732 21292
rect 9692 20874 9720 21286
rect 9876 21010 9904 21422
rect 9968 21350 9996 21440
rect 10048 21422 10100 21428
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 9968 21078 9996 21286
rect 10060 21146 10088 21286
rect 10244 21146 10272 22510
rect 10428 22234 10456 23174
rect 10416 22228 10468 22234
rect 10416 22170 10468 22176
rect 10428 21690 10456 22170
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 10232 21140 10284 21146
rect 10232 21082 10284 21088
rect 9956 21072 10008 21078
rect 9956 21014 10008 21020
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 9864 21004 9916 21010
rect 9864 20946 9916 20952
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9784 20602 9812 20946
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9968 20398 9996 20742
rect 9956 20392 10008 20398
rect 9956 20334 10008 20340
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 9496 20052 9548 20058
rect 9496 19994 9548 20000
rect 9588 20052 9640 20058
rect 9588 19994 9640 20000
rect 9968 19922 9996 20334
rect 10152 19922 10180 20334
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 9956 19780 10008 19786
rect 9956 19722 10008 19728
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 9600 18426 9628 18906
rect 9784 18766 9812 19246
rect 9968 19242 9996 19722
rect 10152 19514 10180 19858
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9968 18970 9996 19178
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 10152 18834 10180 19450
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9588 18284 9640 18290
rect 9692 18272 9720 18634
rect 9784 18358 9812 18702
rect 10152 18426 10180 18770
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10232 18692 10284 18698
rect 10232 18634 10284 18640
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9640 18244 9720 18272
rect 9588 18226 9640 18232
rect 9312 18148 9364 18154
rect 9312 18090 9364 18096
rect 9324 17882 9352 18090
rect 9692 17882 9720 18244
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 8864 17116 8892 17546
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 9324 17134 9352 17818
rect 9784 17746 9812 18294
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9876 18086 9904 18226
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9784 17338 9812 17682
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 8944 17128 8996 17134
rect 8864 17088 8944 17116
rect 8944 17070 8996 17076
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 8956 16726 8984 17070
rect 9324 16794 9352 17070
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 8944 16720 8996 16726
rect 8864 16680 8944 16708
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8864 16046 8892 16680
rect 8944 16662 8996 16668
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 9324 16046 9352 16730
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 8864 15638 8892 15982
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 8852 15632 8904 15638
rect 8852 15574 8904 15580
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8484 15088 8536 15094
rect 8484 15030 8536 15036
rect 8588 14958 8616 15302
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8496 14482 8524 14758
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8588 14278 8616 14894
rect 8864 14618 8892 15574
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 9416 15162 9444 15642
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 9600 14482 9628 15846
rect 9784 15570 9812 16934
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9968 15706 9996 16594
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 10060 16250 10088 16458
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9784 14618 9812 15506
rect 9864 14816 9916 14822
rect 9968 14804 9996 15506
rect 9916 14776 9996 14804
rect 9864 14758 9916 14764
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9876 14550 9904 14758
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9588 14476 9640 14482
rect 9508 14436 9588 14464
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8404 13786 8524 13814
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8404 12986 8432 13670
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8404 12646 8432 12922
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8496 9518 8524 13786
rect 8588 12594 8616 14214
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 9508 14074 9536 14436
rect 9588 14418 9640 14424
rect 9876 14074 9904 14486
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 10152 14006 10180 16526
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9312 13796 9364 13802
rect 9364 13756 9444 13784
rect 9312 13738 9364 13744
rect 9416 13705 9444 13756
rect 9402 13696 9458 13705
rect 9402 13631 9458 13640
rect 9508 13410 9536 13874
rect 10244 13814 10272 18634
rect 10428 18222 10456 18702
rect 10416 18216 10468 18222
rect 10416 18158 10468 18164
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10336 15162 10364 16662
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10520 13814 10548 23310
rect 10692 23258 10744 23264
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10704 19922 10732 20266
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10612 18970 10640 19790
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10612 17882 10640 18906
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10612 17134 10640 17818
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10612 16590 10640 17070
rect 10704 16658 10732 18702
rect 10796 18698 10824 28920
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10796 17814 10824 18022
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10796 16794 10824 17070
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10152 13786 10272 13814
rect 10336 13786 10548 13814
rect 10612 13802 10640 14758
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10600 13796 10652 13802
rect 10048 13456 10100 13462
rect 9508 13382 9628 13410
rect 10048 13398 10100 13404
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8668 12708 8720 12714
rect 8772 12696 8800 13126
rect 8720 12668 8800 12696
rect 8668 12650 8720 12656
rect 8588 12566 8708 12594
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8588 11354 8616 12174
rect 8680 11558 8708 12566
rect 8772 12170 8800 12668
rect 8864 12374 8892 13262
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 9508 12374 9536 13262
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8680 9586 8708 11494
rect 8772 11082 8800 12106
rect 8864 11812 8892 12310
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 8944 11824 8996 11830
rect 8864 11784 8944 11812
rect 8944 11766 8996 11772
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9508 11354 9536 11562
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8772 10198 8800 11018
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 9404 10736 9456 10742
rect 9404 10678 9456 10684
rect 9416 10538 9444 10678
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9324 10266 9352 10474
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8666 9480 8722 9489
rect 8666 9415 8722 9424
rect 8680 9382 8708 9415
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8220 8498 8248 8774
rect 8312 8634 8340 8978
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8220 8294 8248 8434
rect 8588 8430 8616 9114
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8220 7546 8248 7958
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8220 5914 8248 6802
rect 8496 6662 8524 7822
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8404 6458 8432 6598
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8220 4826 8248 4966
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8220 4282 8248 4762
rect 8404 4758 8432 5034
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 7852 4126 7972 4154
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7668 3738 7696 3946
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7944 2514 7972 4126
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8220 3670 8248 3878
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8220 3194 8248 3606
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8220 2904 8248 3130
rect 8312 3058 8340 3674
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8300 2916 8352 2922
rect 8220 2876 8300 2904
rect 8220 2650 8248 2876
rect 8300 2858 8352 2864
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8680 2582 8708 9318
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8864 8430 8892 8842
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8864 8022 8892 8366
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8864 7460 8892 7958
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 8944 7472 8996 7478
rect 8864 7432 8944 7460
rect 8944 7414 8996 7420
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 9324 6186 9352 7822
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7410 9536 7686
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9496 7268 9548 7274
rect 9496 7210 9548 7216
rect 9508 7002 9536 7210
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9600 6798 9628 13382
rect 10060 12850 10088 13398
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10152 12424 10180 13786
rect 10060 12396 10180 12424
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9968 11626 9996 12242
rect 9956 11620 10008 11626
rect 9956 11562 10008 11568
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9692 9382 9720 10066
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 9110 9720 9318
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9692 7478 9720 9046
rect 9968 8566 9996 11562
rect 10060 10130 10088 12396
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10152 11558 10180 12242
rect 10336 12102 10364 13786
rect 10600 13738 10652 13744
rect 10612 13462 10640 13738
rect 10704 13734 10732 14214
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10704 12782 10732 13670
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10704 12442 10732 12718
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10428 11286 10456 11766
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10244 10810 10272 11222
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10428 10674 10456 11222
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10612 10810 10640 11086
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10888 10606 10916 35430
rect 10980 34610 11008 35498
rect 10968 34604 11020 34610
rect 11020 34564 11100 34592
rect 10968 34546 11020 34552
rect 10968 34128 11020 34134
rect 10968 34070 11020 34076
rect 10980 33658 11008 34070
rect 11072 33930 11100 34564
rect 11060 33924 11112 33930
rect 11060 33866 11112 33872
rect 10968 33652 11020 33658
rect 10968 33594 11020 33600
rect 10980 33046 11008 33594
rect 10968 33040 11020 33046
rect 10968 32982 11020 32988
rect 11072 31346 11100 33866
rect 11256 31890 11284 35702
rect 11348 34746 11376 39630
rect 11532 39630 11942 39658
rect 11428 35080 11480 35086
rect 11428 35022 11480 35028
rect 11336 34740 11388 34746
rect 11336 34682 11388 34688
rect 11336 33992 11388 33998
rect 11336 33934 11388 33940
rect 11348 32774 11376 33934
rect 11440 33538 11468 35022
rect 11532 33658 11560 39630
rect 11886 39520 11942 39630
rect 12636 39630 12862 39658
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 12440 36712 12492 36718
rect 12440 36654 12492 36660
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 12164 35148 12216 35154
rect 12164 35090 12216 35096
rect 12176 34678 12204 35090
rect 12164 34672 12216 34678
rect 12164 34614 12216 34620
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 12176 34066 12204 34614
rect 12452 34542 12480 36654
rect 12636 35018 12664 39630
rect 12806 39520 12862 39630
rect 13464 39630 13782 39658
rect 13464 35834 13492 39630
rect 13726 39520 13782 39630
rect 14554 39658 14610 40000
rect 15474 39658 15530 40000
rect 14554 39630 14688 39658
rect 14554 39520 14610 39630
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 13452 35828 13504 35834
rect 13452 35770 13504 35776
rect 14660 35290 14688 39630
rect 15474 39630 15608 39658
rect 15474 39520 15530 39630
rect 15474 38176 15530 38185
rect 15474 38111 15530 38120
rect 14648 35284 14700 35290
rect 14648 35226 14700 35232
rect 12992 35148 13044 35154
rect 12992 35090 13044 35096
rect 12624 35012 12676 35018
rect 12624 34954 12676 34960
rect 12532 34944 12584 34950
rect 12532 34886 12584 34892
rect 12440 34536 12492 34542
rect 12440 34478 12492 34484
rect 12164 34060 12216 34066
rect 12164 34002 12216 34008
rect 12440 34060 12492 34066
rect 12440 34002 12492 34008
rect 12164 33856 12216 33862
rect 12164 33798 12216 33804
rect 11520 33652 11572 33658
rect 11520 33594 11572 33600
rect 11440 33510 11560 33538
rect 11532 33114 11560 33510
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11520 33108 11572 33114
rect 11440 33068 11520 33096
rect 11336 32768 11388 32774
rect 11336 32710 11388 32716
rect 11440 31940 11468 33068
rect 11520 33050 11572 33056
rect 11704 33040 11756 33046
rect 11704 32982 11756 32988
rect 11520 32904 11572 32910
rect 11520 32846 11572 32852
rect 11532 32026 11560 32846
rect 11716 32570 11744 32982
rect 12176 32570 12204 33798
rect 12256 33380 12308 33386
rect 12256 33322 12308 33328
rect 11704 32564 11756 32570
rect 11704 32506 11756 32512
rect 12164 32564 12216 32570
rect 12164 32506 12216 32512
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11520 32020 11572 32026
rect 11520 31962 11572 31968
rect 11348 31912 11468 31940
rect 11244 31884 11296 31890
rect 11244 31826 11296 31832
rect 11060 31340 11112 31346
rect 11060 31282 11112 31288
rect 10968 31204 11020 31210
rect 10968 31146 11020 31152
rect 10980 29850 11008 31146
rect 11072 30938 11100 31282
rect 11256 31142 11284 31826
rect 11244 31136 11296 31142
rect 11244 31078 11296 31084
rect 11060 30932 11112 30938
rect 11060 30874 11112 30880
rect 11348 30734 11376 31912
rect 11520 31884 11572 31890
rect 11520 31826 11572 31832
rect 11428 30864 11480 30870
rect 11428 30806 11480 30812
rect 11336 30728 11388 30734
rect 11336 30670 11388 30676
rect 11348 30258 11376 30670
rect 11440 30394 11468 30806
rect 11428 30388 11480 30394
rect 11428 30330 11480 30336
rect 11336 30252 11388 30258
rect 11336 30194 11388 30200
rect 10968 29844 11020 29850
rect 10968 29786 11020 29792
rect 10968 28620 11020 28626
rect 10968 28562 11020 28568
rect 10980 27946 11008 28562
rect 11060 28552 11112 28558
rect 11060 28494 11112 28500
rect 11072 28218 11100 28494
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 10968 27940 11020 27946
rect 10968 27882 11020 27888
rect 10980 19990 11008 27882
rect 11532 27656 11560 31826
rect 12072 31408 12124 31414
rect 12072 31350 12124 31356
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11980 29776 12032 29782
rect 11980 29718 12032 29724
rect 11888 29640 11940 29646
rect 11888 29582 11940 29588
rect 11900 29306 11928 29582
rect 11888 29300 11940 29306
rect 11888 29242 11940 29248
rect 11992 29102 12020 29718
rect 12084 29458 12112 31350
rect 12164 31204 12216 31210
rect 12164 31146 12216 31152
rect 12176 30734 12204 31146
rect 12164 30728 12216 30734
rect 12164 30670 12216 30676
rect 12176 30326 12204 30670
rect 12164 30320 12216 30326
rect 12164 30262 12216 30268
rect 12176 29646 12204 30262
rect 12164 29640 12216 29646
rect 12164 29582 12216 29588
rect 12084 29430 12204 29458
rect 11980 29096 12032 29102
rect 11980 29038 12032 29044
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11440 27628 11560 27656
rect 11152 27464 11204 27470
rect 11152 27406 11204 27412
rect 11164 27062 11192 27406
rect 11152 27056 11204 27062
rect 11058 27024 11114 27033
rect 11152 26998 11204 27004
rect 11058 26959 11114 26968
rect 11072 26926 11100 26959
rect 11060 26920 11112 26926
rect 11060 26862 11112 26868
rect 11060 26784 11112 26790
rect 11060 26726 11112 26732
rect 11072 26382 11100 26726
rect 11060 26376 11112 26382
rect 11060 26318 11112 26324
rect 11164 26246 11192 26998
rect 11244 26308 11296 26314
rect 11244 26250 11296 26256
rect 11152 26240 11204 26246
rect 11152 26182 11204 26188
rect 11164 25974 11192 26182
rect 11152 25968 11204 25974
rect 11152 25910 11204 25916
rect 11256 24818 11284 26250
rect 11336 25764 11388 25770
rect 11336 25706 11388 25712
rect 11348 25498 11376 25706
rect 11336 25492 11388 25498
rect 11336 25434 11388 25440
rect 11440 25378 11468 27628
rect 11980 27600 12032 27606
rect 11980 27542 12032 27548
rect 11520 27464 11572 27470
rect 11520 27406 11572 27412
rect 11532 26858 11560 27406
rect 11520 26852 11572 26858
rect 11520 26794 11572 26800
rect 11348 25350 11468 25378
rect 11244 24812 11296 24818
rect 11244 24754 11296 24760
rect 11256 24206 11284 24754
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 11256 23662 11284 24142
rect 11244 23656 11296 23662
rect 11150 23624 11206 23633
rect 11244 23598 11296 23604
rect 11150 23559 11206 23568
rect 11164 21146 11192 23559
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 11072 19514 11100 20470
rect 11164 20398 11192 21082
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 11256 20602 11284 20946
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11152 20392 11204 20398
rect 11152 20334 11204 20340
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10980 16726 11008 18022
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11256 17134 11284 17614
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 10968 15972 11020 15978
rect 10968 15914 11020 15920
rect 10980 15162 11008 15914
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 11072 14414 11100 16934
rect 11348 16794 11376 25350
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 11440 24342 11468 24550
rect 11428 24336 11480 24342
rect 11428 24278 11480 24284
rect 11440 23866 11468 24278
rect 11532 24206 11560 26794
rect 11992 26790 12020 27542
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 12072 26784 12124 26790
rect 12072 26726 12124 26732
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11704 26376 11756 26382
rect 11704 26318 11756 26324
rect 11716 26042 11744 26318
rect 11704 26036 11756 26042
rect 11704 25978 11756 25984
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11796 25424 11848 25430
rect 11796 25366 11848 25372
rect 11808 24954 11836 25366
rect 11992 25362 12020 26726
rect 12084 26382 12112 26726
rect 12072 26376 12124 26382
rect 12176 26364 12204 29430
rect 12268 26926 12296 33322
rect 12452 32842 12480 34002
rect 12544 33522 12572 34886
rect 13004 34542 13032 35090
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 12992 34536 13044 34542
rect 12992 34478 13044 34484
rect 13634 34504 13690 34513
rect 12532 33516 12584 33522
rect 12532 33458 12584 33464
rect 12808 33516 12860 33522
rect 12808 33458 12860 33464
rect 12544 33114 12572 33458
rect 12532 33108 12584 33114
rect 12532 33050 12584 33056
rect 12820 33046 12848 33458
rect 12808 33040 12860 33046
rect 12808 32982 12860 32988
rect 13004 32978 13032 34478
rect 13634 34439 13690 34448
rect 13452 34060 13504 34066
rect 13452 34002 13504 34008
rect 13464 33658 13492 34002
rect 13452 33652 13504 33658
rect 13452 33594 13504 33600
rect 12992 32972 13044 32978
rect 12992 32914 13044 32920
rect 12440 32836 12492 32842
rect 12440 32778 12492 32784
rect 12348 32224 12400 32230
rect 12348 32166 12400 32172
rect 12256 26920 12308 26926
rect 12256 26862 12308 26868
rect 12256 26376 12308 26382
rect 12176 26336 12256 26364
rect 12072 26318 12124 26324
rect 12256 26318 12308 26324
rect 12268 25702 12296 26318
rect 12256 25696 12308 25702
rect 12256 25638 12308 25644
rect 11980 25356 12032 25362
rect 11980 25298 12032 25304
rect 12072 25288 12124 25294
rect 12072 25230 12124 25236
rect 11796 24948 11848 24954
rect 11796 24890 11848 24896
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 11808 23594 11836 24142
rect 12084 24070 12112 25230
rect 12072 24064 12124 24070
rect 12072 24006 12124 24012
rect 12084 23730 12112 24006
rect 12268 23730 12296 25638
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 12360 23610 12388 32166
rect 12452 31226 12480 32778
rect 13004 32230 13032 32914
rect 12992 32224 13044 32230
rect 12992 32166 13044 32172
rect 12452 31198 12572 31226
rect 12440 31136 12492 31142
rect 12440 31078 12492 31084
rect 12452 27538 12480 31078
rect 12440 27532 12492 27538
rect 12440 27474 12492 27480
rect 12544 27418 12572 31198
rect 13268 27532 13320 27538
rect 13268 27474 13320 27480
rect 12452 27390 12572 27418
rect 12452 24256 12480 27390
rect 12532 27328 12584 27334
rect 12532 27270 12584 27276
rect 12544 25906 12572 27270
rect 12716 26920 12768 26926
rect 12716 26862 12768 26868
rect 12624 26512 12676 26518
rect 12624 26454 12676 26460
rect 12636 26246 12664 26454
rect 12624 26240 12676 26246
rect 12624 26182 12676 26188
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12544 25498 12572 25842
rect 12636 25770 12664 26182
rect 12624 25764 12676 25770
rect 12624 25706 12676 25712
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12544 24410 12572 24550
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12624 24268 12676 24274
rect 12452 24228 12624 24256
rect 12624 24210 12676 24216
rect 12636 23798 12664 24210
rect 12624 23792 12676 23798
rect 12624 23734 12676 23740
rect 12440 23724 12492 23730
rect 12440 23666 12492 23672
rect 11796 23588 11848 23594
rect 11796 23530 11848 23536
rect 11992 23582 12388 23610
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11520 23248 11572 23254
rect 11520 23190 11572 23196
rect 11428 23112 11480 23118
rect 11428 23054 11480 23060
rect 11440 22778 11468 23054
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11532 22438 11560 23190
rect 11520 22432 11572 22438
rect 11520 22374 11572 22380
rect 11532 22234 11560 22374
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11520 22228 11572 22234
rect 11520 22170 11572 22176
rect 11520 22092 11572 22098
rect 11520 22034 11572 22040
rect 11532 21350 11560 22034
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11532 20330 11560 20946
rect 11520 20324 11572 20330
rect 11520 20266 11572 20272
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11532 19514 11560 19858
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11428 19440 11480 19446
rect 11428 19382 11480 19388
rect 11440 18834 11468 19382
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11440 18426 11468 18770
rect 11428 18420 11480 18426
rect 11428 18362 11480 18368
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 11532 17746 11560 18226
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11532 17338 11560 17682
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11992 17202 12020 23582
rect 12164 23520 12216 23526
rect 12452 23474 12480 23666
rect 12164 23462 12216 23468
rect 12176 23254 12204 23462
rect 12360 23446 12480 23474
rect 12360 23322 12388 23446
rect 12348 23316 12400 23322
rect 12348 23258 12400 23264
rect 12164 23248 12216 23254
rect 12164 23190 12216 23196
rect 12360 22778 12388 23258
rect 12348 22772 12400 22778
rect 12348 22714 12400 22720
rect 12072 22568 12124 22574
rect 12072 22510 12124 22516
rect 12532 22568 12584 22574
rect 12532 22510 12584 22516
rect 12084 22098 12112 22510
rect 12544 22166 12572 22510
rect 12624 22500 12676 22506
rect 12624 22442 12676 22448
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 12084 21146 12112 22034
rect 12164 21956 12216 21962
rect 12164 21898 12216 21904
rect 12176 21350 12204 21898
rect 12636 21690 12664 22442
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 12072 21140 12124 21146
rect 12072 21082 12124 21088
rect 12072 20868 12124 20874
rect 12176 20856 12204 21286
rect 12124 20828 12204 20856
rect 12072 20810 12124 20816
rect 12084 20262 12112 20810
rect 12256 20324 12308 20330
rect 12256 20266 12308 20272
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11532 17066 11560 17138
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11164 15706 11192 16050
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10980 14074 11008 14214
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 9968 7954 9996 8502
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9784 6798 9812 7210
rect 9876 6798 9904 7754
rect 9968 7546 9996 7890
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9416 6186 9444 6394
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9324 5914 9352 6122
rect 9508 5914 9536 6598
rect 9784 6118 9812 6734
rect 9876 6390 9904 6734
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9968 6322 9996 6870
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 9324 5234 9352 5850
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9692 5370 9720 5714
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 8772 3126 8800 5170
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8864 4214 8892 4422
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9232 3670 9260 4082
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9416 3534 9444 5238
rect 9784 4214 9812 6054
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9968 4282 9996 4626
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9678 4040 9734 4049
rect 9678 3975 9734 3984
rect 9692 3602 9720 3975
rect 10060 3641 10088 5102
rect 10888 4282 10916 10542
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10980 4282 11008 4558
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 11072 4154 11100 14010
rect 11256 11694 11284 16526
rect 11336 14476 11388 14482
rect 11388 14436 11468 14464
rect 11336 14418 11388 14424
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 11348 12288 11376 14282
rect 11440 13734 11468 14436
rect 11532 14074 11560 17002
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11716 14890 11744 15438
rect 11808 15162 11836 15574
rect 11992 15502 12020 15914
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11808 14958 11836 15098
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11428 13728 11480 13734
rect 11426 13696 11428 13705
rect 11480 13696 11482 13705
rect 11426 13631 11482 13640
rect 11440 13605 11468 13631
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11440 13297 11468 13330
rect 11426 13288 11482 13297
rect 11426 13223 11482 13232
rect 11440 12986 11468 13223
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 12084 12753 12112 20198
rect 12164 16176 12216 16182
rect 12164 16118 12216 16124
rect 12070 12744 12126 12753
rect 12070 12679 12126 12688
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11428 12300 11480 12306
rect 11348 12260 11428 12288
rect 11428 12242 11480 12248
rect 11440 11694 11468 12242
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11348 9625 11376 11494
rect 11334 9616 11390 9625
rect 11334 9551 11390 9560
rect 11072 4126 11284 4154
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10046 3632 10102 3641
rect 9680 3596 9732 3602
rect 10046 3567 10102 3576
rect 10232 3596 10284 3602
rect 9680 3538 9732 3544
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 7470 82 7526 480
rect 7208 54 7526 82
rect 8312 82 8340 2246
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 8390 82 8446 480
rect 8312 54 8446 82
rect 6550 0 6606 54
rect 7470 0 7526 54
rect 8390 0 8446 54
rect 9218 82 9274 480
rect 9324 82 9352 3334
rect 9416 3194 9444 3470
rect 10060 3194 10088 3567
rect 10232 3538 10284 3544
rect 10244 3194 10272 3538
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 9692 2990 9720 3130
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 9218 54 9352 82
rect 9876 82 9904 2790
rect 10428 2446 10456 2790
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10138 82 10194 480
rect 9876 54 10194 82
rect 10704 82 10732 3878
rect 11256 3466 11284 4126
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11440 2514 11468 11630
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11624 10810 11652 11222
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11992 10470 12020 11086
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11992 9722 12020 10406
rect 11980 9716 12032 9722
rect 11980 9658 12032 9664
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 12176 5953 12204 16118
rect 12268 9081 12296 20266
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12452 18222 12480 19314
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12360 15910 12388 16594
rect 12728 16590 12756 26862
rect 13280 26790 13308 27474
rect 13648 27130 13676 34439
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 15488 31890 15516 38111
rect 15580 34202 15608 39630
rect 15568 34196 15620 34202
rect 15568 34138 15620 34144
rect 15476 31884 15528 31890
rect 15476 31826 15528 31832
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14738 27296 14794 27305
rect 14289 27228 14585 27248
rect 14738 27231 14794 27240
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 13636 27124 13688 27130
rect 13636 27066 13688 27072
rect 13268 26784 13320 26790
rect 13268 26726 13320 26732
rect 13084 26444 13136 26450
rect 13084 26386 13136 26392
rect 13096 26042 13124 26386
rect 13084 26036 13136 26042
rect 13084 25978 13136 25984
rect 13096 24818 13124 25978
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 12900 24744 12952 24750
rect 12900 24686 12952 24692
rect 12912 24206 12940 24686
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 13082 19952 13138 19961
rect 13082 19887 13138 19896
rect 13096 18834 13124 19887
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 13096 17746 13124 18770
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 12820 17338 12848 17682
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12820 16726 12848 17274
rect 12912 17066 12940 17546
rect 13096 17270 13124 17682
rect 13084 17264 13136 17270
rect 13084 17206 13136 17212
rect 12900 17060 12952 17066
rect 12900 17002 12952 17008
rect 12808 16720 12860 16726
rect 12808 16662 12860 16668
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12912 16522 12940 17002
rect 12900 16516 12952 16522
rect 12900 16458 12952 16464
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12254 9072 12310 9081
rect 12254 9007 12310 9016
rect 12162 5944 12218 5953
rect 12162 5879 12218 5888
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 11624 3194 11652 3402
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 12360 2417 12388 15846
rect 13280 14346 13308 26726
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 13544 25356 13596 25362
rect 13544 25298 13596 25304
rect 13556 24954 13584 25298
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 13544 24948 13596 24954
rect 13544 24890 13596 24896
rect 13556 23769 13584 24890
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 13542 23760 13598 23769
rect 13542 23695 13598 23704
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 13452 22568 13504 22574
rect 13452 22510 13504 22516
rect 13464 21418 13492 22510
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 13452 21412 13504 21418
rect 13452 21354 13504 21360
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14752 20534 14780 27231
rect 14740 20528 14792 20534
rect 14740 20470 14792 20476
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13556 15978 13584 16594
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14752 16289 14780 17002
rect 14738 16280 14794 16289
rect 14738 16215 14794 16224
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 13268 14340 13320 14346
rect 13268 14282 13320 14288
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12346 2408 12402 2417
rect 11704 2372 11756 2378
rect 12346 2343 12402 2352
rect 11704 2314 11756 2320
rect 11058 82 11114 480
rect 10704 54 11114 82
rect 11716 82 11744 2314
rect 11886 82 11942 480
rect 11716 54 11942 82
rect 12544 82 12572 2858
rect 13188 2514 13216 5306
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 12806 82 12862 480
rect 12544 54 12862 82
rect 9218 0 9274 54
rect 10138 0 10194 54
rect 11058 0 11114 54
rect 11886 0 11942 54
rect 12806 0 12862 54
rect 13726 128 13782 480
rect 13726 76 13728 128
rect 13780 76 13782 128
rect 13726 0 13782 76
rect 14554 82 14610 480
rect 14660 82 14688 2314
rect 14554 54 14688 82
rect 15474 82 15530 480
rect 15580 82 15608 2586
rect 15474 54 15608 82
rect 14554 0 14610 54
rect 15474 0 15530 54
<< via2 >>
rect 110 12416 166 12472
rect 110 2488 166 2544
rect 2318 6840 2374 6896
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3146 23604 3148 23624
rect 3148 23604 3200 23624
rect 3200 23604 3202 23624
rect 3146 23568 3202 23604
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 5814 37168 5870 37224
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 4158 21936 4214 21992
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3974 19352 4030 19408
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3514 16904 3570 16960
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 2594 3032 2650 3088
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3514 11736 3570 11792
rect 4250 19352 4306 19408
rect 3974 11328 4030 11384
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 5814 26968 5870 27024
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6734 26832 6790 26888
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 4434 11736 4490 11792
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3974 9560 4030 9616
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 3514 3576 3570 3632
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 4894 13232 4950 13288
rect 5262 13232 5318 13288
rect 5078 9460 5080 9480
rect 5080 9460 5132 9480
rect 5132 9460 5134 9480
rect 5078 9424 5134 9460
rect 4618 3984 4674 4040
rect 4618 3032 4674 3088
rect 6734 23432 6790 23488
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 7378 23704 7434 23760
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6182 14864 6238 14920
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 8482 31864 8538 31920
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 10230 30776 10286 30832
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8206 23704 8262 23760
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6734 11192 6790 11248
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 8206 14900 8208 14920
rect 8208 14900 8260 14920
rect 8260 14900 8262 14920
rect 8206 14864 8262 14900
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 9678 23432 9734 23488
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 10690 23568 10746 23624
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 9402 13640 9458 13696
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8666 9424 8722 9480
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 15474 38120 15530 38176
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11058 26968 11114 27024
rect 11150 23568 11206 23624
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 13634 34448 13690 34504
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 9678 3984 9734 4040
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11426 13676 11428 13696
rect 11428 13676 11480 13696
rect 11480 13676 11482 13696
rect 11426 13640 11482 13676
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11426 13232 11482 13288
rect 12070 12688 12126 12744
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 11334 9560 11390 9616
rect 10046 3576 10102 3632
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14738 27240 14794 27296
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 13082 19896 13138 19952
rect 12254 9016 12310 9072
rect 12162 5888 12218 5944
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 13542 23704 13598 23760
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14738 16224 14794 16280
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 12346 2352 12402 2408
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
<< metal3 >>
rect 15520 38181 16000 38208
rect 15469 38178 16000 38181
rect 15388 38176 16000 38178
rect 15388 38120 15474 38176
rect 15530 38120 16000 38176
rect 15388 38118 16000 38120
rect 15469 38115 16000 38118
rect 15520 38088 16000 38115
rect 6277 37568 6597 37569
rect 0 37408 480 37528
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 62 37226 122 37408
rect 5809 37226 5875 37229
rect 62 37224 5875 37226
rect 62 37168 5814 37224
rect 5870 37168 5875 37224
rect 62 37166 5875 37168
rect 5809 37163 5875 37166
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 13629 34506 13695 34509
rect 15520 34506 16000 34536
rect 13629 34504 16000 34506
rect 13629 34448 13634 34504
rect 13690 34448 16000 34504
rect 13629 34446 16000 34448
rect 13629 34443 13695 34446
rect 15520 34416 16000 34446
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 0 32376 480 32496
rect 62 31922 122 32376
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 8477 31922 8543 31925
rect 62 31920 8543 31922
rect 62 31864 8482 31920
rect 8538 31864 8543 31920
rect 62 31862 8543 31864
rect 8477 31859 8543 31862
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 10225 30834 10291 30837
rect 15520 30834 16000 30864
rect 10225 30832 16000 30834
rect 10225 30776 10230 30832
rect 10286 30776 16000 30832
rect 10225 30774 16000 30776
rect 10225 30771 10291 30774
rect 15520 30744 16000 30774
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 29887 11930 29888
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 0 27344 480 27464
rect 62 26890 122 27344
rect 14733 27298 14799 27301
rect 15520 27298 16000 27328
rect 14733 27296 16000 27298
rect 14733 27240 14738 27296
rect 14794 27240 16000 27296
rect 14733 27238 16000 27240
rect 14733 27235 14799 27238
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 15520 27208 16000 27238
rect 14277 27167 14597 27168
rect 5809 27026 5875 27029
rect 11053 27026 11119 27029
rect 5809 27024 11119 27026
rect 5809 26968 5814 27024
rect 5870 26968 11058 27024
rect 11114 26968 11119 27024
rect 5809 26966 11119 26968
rect 5809 26963 5875 26966
rect 11053 26963 11119 26966
rect 6729 26890 6795 26893
rect 62 26888 6795 26890
rect 62 26832 6734 26888
rect 6790 26832 6795 26888
rect 62 26830 6795 26832
rect 6729 26827 6795 26830
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 7373 23762 7439 23765
rect 8201 23762 8267 23765
rect 13537 23762 13603 23765
rect 7373 23760 13603 23762
rect 7373 23704 7378 23760
rect 7434 23704 8206 23760
rect 8262 23704 13542 23760
rect 13598 23704 13603 23760
rect 7373 23702 13603 23704
rect 7373 23699 7439 23702
rect 8201 23699 8267 23702
rect 13537 23699 13603 23702
rect 3141 23626 3207 23629
rect 10685 23626 10751 23629
rect 3141 23624 10751 23626
rect 3141 23568 3146 23624
rect 3202 23568 10690 23624
rect 10746 23568 10751 23624
rect 3141 23566 10751 23568
rect 3141 23563 3207 23566
rect 10685 23563 10751 23566
rect 11145 23626 11211 23629
rect 15520 23626 16000 23656
rect 11145 23624 16000 23626
rect 11145 23568 11150 23624
rect 11206 23568 16000 23624
rect 11145 23566 16000 23568
rect 11145 23563 11211 23566
rect 15520 23536 16000 23566
rect 6729 23490 6795 23493
rect 9673 23490 9739 23493
rect 6729 23488 9739 23490
rect 6729 23432 6734 23488
rect 6790 23432 9678 23488
rect 9734 23432 9739 23488
rect 6729 23430 9739 23432
rect 6729 23427 6795 23430
rect 9673 23427 9739 23430
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 0 22448 480 22568
rect 62 21994 122 22448
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 4153 21994 4219 21997
rect 62 21992 4219 21994
rect 62 21936 4158 21992
rect 4214 21936 4219 21992
rect 62 21934 4219 21936
rect 4153 21931 4219 21934
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 13077 19954 13143 19957
rect 15520 19954 16000 19984
rect 13077 19952 16000 19954
rect 13077 19896 13082 19952
rect 13138 19896 16000 19952
rect 13077 19894 16000 19896
rect 13077 19891 13143 19894
rect 15520 19864 16000 19894
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 3969 19410 4035 19413
rect 4245 19410 4311 19413
rect 3969 19408 4311 19410
rect 3969 19352 3974 19408
rect 4030 19352 4250 19408
rect 4306 19352 4311 19408
rect 3969 19350 4311 19352
rect 3969 19347 4035 19350
rect 4245 19347 4311 19350
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 0 17416 480 17536
rect 3610 17440 3930 17441
rect 62 16962 122 17416
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 3509 16962 3575 16965
rect 62 16960 3575 16962
rect 62 16904 3514 16960
rect 3570 16904 3575 16960
rect 62 16902 3575 16904
rect 3509 16899 3575 16902
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 14733 16282 14799 16285
rect 15520 16282 16000 16312
rect 14733 16280 16000 16282
rect 14733 16224 14738 16280
rect 14794 16224 16000 16280
rect 14733 16222 16000 16224
rect 14733 16219 14799 16222
rect 15520 16192 16000 16222
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 6177 14922 6243 14925
rect 8201 14922 8267 14925
rect 6177 14920 8267 14922
rect 6177 14864 6182 14920
rect 6238 14864 8206 14920
rect 8262 14864 8267 14920
rect 6177 14862 8267 14864
rect 6177 14859 6243 14862
rect 8201 14859 8267 14862
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 9397 13698 9463 13701
rect 11421 13698 11487 13701
rect 9397 13696 11487 13698
rect 9397 13640 9402 13696
rect 9458 13640 11426 13696
rect 11482 13640 11487 13696
rect 9397 13638 11487 13640
rect 9397 13635 9463 13638
rect 11421 13635 11487 13638
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 4889 13290 4955 13293
rect 5257 13290 5323 13293
rect 11421 13290 11487 13293
rect 4889 13288 11487 13290
rect 4889 13232 4894 13288
rect 4950 13232 5262 13288
rect 5318 13232 11426 13288
rect 11482 13232 11487 13288
rect 4889 13230 11487 13232
rect 4889 13227 4955 13230
rect 5257 13227 5323 13230
rect 11421 13227 11487 13230
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 12065 12746 12131 12749
rect 15520 12746 16000 12776
rect 12065 12744 16000 12746
rect 12065 12688 12070 12744
rect 12126 12688 16000 12744
rect 12065 12686 16000 12688
rect 12065 12683 12131 12686
rect 15520 12656 16000 12686
rect 6277 12544 6597 12545
rect 0 12472 480 12504
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 0 12416 110 12472
rect 166 12416 480 12472
rect 0 12384 480 12416
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 3509 11794 3575 11797
rect 4429 11794 4495 11797
rect 3509 11792 4495 11794
rect 3509 11736 3514 11792
rect 3570 11736 4434 11792
rect 4490 11736 4495 11792
rect 3509 11734 4495 11736
rect 3509 11731 3575 11734
rect 4429 11731 4495 11734
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 3969 11386 4035 11389
rect 3969 11384 4170 11386
rect 3969 11328 3974 11384
rect 4030 11328 4170 11384
rect 3969 11326 4170 11328
rect 3969 11323 4035 11326
rect 4110 11250 4170 11326
rect 6729 11250 6795 11253
rect 4110 11248 6795 11250
rect 4110 11192 6734 11248
rect 6790 11192 6795 11248
rect 4110 11190 6795 11192
rect 6729 11187 6795 11190
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 3969 9618 4035 9621
rect 11329 9618 11395 9621
rect 3969 9616 11395 9618
rect 3969 9560 3974 9616
rect 4030 9560 11334 9616
rect 11390 9560 11395 9616
rect 3969 9558 11395 9560
rect 3969 9555 4035 9558
rect 11329 9555 11395 9558
rect 5073 9482 5139 9485
rect 8661 9482 8727 9485
rect 5073 9480 8727 9482
rect 5073 9424 5078 9480
rect 5134 9424 8666 9480
rect 8722 9424 8727 9480
rect 5073 9422 8727 9424
rect 5073 9419 5139 9422
rect 8661 9419 8727 9422
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 12249 9074 12315 9077
rect 15520 9074 16000 9104
rect 12249 9072 16000 9074
rect 12249 9016 12254 9072
rect 12310 9016 16000 9072
rect 12249 9014 16000 9016
rect 12249 9011 12315 9014
rect 15520 8984 16000 9014
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 0 7352 480 7472
rect 62 6898 122 7352
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 2313 6898 2379 6901
rect 62 6896 2379 6898
rect 62 6840 2318 6896
rect 2374 6840 2379 6896
rect 62 6838 2379 6840
rect 2313 6835 2379 6838
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 12157 5946 12223 5949
rect 12157 5944 15578 5946
rect 12157 5888 12162 5944
rect 12218 5888 15578 5944
rect 12157 5886 15578 5888
rect 12157 5883 12223 5886
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 15518 5432 15578 5886
rect 15518 5342 16000 5432
rect 15520 5312 16000 5342
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 4613 4042 4679 4045
rect 9673 4042 9739 4045
rect 4613 4040 9739 4042
rect 4613 3984 4618 4040
rect 4674 3984 9678 4040
rect 9734 3984 9739 4040
rect 4613 3982 9739 3984
rect 4613 3979 4679 3982
rect 9673 3979 9739 3982
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 3509 3634 3575 3637
rect 10041 3634 10107 3637
rect 3509 3632 10107 3634
rect 3509 3576 3514 3632
rect 3570 3576 10046 3632
rect 10102 3576 10107 3632
rect 3509 3574 10107 3576
rect 3509 3571 3575 3574
rect 10041 3571 10107 3574
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 2589 3090 2655 3093
rect 4613 3090 4679 3093
rect 2589 3088 4679 3090
rect 2589 3032 2594 3088
rect 2650 3032 4618 3088
rect 4674 3032 4679 3088
rect 2589 3030 4679 3032
rect 2589 3027 2655 3030
rect 4613 3027 4679 3030
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 0 2544 480 2576
rect 0 2488 110 2544
rect 166 2488 480 2544
rect 0 2456 480 2488
rect 12341 2410 12407 2413
rect 12341 2408 15578 2410
rect 12341 2352 12346 2408
rect 12402 2352 15578 2408
rect 12341 2350 15578 2352
rect 12341 2347 12407 2350
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 15518 1896 15578 2350
rect 15518 1806 16000 1896
rect 15520 1776 16000 1806
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_8
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_12
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_25
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_36
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_29
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_50
timestamp 1586364061
transform 1 0 5704 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_44
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_48
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _183_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_buf_2  _188_
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_77
timestamp 1586364061
transform 1 0 8188 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_70
timestamp 1586364061
transform 1 0 7544 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_89
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_85
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_94 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_92 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _186_
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _184_
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_104
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_108
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_108
timestamp 1586364061
transform 1 0 11040 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_116
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _180_
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_123 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _181_
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_135
timestamp 1586364061
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_135 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_139
timestamp 1586364061
transform 1 0 13892 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_2_12
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 406 592
use scs8hd_conb_1  _172_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_29
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_43
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_47
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _187_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_108
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_120
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_132
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_8
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_12
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_23
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_41
timestamp 1586364061
transform 1 0 4876 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_76
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_93
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _185_
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_121
timestamp 1586364061
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4692 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_29
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_58
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_82
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_86
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_8  FILLER_4_96
timestamp 1586364061
transform 1 0 9936 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_nor2_4  _074_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_23
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _182_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8280 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_70
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_87
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_102
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_11
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_17
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_21
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_24
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_16
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 774 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_47
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_58
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_75
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_79
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_80
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_90
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_96
timestamp 1586364061
transform 1 0 9936 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_84
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_108
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_97
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_105
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_120
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_117
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_121
timestamp 1586364061
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_11
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_1  _069_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_37
timestamp 1586364061
transform 1 0 4508 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_8_43
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_60
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_114
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_126
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_50
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_66
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_9_82
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_103
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_21
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_24
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_29
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_114
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_126
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_138
timestamp 1586364061
transform 1 0 13800 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_23
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_78
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_90
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_102
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_43
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_47
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_51
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _083_
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_72
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_79
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_87
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_26
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_29
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_37
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_54
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_conb_1  _173_
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_65
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_82
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_71
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_90
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_90
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_96
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_107
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_119
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_132
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_20
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_24
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_28
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_32
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_47
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_80
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_84
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_97
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_120
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_11
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_28
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_49
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_55
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_119
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_131
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_22
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_66
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_99
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_103
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_19
timestamp 1586364061
transform 1 0 2852 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_29
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_38
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_50
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_54
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_18_67
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_73
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_137
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_22
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_29
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_35
timestamp 1586364061
transform 1 0 4324 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_39
timestamp 1586364061
transform 1 0 4692 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_54
timestamp 1586364061
transform 1 0 6072 0 -1 13600
box -38 -48 774 592
use scs8hd_conb_1  _174_
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_65
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_69
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_73
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_73
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_8  _146_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_104
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_115
timestamp 1586364061
transform 1 0 11684 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_127
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_139
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_23
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 6256 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_58
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_78
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_82
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_87
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_91
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_104
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_108
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_143
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_11
timestamp 1586364061
transform 1 0 2116 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_16
timestamp 1586364061
transform 1 0 2576 0 -1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_28
timestamp 1586364061
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__082__C
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_59
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_63
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_78
timestamp 1586364061
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_86
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_115
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_127
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_22_139
timestamp 1586364061
transform 1 0 13892 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_42
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_46
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_88
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_92
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 314 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _175_
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_49
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_or3_4  _082_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_87
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_110
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_123
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_143
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_23
timestamp 1586364061
transform 1 0 3220 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_30
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_49
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_25_55
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_nor3_4  _144_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__144__C
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_95
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_99
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 406 592
use scs8hd_conb_1  _171_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_126
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_25_134
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_137
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_22
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 590 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 4232 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_47
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_43
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_43
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 866 592
use scs8hd_or3_4  _110_
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_62
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_67
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_or3_4  _118_
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 866 592
use scs8hd_nor3_4  _143_
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_79
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use scs8hd_or3_4  _068_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_95
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 866 592
use scs8hd_inv_8  _152_
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_99
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_112
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_116
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 590 592
use scs8hd_decap_4  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 13156 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_129
timestamp 1586364061
transform 1 0 12972 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_133
timestamp 1586364061
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_137
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_145
timestamp 1586364061
transform 1 0 14444 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_11
timestamp 1586364061
transform 1 0 2116 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_16
timestamp 1586364061
transform 1 0 2576 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 4508 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_35
timestamp 1586364061
transform 1 0 4324 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_39
timestamp 1586364061
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_52
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8188 0 -1 17952
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_73
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use scs8hd_or3_4  _099_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__D
timestamp 1586364061
transform 1 0 9292 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_91
timestamp 1586364061
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_119
timestamp 1586364061
transform 1 0 12052 0 -1 17952
box -38 -48 774 592
use scs8hd_or3_4  _153_
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_136
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_144
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 590 592
use scs8hd_decap_3  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 3404 0 1 17952
box -38 -48 866 592
use scs8hd_buf_1  _119_
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_17
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_22
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_55
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_73
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_77
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_81
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_or4_4  _135_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_85
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _067_
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_102
timestamp 1586364061
transform 1 0 10488 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_109
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _101_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_113
timestamp 1586364061
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_117
timestamp 1586364061
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 12880 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_126
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_130
timestamp 1586364061
transform 1 0 13064 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_142
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_4  FILLER_30_12
timestamp 1586364061
transform 1 0 2208 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_16
timestamp 1586364061
transform 1 0 2576 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_40
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 4968 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_59
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_64
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_76
timestamp 1586364061
transform 1 0 8096 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 406 592
use scs8hd_or3_4  _066_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__C
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_87
timestamp 1586364061
transform 1 0 9108 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_119
timestamp 1586364061
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_131
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_143
timestamp 1586364061
transform 1 0 14260 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 2668 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_26
timestamp 1586364061
transform 1 0 3496 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_30
timestamp 1586364061
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5520 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_45
timestamp 1586364061
transform 1 0 5244 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_50
timestamp 1586364061
transform 1 0 5704 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_54
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_58
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 130 592
use scs8hd_or2_4  _100_
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _126_
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_90
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_103
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_107
timestamp 1586364061
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_111
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_115
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_conb_1  _176_
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_37
timestamp 1586364061
transform 1 0 4508 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_41
timestamp 1586364061
transform 1 0 4876 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_45
timestamp 1586364061
transform 1 0 5244 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_59
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_76
timestamp 1586364061
transform 1 0 8096 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 774 592
use scs8hd_or3_4  _127_
timestamp 1586364061
transform 1 0 9844 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_104
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_115
timestamp 1586364061
transform 1 0 11684 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_127
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_32_139
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 4140 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_35
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_48
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_54
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_42
timestamp 1586364061
transform 1 0 4968 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_54
timestamp 1586364061
transform 1 0 6072 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_58
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_72
timestamp 1586364061
transform 1 0 7728 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_75
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_71
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_34_83
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_79
timestamp 1586364061
transform 1 0 8372 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_inv_8  _148_
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 866 592
use scs8hd_or3_4  _154_
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 866 592
use scs8hd_inv_8  _160_
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__C
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_88
timestamp 1586364061
transform 1 0 9200 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_92
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_95
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_89
timestamp 1586364061
transform 1 0 9292 0 -1 21216
box -38 -48 130 592
use scs8hd_or3_4  _167_
timestamp 1586364061
transform 1 0 11224 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_105
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_109
timestamp 1586364061
transform 1 0 11132 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_102
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_106
timestamp 1586364061
transform 1 0 10856 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_116
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_112
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_119
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_120
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 12236 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_123
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_34_135
timestamp 1586364061
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_143
timestamp 1586364061
transform 1 0 14260 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 130 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_30
timestamp 1586364061
transform 1 0 3864 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 5244 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_43
timestamp 1586364061
transform 1 0 5060 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_47
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_or3_4  _157_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_or3_4  _062_
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_71
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_or3_4  _149_
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_92
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_105
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_109
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  _150_
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_113
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_126
timestamp 1586364061
transform 1 0 12696 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_130
timestamp 1586364061
transform 1 0 13064 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_142
timestamp 1586364061
transform 1 0 14168 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4508 0 -1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_36
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_48
timestamp 1586364061
transform 1 0 5520 0 -1 22304
box -38 -48 774 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 7268 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_65
timestamp 1586364061
transform 1 0 7084 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_69
timestamp 1586364061
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_8  _147_
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_73
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 9844 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 22304
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_36_108
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 774 592
use scs8hd_or3_4  _164_
timestamp 1586364061
transform 1 0 11776 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_12  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_137
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_buf_1  _073_
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_19
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_22
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4600 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_30
timestamp 1586364061
transform 1 0 3864 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_34
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_49
timestamp 1586364061
transform 1 0 5612 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 8096 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_78
timestamp 1586364061
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use scs8hd_or3_4  _161_
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 9384 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_88
timestamp 1586364061
transform 1 0 9200 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 10948 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_105
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_109
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_117
timestamp 1586364061
transform 1 0 11868 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_121
timestamp 1586364061
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use scs8hd_buf_1  _063_
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_126
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_137
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_141
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_145
timestamp 1586364061
transform 1 0 14444 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 2944 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 4232 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_29
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_36
timestamp 1586364061
transform 1 0 4416 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_49
timestamp 1586364061
transform 1 0 5612 0 -1 23392
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 23392
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_1  _151_
timestamp 1586364061
transform 1 0 8096 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_72
timestamp 1586364061
transform 1 0 7728 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_79
timestamp 1586364061
transform 1 0 8372 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_83
timestamp 1586364061
transform 1 0 8740 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_1  _158_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 8924 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_87
timestamp 1586364061
transform 1 0 9108 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_91
timestamp 1586364061
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_96
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 10120 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_100
timestamp 1586364061
transform 1 0 10304 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 774 592
use scs8hd_conb_1  _170_
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_128
timestamp 1586364061
transform 1 0 12880 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_38_140
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_19
timestamp 1586364061
transform 1 0 2852 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_19
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 222 592
use scs8hd_buf_1  _079_
timestamp 1586364061
transform 1 0 2944 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 2576 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_23
timestamp 1586364061
transform 1 0 3220 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_23
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 866 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_36
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_40
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_29
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_41
timestamp 1586364061
transform 1 0 4876 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_1  _071_
timestamp 1586364061
transform 1 0 5980 0 -1 24480
box -38 -48 314 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 5152 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 5520 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_46
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_50
timestamp 1586364061
transform 1 0 5704 0 -1 24480
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_60
timestamp 1586364061
transform 1 0 6624 0 -1 24480
box -38 -48 222 592
use scs8hd_buf_1  _168_
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_73
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_77
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_73
timestamp 1586364061
transform 1 0 7820 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_88
timestamp 1586364061
transform 1 0 9200 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_90
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 9568 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_96
timestamp 1586364061
transform 1 0 9936 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_94
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use scs8hd_buf_1  _162_
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 314 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 10120 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_107
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_100
timestamp 1586364061
transform 1 0 10304 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_104
timestamp 1586364061
transform 1 0 10672 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_121
timestamp 1586364061
transform 1 0 12236 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12052 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_127
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_128
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_39_139
timestamp 1586364061
transform 1 0 13892 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_145
timestamp 1586364061
transform 1 0 14444 0 1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_140
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_41_11
timestamp 1586364061
transform 1 0 2116 0 1 24480
box -38 -48 314 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 2392 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 2760 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_16
timestamp 1586364061
transform 1 0 2576 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_20
timestamp 1586364061
transform 1 0 2944 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_24
timestamp 1586364061
transform 1 0 3312 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4876 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_36
timestamp 1586364061
transform 1 0 4416 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_40
timestamp 1586364061
transform 1 0 4784 0 1 24480
box -38 -48 130 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_43
timestamp 1586364061
transform 1 0 5060 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_53
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_78
timestamp 1586364061
transform 1 0 8280 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_92
timestamp 1586364061
transform 1 0 9568 0 1 24480
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10488 0 1 24480
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 222 592
use scs8hd_nor2_4  _163_
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_113
timestamp 1586364061
transform 1 0 11500 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_132
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_137
timestamp 1586364061
transform 1 0 13708 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_41_145
timestamp 1586364061
transform 1 0 14444 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  FILLER_42_11
timestamp 1586364061
transform 1 0 2116 0 -1 25568
box -38 -48 314 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 2392 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_8  FILLER_42_23
timestamp 1586364061
transform 1 0 3220 0 -1 25568
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 25568
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4232 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_36
timestamp 1586364061
transform 1 0 4416 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_42_52
timestamp 1586364061
transform 1 0 5888 0 -1 25568
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_58
timestamp 1586364061
transform 1 0 6440 0 -1 25568
box -38 -48 130 592
use scs8hd_conb_1  _177_
timestamp 1586364061
transform 1 0 8464 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_72
timestamp 1586364061
transform 1 0 7728 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_76
timestamp 1586364061
transform 1 0 8096 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_83
timestamp 1586364061
transform 1 0 8740 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_91
timestamp 1586364061
transform 1 0 9476 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 25568
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_42_108
timestamp 1586364061
transform 1 0 11040 0 -1 25568
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11776 0 -1 25568
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_127
timestamp 1586364061
transform 1 0 12788 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_131
timestamp 1586364061
transform 1 0 13156 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_8  FILLER_42_138
timestamp 1586364061
transform 1 0 13800 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4232 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_30
timestamp 1586364061
transform 1 0 3864 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6072 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_45
timestamp 1586364061
transform 1 0 5244 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_49
timestamp 1586364061
transform 1 0 5612 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_53
timestamp 1586364061
transform 1 0 5980 0 1 25568
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 7360 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_56
timestamp 1586364061
transform 1 0 6256 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_60
timestamp 1586364061
transform 1 0 6624 0 1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_43_65
timestamp 1586364061
transform 1 0 7084 0 1 25568
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8280 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 7728 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_70
timestamp 1586364061
transform 1 0 7544 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_74
timestamp 1586364061
transform 1 0 7912 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_89
timestamp 1586364061
transform 1 0 9292 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_93
timestamp 1586364061
transform 1 0 9660 0 1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10028 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_108
timestamp 1586364061
transform 1 0 11040 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 12144 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_112
timestamp 1586364061
transform 1 0 11408 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_116
timestamp 1586364061
transform 1 0 11776 0 1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 13432 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_132
timestamp 1586364061
transform 1 0 13248 0 1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_43_136
timestamp 1586364061
transform 1 0 13616 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_144
timestamp 1586364061
transform 1 0 14352 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4324 0 -1 26656
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6072 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_46
timestamp 1586364061
transform 1 0 5336 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_50
timestamp 1586364061
transform 1 0 5704 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_63
timestamp 1586364061
transform 1 0 6900 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_67
timestamp 1586364061
transform 1 0 7268 0 -1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _064_
timestamp 1586364061
transform 1 0 7820 0 -1 26656
box -38 -48 866 592
use scs8hd_fill_2  FILLER_44_71
timestamp 1586364061
transform 1 0 7636 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_82
timestamp 1586364061
transform 1 0 8648 0 -1 26656
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_88
timestamp 1586364061
transform 1 0 9200 0 -1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_102
timestamp 1586364061
transform 1 0 10488 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_106
timestamp 1586364061
transform 1 0 10856 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_119
timestamp 1586364061
transform 1 0 12052 0 -1 26656
box -38 -48 406 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 12788 0 -1 26656
box -38 -48 866 592
use scs8hd_fill_2  FILLER_44_125
timestamp 1586364061
transform 1 0 12604 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_136
timestamp 1586364061
transform 1 0 13616 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_44_144
timestamp 1586364061
transform 1 0 14352 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3036 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3496 0 1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 590 592
use scs8hd_fill_2  FILLER_45_24
timestamp 1586364061
transform 1 0 3312 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_28
timestamp 1586364061
transform 1 0 3680 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_35
timestamp 1586364061
transform 1 0 4324 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_52
timestamp 1586364061
transform 1 0 5888 0 1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_57
timestamp 1586364061
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_71
timestamp 1586364061
transform 1 0 7636 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_75
timestamp 1586364061
transform 1 0 8004 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_82
timestamp 1586364061
transform 1 0 8648 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_86
timestamp 1586364061
transform 1 0 9016 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_90
timestamp 1586364061
transform 1 0 9384 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_101
timestamp 1586364061
transform 1 0 10396 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_105
timestamp 1586364061
transform 1 0 10764 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11960 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_112
timestamp 1586364061
transform 1 0 11408 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_116
timestamp 1586364061
transform 1 0 11776 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_120
timestamp 1586364061
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_126
timestamp 1586364061
transform 1 0 12696 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_130
timestamp 1586364061
transform 1 0 13064 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_137
timestamp 1586364061
transform 1 0 13708 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_141
timestamp 1586364061
transform 1 0 14076 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_145
timestamp 1586364061
transform 1 0 14444 0 1 26656
box -38 -48 130 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_47_27
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3956 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_34
timestamp 1586364061
transform 1 0 4232 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_38
timestamp 1586364061
transform 1 0 4600 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_37
timestamp 1586364061
transform 1 0 4508 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_41
timestamp 1586364061
transform 1 0 4876 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4784 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 27744
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 27744
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 6072 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_54
timestamp 1586364061
transform 1 0 6072 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_51
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 27744
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 6256 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6624 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_58
timestamp 1586364061
transform 1 0 6440 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_56
timestamp 1586364061
transform 1 0 6256 0 1 27744
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 8740 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_71
timestamp 1586364061
transform 1 0 7636 0 -1 27744
box -38 -48 774 592
use scs8hd_decap_6  FILLER_46_82
timestamp 1586364061
transform 1 0 8648 0 -1 27744
box -38 -48 590 592
use scs8hd_fill_2  FILLER_47_73
timestamp 1586364061
transform 1 0 7820 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_77
timestamp 1586364061
transform 1 0 8188 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_81
timestamp 1586364061
transform 1 0 8556 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 9292 0 1 27744
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 9108 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 9292 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_88
timestamp 1586364061
transform 1 0 9200 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_1  FILLER_46_91
timestamp 1586364061
transform 1 0 9476 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_85
timestamp 1586364061
transform 1 0 8924 0 1 27744
box -38 -48 222 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 10856 0 1 27744
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 27744
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 10304 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_102
timestamp 1586364061
transform 1 0 10488 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_98
timestamp 1586364061
transform 1 0 10120 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_47_102
timestamp 1586364061
transform 1 0 10488 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_109
timestamp 1586364061
transform 1 0 11132 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 11316 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 11684 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_119
timestamp 1586364061
transform 1 0 12052 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_113
timestamp 1586364061
transform 1 0 11500 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_47_117
timestamp 1586364061
transform 1 0 11868 0 1 27744
box -38 -48 406 592
use scs8hd_fill_1  FILLER_47_121
timestamp 1586364061
transform 1 0 12236 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_130
timestamp 1586364061
transform 1 0 13064 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_135
timestamp 1586364061
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use scs8hd_decap_4  FILLER_46_142
timestamp 1586364061
transform 1 0 14168 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_3  FILLER_47_143
timestamp 1586364061
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 774 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 6072 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_43
timestamp 1586364061
transform 1 0 5060 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_47
timestamp 1586364061
transform 1 0 5428 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_51
timestamp 1586364061
transform 1 0 5796 0 -1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 7084 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_63
timestamp 1586364061
transform 1 0 6900 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_67
timestamp 1586364061
transform 1 0 7268 0 -1 28832
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 28832
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_48_82
timestamp 1586364061
transform 1 0 8648 0 -1 28832
box -38 -48 222 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 8832 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_48_86
timestamp 1586364061
transform 1 0 9016 0 -1 28832
box -38 -48 590 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 11224 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_8  FILLER_48_102
timestamp 1586364061
transform 1 0 10488 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_12  FILLER_48_113
timestamp 1586364061
transform 1 0 11500 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_125
timestamp 1586364061
transform 1 0 12604 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_48_137
timestamp 1586364061
transform 1 0 13708 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_1  FILLER_48_145
timestamp 1586364061
transform 1 0 14444 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_49_39
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_53
timestamp 1586364061
transform 1 0 5980 0 1 28832
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7360 0 1 28832
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 6440 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_57
timestamp 1586364061
transform 1 0 6348 0 1 28832
box -38 -48 130 592
use scs8hd_fill_1  FILLER_49_60
timestamp 1586364061
transform 1 0 6624 0 1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_49_62
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 8556 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_79
timestamp 1586364061
transform 1 0 8372 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_83
timestamp 1586364061
transform 1 0 8740 0 1 28832
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9108 0 1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 28832
box -38 -48 222 592
use scs8hd_conb_1  _178_
timestamp 1586364061
transform 1 0 10856 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_98
timestamp 1586364061
transform 1 0 10120 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_102
timestamp 1586364061
transform 1 0 10488 0 1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_49_109
timestamp 1586364061
transform 1 0 11132 0 1 28832
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_115
timestamp 1586364061
transform 1 0 11684 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_118
timestamp 1586364061
transform 1 0 11960 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_135
timestamp 1586364061
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_143
timestamp 1586364061
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_50_46
timestamp 1586364061
transform 1 0 5336 0 -1 29920
box -38 -48 1142 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 6440 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 7452 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_67
timestamp 1586364061
transform 1 0 7268 0 -1 29920
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 8004 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_71
timestamp 1586364061
transform 1 0 7636 0 -1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_50_84
timestamp 1586364061
transform 1 0 8832 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_50_89
timestamp 1586364061
transform 1 0 9292 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 29920
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_50_108
timestamp 1586364061
transform 1 0 11040 0 -1 29920
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 29920
box -38 -48 866 592
use scs8hd_decap_12  FILLER_50_125
timestamp 1586364061
transform 1 0 12604 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_50_137
timestamp 1586364061
transform 1 0 13708 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_50_145
timestamp 1586364061
transform 1 0 14444 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_39
timestamp 1586364061
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_51
timestamp 1586364061
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 7268 0 1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 7084 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_59
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8648 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_76
timestamp 1586364061
transform 1 0 8096 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_80
timestamp 1586364061
transform 1 0 8464 0 1 29920
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9844 0 1 29920
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8832 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_87
timestamp 1586364061
transform 1 0 9108 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_91
timestamp 1586364061
transform 1 0 9476 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_106
timestamp 1586364061
transform 1 0 10856 0 1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_112
timestamp 1586364061
transform 1 0 11408 0 1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_51_116
timestamp 1586364061
transform 1 0 11776 0 1 29920
box -38 -48 590 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_143
timestamp 1586364061
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 6072 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 5704 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_53_47
timestamp 1586364061
transform 1 0 5428 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_52
timestamp 1586364061
transform 1 0 5888 0 1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 866 592
use scs8hd_conb_1  _179_
timestamp 1586364061
transform 1 0 6992 0 -1 31008
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 6808 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 590 592
use scs8hd_decap_4  FILLER_52_67
timestamp 1586364061
transform 1 0 7268 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_3  FILLER_53_56
timestamp 1586364061
transform 1 0 6256 0 1 31008
box -38 -48 314 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 8648 0 1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 8464 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 7820 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 7636 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_73
timestamp 1586364061
transform 1 0 7820 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_71
timestamp 1586364061
transform 1 0 7636 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_75
timestamp 1586364061
transform 1 0 8004 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_79
timestamp 1586364061
transform 1 0 8372 0 1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 9660 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_84
timestamp 1586364061
transform 1 0 8832 0 -1 31008
box -38 -48 590 592
use scs8hd_fill_2  FILLER_53_91
timestamp 1586364061
transform 1 0 9476 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_95
timestamp 1586364061
transform 1 0 9844 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 10028 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_102
timestamp 1586364061
transform 1 0 10488 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_106
timestamp 1586364061
transform 1 0 10856 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_99
timestamp 1586364061
transform 1 0 10212 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_119
timestamp 1586364061
transform 1 0 12052 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_112
timestamp 1586364061
transform 1 0 11408 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_53_116
timestamp 1586364061
transform 1 0 11776 0 1 31008
box -38 -48 590 592
use scs8hd_decap_12  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_131
timestamp 1586364061
transform 1 0 13156 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_135
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  FILLER_52_143
timestamp 1586364061
transform 1 0 14260 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  FILLER_53_143
timestamp 1586364061
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 6072 0 -1 32096
box -38 -48 866 592
use scs8hd_decap_8  FILLER_54_44
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 774 592
use scs8hd_fill_2  FILLER_54_52
timestamp 1586364061
transform 1 0 5888 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_63
timestamp 1586364061
transform 1 0 6900 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_67
timestamp 1586364061
transform 1 0 7268 0 -1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 7636 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 8648 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_80
timestamp 1586364061
transform 1 0 8464 0 -1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_84
timestamp 1586364061
transform 1 0 8832 0 -1 32096
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 10672 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_102
timestamp 1586364061
transform 1 0 10488 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_106
timestamp 1586364061
transform 1 0 10856 0 -1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_113
timestamp 1586364061
transform 1 0 11500 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_54_117
timestamp 1586364061
transform 1 0 11868 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_129
timestamp 1586364061
transform 1 0 12972 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_4  FILLER_54_141
timestamp 1586364061
transform 1 0 14076 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_145
timestamp 1586364061
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_39
timestamp 1586364061
transform 1 0 4692 0 1 32096
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_47
timestamp 1586364061
transform 1 0 5428 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_52
timestamp 1586364061
transform 1 0 5888 0 1 32096
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_57
timestamp 1586364061
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8556 0 1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_73
timestamp 1586364061
transform 1 0 7820 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_77
timestamp 1586364061
transform 1 0 8188 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_92
timestamp 1586364061
transform 1 0 9568 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_96
timestamp 1586364061
transform 1 0 9936 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 10304 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 10120 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_109
timestamp 1586364061
transform 1 0 11132 0 1 32096
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_113
timestamp 1586364061
transform 1 0 11500 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_117
timestamp 1586364061
transform 1 0 11868 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_126
timestamp 1586364061
transform 1 0 12696 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_131
timestamp 1586364061
transform 1 0 13156 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_143
timestamp 1586364061
transform 1 0 14260 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 -1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_44
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 590 592
use scs8hd_fill_2  FILLER_56_53
timestamp 1586364061
transform 1 0 5980 0 -1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 33184
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_56_57
timestamp 1586364061
transform 1 0 6348 0 -1 33184
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_72
timestamp 1586364061
transform 1 0 7728 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_76
timestamp 1586364061
transform 1 0 8096 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_83
timestamp 1586364061
transform 1 0 8740 0 -1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_87
timestamp 1586364061
transform 1 0 9108 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_91
timestamp 1586364061
transform 1 0 9476 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_104
timestamp 1586364061
transform 1 0 10672 0 -1 33184
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_121
timestamp 1586364061
transform 1 0 12236 0 -1 33184
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12972 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_4  FILLER_56_125
timestamp 1586364061
transform 1 0 12604 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_132
timestamp 1586364061
transform 1 0 13248 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_56_144
timestamp 1586364061
transform 1 0 14352 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 33184
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_42
timestamp 1586364061
transform 1 0 4968 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_46
timestamp 1586364061
transform 1 0 5336 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_53
timestamp 1586364061
transform 1 0 5980 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_57
timestamp 1586364061
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_57_66
timestamp 1586364061
transform 1 0 7176 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_78
timestamp 1586364061
transform 1 0 8280 0 1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_57_82
timestamp 1586364061
transform 1 0 8648 0 1 33184
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9292 0 1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_85
timestamp 1586364061
transform 1 0 8924 0 1 33184
box -38 -48 222 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 11040 0 1 33184
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10488 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_100
timestamp 1586364061
transform 1 0 10304 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_104
timestamp 1586364061
transform 1 0 10672 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 11592 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_112
timestamp 1586364061
transform 1 0 11408 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_116
timestamp 1586364061
transform 1 0 11776 0 1 33184
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 13432 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_132
timestamp 1586364061
transform 1 0 13248 0 1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_57_136
timestamp 1586364061
transform 1 0 13616 0 1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_144
timestamp 1586364061
transform 1 0 14352 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 34272
box -38 -48 866 592
use scs8hd_decap_8  FILLER_58_47
timestamp 1586364061
transform 1 0 5428 0 -1 34272
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_64
timestamp 1586364061
transform 1 0 6992 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 34272
box -38 -48 866 592
use scs8hd_fill_1  FILLER_58_71
timestamp 1586364061
transform 1 0 7636 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_58_81
timestamp 1586364061
transform 1 0 8556 0 -1 34272
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  FILLER_58_89
timestamp 1586364061
transform 1 0 9292 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_104
timestamp 1586364061
transform 1 0 10672 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_108
timestamp 1586364061
transform 1 0 11040 0 -1 34272
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 34272
box -38 -48 866 592
use scs8hd_decap_8  FILLER_58_121
timestamp 1586364061
transform 1 0 12236 0 -1 34272
box -38 -48 774 592
use scs8hd_buf_2  _189_
timestamp 1586364061
transform 1 0 12972 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_133
timestamp 1586364061
transform 1 0 13340 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_58_145
timestamp 1586364061
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_59_39
timestamp 1586364061
transform 1 0 4692 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 5612 0 1 34272
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5888 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 6164 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_47
timestamp 1586364061
transform 1 0 5428 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_53
timestamp 1586364061
transform 1 0 5980 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_8  FILLER_60_55
timestamp 1586364061
transform 1 0 6164 0 -1 35360
box -38 -48 774 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 6900 0 -1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 6992 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_57
timestamp 1586364061
transform 1 0 6348 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_66
timestamp 1586364061
transform 1 0 7176 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_60_67
timestamp 1586364061
transform 1 0 7268 0 -1 35360
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 34272
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_79
timestamp 1586364061
transform 1 0 8372 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_83
timestamp 1586364061
transform 1 0 8740 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_60_72
timestamp 1586364061
transform 1 0 7728 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_4  FILLER_60_88
timestamp 1586364061
transform 1 0 9200 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_60_84
timestamp 1586364061
transform 1 0 8832 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 1 34272
box -38 -48 222 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 9108 0 1 34272
box -38 -48 406 592
use scs8hd_decap_6  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 590 592
use scs8hd_fill_2  FILLER_59_95
timestamp 1586364061
transform 1 0 9844 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_91
timestamp 1586364061
transform 1 0 9476 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 9660 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 34272
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_108
timestamp 1586364061
transform 1 0 11040 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_110
timestamp 1586364061
transform 1 0 11224 0 -1 35360
box -38 -48 774 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11960 0 -1 35360
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_59_112
timestamp 1586364061
transform 1 0 11408 0 1 34272
box -38 -48 590 592
use scs8hd_fill_2  FILLER_59_120
timestamp 1586364061
transform 1 0 12144 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_121
timestamp 1586364061
transform 1 0 12236 0 -1 35360
box -38 -48 774 592
use scs8hd_buf_2  _190_
timestamp 1586364061
transform 1 0 12972 0 -1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 12972 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 13340 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_127
timestamp 1586364061
transform 1 0 12788 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_131
timestamp 1586364061
transform 1 0 13156 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_59_135
timestamp 1586364061
transform 1 0 13524 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_133
timestamp 1586364061
transform 1 0 13340 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_59_143
timestamp 1586364061
transform 1 0 14260 0 1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_60_145
timestamp 1586364061
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_buf_2  _191_
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 7360 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_66
timestamp 1586364061
transform 1 0 7176 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_70
timestamp 1586364061
transform 1 0 7544 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 9200 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_86
timestamp 1586364061
transform 1 0 9016 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_90
timestamp 1586364061
transform 1 0 9384 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_95
timestamp 1586364061
transform 1 0 9844 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_108
timestamp 1586364061
transform 1 0 11040 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_120
timestamp 1586364061
transform 1 0 12144 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_135
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_143
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7452 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 130 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_72
timestamp 1586364061
transform 1 0 7728 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_76
timestamp 1586364061
transform 1 0 8096 0 -1 36448
box -38 -48 130 592
use scs8hd_fill_1  FILLER_62_79
timestamp 1586364061
transform 1 0 8372 0 -1 36448
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_62_84
timestamp 1586364061
transform 1 0 8832 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_3  FILLER_62_96
timestamp 1586364061
transform 1 0 9936 0 -1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_62_101
timestamp 1586364061
transform 1 0 10396 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_113
timestamp 1586364061
transform 1 0 11500 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_125
timestamp 1586364061
transform 1 0 12604 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_62_137
timestamp 1586364061
transform 1 0 13708 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_1  FILLER_62_145
timestamp 1586364061
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 36448
box -38 -48 314 592
use scs8hd_decap_6  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 590 592
use scs8hd_fill_2  FILLER_63_95
timestamp 1586364061
transform 1 0 9844 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_99
timestamp 1586364061
transform 1 0 10212 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_63_111
timestamp 1586364061
transform 1 0 11316 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  FILLER_63_119
timestamp 1586364061
transform 1 0 12052 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_143
timestamp 1586364061
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_75
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_87
timestamp 1586364061
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal3 s 15520 5312 16000 5432 6 address[0]
port 0 nsew default input
rlabel metal3 s 15520 8984 16000 9104 6 address[1]
port 1 nsew default input
rlabel metal3 s 15520 12656 16000 12776 6 address[2]
port 2 nsew default input
rlabel metal3 s 15520 16192 16000 16312 6 address[3]
port 3 nsew default input
rlabel metal3 s 15520 19864 16000 19984 6 address[4]
port 4 nsew default input
rlabel metal3 s 15520 23536 16000 23656 6 address[5]
port 5 nsew default input
rlabel metal3 s 15520 27208 16000 27328 6 address[6]
port 6 nsew default input
rlabel metal2 s 386 0 442 480 6 chany_bottom_in[0]
port 7 nsew default input
rlabel metal2 s 1214 0 1270 480 6 chany_bottom_in[1]
port 8 nsew default input
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_in[2]
port 9 nsew default input
rlabel metal2 s 3054 0 3110 480 6 chany_bottom_in[3]
port 10 nsew default input
rlabel metal2 s 3882 0 3938 480 6 chany_bottom_in[4]
port 11 nsew default input
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[5]
port 12 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[6]
port 13 nsew default input
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[7]
port 14 nsew default input
rlabel metal2 s 7470 0 7526 480 6 chany_bottom_in[8]
port 15 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_out[0]
port 16 nsew default tristate
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_out[1]
port 17 nsew default tristate
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_out[2]
port 18 nsew default tristate
rlabel metal2 s 11058 0 11114 480 6 chany_bottom_out[3]
port 19 nsew default tristate
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_out[4]
port 20 nsew default tristate
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_out[5]
port 21 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_out[6]
port 22 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[7]
port 23 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[8]
port 24 nsew default tristate
rlabel metal2 s 386 39520 442 40000 6 chany_top_in[0]
port 25 nsew default input
rlabel metal2 s 1214 39520 1270 40000 6 chany_top_in[1]
port 26 nsew default input
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_in[2]
port 27 nsew default input
rlabel metal2 s 3054 39520 3110 40000 6 chany_top_in[3]
port 28 nsew default input
rlabel metal2 s 3882 39520 3938 40000 6 chany_top_in[4]
port 29 nsew default input
rlabel metal2 s 4802 39520 4858 40000 6 chany_top_in[5]
port 30 nsew default input
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_in[6]
port 31 nsew default input
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_in[7]
port 32 nsew default input
rlabel metal2 s 7470 39520 7526 40000 6 chany_top_in[8]
port 33 nsew default input
rlabel metal2 s 8390 39520 8446 40000 6 chany_top_out[0]
port 34 nsew default tristate
rlabel metal2 s 9218 39520 9274 40000 6 chany_top_out[1]
port 35 nsew default tristate
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_out[2]
port 36 nsew default tristate
rlabel metal2 s 11058 39520 11114 40000 6 chany_top_out[3]
port 37 nsew default tristate
rlabel metal2 s 11886 39520 11942 40000 6 chany_top_out[4]
port 38 nsew default tristate
rlabel metal2 s 12806 39520 12862 40000 6 chany_top_out[5]
port 39 nsew default tristate
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_out[6]
port 40 nsew default tristate
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_out[7]
port 41 nsew default tristate
rlabel metal2 s 15474 39520 15530 40000 6 chany_top_out[8]
port 42 nsew default tristate
rlabel metal3 s 15520 30744 16000 30864 6 data_in
port 43 nsew default input
rlabel metal3 s 15520 1776 16000 1896 6 enable
port 44 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_grid_pin_0_
port 45 nsew default tristate
rlabel metal3 s 0 27344 480 27464 6 left_grid_pin_10_
port 46 nsew default tristate
rlabel metal3 s 0 32376 480 32496 6 left_grid_pin_12_
port 47 nsew default tristate
rlabel metal3 s 0 37408 480 37528 6 left_grid_pin_14_
port 48 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 left_grid_pin_2_
port 49 nsew default tristate
rlabel metal3 s 0 12384 480 12504 6 left_grid_pin_4_
port 50 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 left_grid_pin_6_
port 51 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 left_grid_pin_8_
port 52 nsew default tristate
rlabel metal3 s 15520 34416 16000 34536 6 right_grid_pin_3_
port 53 nsew default tristate
rlabel metal3 s 15520 38088 16000 38208 6 right_grid_pin_7_
port 54 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 vpwr
port 55 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 vgnd
port 56 nsew default input
<< end >>
