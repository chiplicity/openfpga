VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_2__1_
  CLASS BLOCK ;
  FOREIGN cby_2__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 85.000 BY 100.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 96.000 1.290 100.000 ;
    END
  END IO_ISOL_N
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 81.000 9.560 85.000 10.160 ;
    END
  END ccff_tail
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 96.000 43.610 100.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 96.000 63.850 100.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 96.000 65.690 100.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.710 96.000 67.990 100.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 96.000 69.830 100.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 96.000 72.130 100.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 96.000 73.970 100.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 96.000 75.810 100.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.830 96.000 78.110 100.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.670 96.000 79.950 100.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.970 96.000 82.250 100.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 96.000 45.450 100.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.470 96.000 47.750 100.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.310 96.000 49.590 100.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.610 96.000 51.890 100.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 96.000 53.730 100.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 96.000 55.570 100.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.590 96.000 57.870 100.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 96.000 59.710 100.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 96.000 62.010 100.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 96.000 3.130 100.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.090 96.000 23.370 100.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 96.000 25.210 100.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.230 96.000 27.510 100.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.070 96.000 29.350 100.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 31.370 96.000 31.650 100.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.210 96.000 33.490 100.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.050 96.000 35.330 100.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.350 96.000 37.630 100.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.190 96.000 39.470 100.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.490 96.000 41.770 100.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.690 96.000 4.970 100.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.990 96.000 7.270 100.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.830 96.000 9.110 100.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.130 96.000 11.410 100.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.970 96.000 13.250 100.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.810 96.000 15.090 100.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.110 96.000 17.390 100.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.950 96.000 19.230 100.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 21.250 96.000 21.530 100.000 ;
    END
  END chany_top_out[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 81.000 49.000 85.000 49.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 81.000 69.400 85.000 70.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 81.000 89.120 85.000 89.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
  PIN left_grid_pin_16_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END left_grid_pin_16_
  PIN left_grid_pin_17_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END left_grid_pin_17_
  PIN left_grid_pin_18_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END left_grid_pin_18_
  PIN left_grid_pin_19_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END left_grid_pin_19_
  PIN left_grid_pin_20_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END left_grid_pin_20_
  PIN left_grid_pin_21_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END left_grid_pin_21_
  PIN left_grid_pin_22_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END left_grid_pin_22_
  PIN left_grid_pin_23_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END left_grid_pin_23_
  PIN left_grid_pin_24_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END left_grid_pin_24_
  PIN left_grid_pin_25_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END left_grid_pin_25_
  PIN left_grid_pin_26_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END left_grid_pin_26_
  PIN left_grid_pin_27_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END left_grid_pin_27_
  PIN left_grid_pin_28_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END left_grid_pin_28_
  PIN left_grid_pin_29_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END left_grid_pin_29_
  PIN left_grid_pin_30_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END left_grid_pin_30_
  PIN left_grid_pin_31_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END left_grid_pin_31_
  PIN left_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END left_width_0_height_0__pin_0_
  PIN left_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END left_width_0_height_0__pin_1_lower
  PIN left_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END left_width_0_height_0__pin_1_upper
  PIN prog_clk_0_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 96.000 84.090 100.000 ;
    END
  END prog_clk_0_N_out
  PIN prog_clk_0_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END prog_clk_0_S_out
  PIN prog_clk_0_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END prog_clk_0_W_in
  PIN right_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 81.000 29.280 85.000 29.880 ;
    END
  END right_grid_pin_0_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.045 10.640 18.645 87.280 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 29.375 10.640 30.975 87.280 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 79.120 87.125 ;
      LAYER met1 ;
        RECT 0.990 6.500 84.110 95.840 ;
      LAYER met2 ;
        RECT 1.570 95.720 2.570 97.765 ;
        RECT 3.410 95.720 4.410 97.765 ;
        RECT 5.250 95.720 6.710 97.765 ;
        RECT 7.550 95.720 8.550 97.765 ;
        RECT 9.390 95.720 10.850 97.765 ;
        RECT 11.690 95.720 12.690 97.765 ;
        RECT 13.530 95.720 14.530 97.765 ;
        RECT 15.370 95.720 16.830 97.765 ;
        RECT 17.670 95.720 18.670 97.765 ;
        RECT 19.510 95.720 20.970 97.765 ;
        RECT 21.810 95.720 22.810 97.765 ;
        RECT 23.650 95.720 24.650 97.765 ;
        RECT 25.490 95.720 26.950 97.765 ;
        RECT 27.790 95.720 28.790 97.765 ;
        RECT 29.630 95.720 31.090 97.765 ;
        RECT 31.930 95.720 32.930 97.765 ;
        RECT 33.770 95.720 34.770 97.765 ;
        RECT 35.610 95.720 37.070 97.765 ;
        RECT 37.910 95.720 38.910 97.765 ;
        RECT 39.750 95.720 41.210 97.765 ;
        RECT 42.050 95.720 43.050 97.765 ;
        RECT 43.890 95.720 44.890 97.765 ;
        RECT 45.730 95.720 47.190 97.765 ;
        RECT 48.030 95.720 49.030 97.765 ;
        RECT 49.870 95.720 51.330 97.765 ;
        RECT 52.170 95.720 53.170 97.765 ;
        RECT 54.010 95.720 55.010 97.765 ;
        RECT 55.850 95.720 57.310 97.765 ;
        RECT 58.150 95.720 59.150 97.765 ;
        RECT 59.990 95.720 61.450 97.765 ;
        RECT 62.290 95.720 63.290 97.765 ;
        RECT 64.130 95.720 65.130 97.765 ;
        RECT 65.970 95.720 67.430 97.765 ;
        RECT 68.270 95.720 69.270 97.765 ;
        RECT 70.110 95.720 71.570 97.765 ;
        RECT 72.410 95.720 73.410 97.765 ;
        RECT 74.250 95.720 75.250 97.765 ;
        RECT 76.090 95.720 77.550 97.765 ;
        RECT 78.390 95.720 79.390 97.765 ;
        RECT 80.230 95.720 81.690 97.765 ;
        RECT 82.530 95.720 83.530 97.765 ;
        RECT 1.010 4.280 84.080 95.720 ;
        RECT 1.570 4.000 2.570 4.280 ;
        RECT 3.410 4.000 4.870 4.280 ;
        RECT 5.710 4.000 6.710 4.280 ;
        RECT 7.550 4.000 9.010 4.280 ;
        RECT 9.850 4.000 10.850 4.280 ;
        RECT 11.690 4.000 13.150 4.280 ;
        RECT 13.990 4.000 14.990 4.280 ;
        RECT 15.830 4.000 17.290 4.280 ;
        RECT 18.130 4.000 19.130 4.280 ;
        RECT 19.970 4.000 21.430 4.280 ;
        RECT 22.270 4.000 23.270 4.280 ;
        RECT 24.110 4.000 25.570 4.280 ;
        RECT 26.410 4.000 27.410 4.280 ;
        RECT 28.250 4.000 29.710 4.280 ;
        RECT 30.550 4.000 31.550 4.280 ;
        RECT 32.390 4.000 33.850 4.280 ;
        RECT 34.690 4.000 35.690 4.280 ;
        RECT 36.530 4.000 37.990 4.280 ;
        RECT 38.830 4.000 39.830 4.280 ;
        RECT 40.670 4.000 42.130 4.280 ;
        RECT 42.970 4.000 43.970 4.280 ;
        RECT 44.810 4.000 46.270 4.280 ;
        RECT 47.110 4.000 48.110 4.280 ;
        RECT 48.950 4.000 50.410 4.280 ;
        RECT 51.250 4.000 52.250 4.280 ;
        RECT 53.090 4.000 54.550 4.280 ;
        RECT 55.390 4.000 56.390 4.280 ;
        RECT 57.230 4.000 58.690 4.280 ;
        RECT 59.530 4.000 60.530 4.280 ;
        RECT 61.370 4.000 62.830 4.280 ;
        RECT 63.670 4.000 64.670 4.280 ;
        RECT 65.510 4.000 66.970 4.280 ;
        RECT 67.810 4.000 68.810 4.280 ;
        RECT 69.650 4.000 71.110 4.280 ;
        RECT 71.950 4.000 72.950 4.280 ;
        RECT 73.790 4.000 75.250 4.280 ;
        RECT 76.090 4.000 77.090 4.280 ;
        RECT 77.930 4.000 79.390 4.280 ;
        RECT 80.230 4.000 81.230 4.280 ;
        RECT 82.070 4.000 83.530 4.280 ;
      LAYER met3 ;
        RECT 4.400 96.880 81.000 97.745 ;
        RECT 0.985 93.520 81.000 96.880 ;
        RECT 4.400 92.120 81.000 93.520 ;
        RECT 0.985 90.120 81.000 92.120 ;
        RECT 0.985 88.760 80.600 90.120 ;
        RECT 4.400 88.720 80.600 88.760 ;
        RECT 4.400 87.360 81.000 88.720 ;
        RECT 0.985 84.000 81.000 87.360 ;
        RECT 4.400 82.600 81.000 84.000 ;
        RECT 0.985 79.240 81.000 82.600 ;
        RECT 4.400 77.840 81.000 79.240 ;
        RECT 0.985 74.480 81.000 77.840 ;
        RECT 4.400 73.080 81.000 74.480 ;
        RECT 0.985 70.400 81.000 73.080 ;
        RECT 0.985 69.720 80.600 70.400 ;
        RECT 4.400 69.000 80.600 69.720 ;
        RECT 4.400 68.320 81.000 69.000 ;
        RECT 0.985 64.960 81.000 68.320 ;
        RECT 4.400 63.560 81.000 64.960 ;
        RECT 0.985 60.200 81.000 63.560 ;
        RECT 4.400 58.800 81.000 60.200 ;
        RECT 0.985 55.440 81.000 58.800 ;
        RECT 4.400 54.040 81.000 55.440 ;
        RECT 0.985 50.680 81.000 54.040 ;
        RECT 4.400 50.000 81.000 50.680 ;
        RECT 4.400 49.280 80.600 50.000 ;
        RECT 0.985 48.600 80.600 49.280 ;
        RECT 0.985 45.920 81.000 48.600 ;
        RECT 4.400 44.520 81.000 45.920 ;
        RECT 0.985 41.160 81.000 44.520 ;
        RECT 4.400 39.760 81.000 41.160 ;
        RECT 0.985 36.400 81.000 39.760 ;
        RECT 4.400 35.000 81.000 36.400 ;
        RECT 0.985 31.640 81.000 35.000 ;
        RECT 4.400 30.280 81.000 31.640 ;
        RECT 4.400 30.240 80.600 30.280 ;
        RECT 0.985 28.880 80.600 30.240 ;
        RECT 0.985 26.880 81.000 28.880 ;
        RECT 4.400 25.480 81.000 26.880 ;
        RECT 0.985 22.120 81.000 25.480 ;
        RECT 4.400 20.720 81.000 22.120 ;
        RECT 0.985 17.360 81.000 20.720 ;
        RECT 4.400 15.960 81.000 17.360 ;
        RECT 0.985 12.600 81.000 15.960 ;
        RECT 4.400 11.200 81.000 12.600 ;
        RECT 0.985 10.560 81.000 11.200 ;
        RECT 0.985 9.160 80.600 10.560 ;
        RECT 0.985 7.840 81.000 9.160 ;
        RECT 4.400 6.440 81.000 7.840 ;
        RECT 0.985 3.080 81.000 6.440 ;
        RECT 4.400 2.220 81.000 3.080 ;
      LAYER met4 ;
        RECT 14.095 10.240 16.645 87.280 ;
        RECT 19.045 10.240 28.975 87.280 ;
        RECT 31.375 10.240 73.305 87.280 ;
        RECT 14.095 2.215 73.305 10.240 ;
  END
END cby_2__1_
END LIBRARY

