magic
tech sky130A
magscale 1 2
timestamp 1606929242
<< locali >>
rect 9229 17867 9263 17969
rect 10149 17867 10183 17969
rect 9505 13311 9539 13481
rect 12265 10523 12299 10693
rect 12265 2839 12299 3145
<< viali >>
rect 9229 17969 9263 18003
rect 9229 17833 9263 17867
rect 10149 17969 10183 18003
rect 10149 17833 10183 17867
rect 11437 17289 11471 17323
rect 8125 17221 8159 17255
rect 9321 17221 9355 17255
rect 12817 17221 12851 17255
rect 1777 17153 1811 17187
rect 2605 17153 2639 17187
rect 4261 17153 4295 17187
rect 4905 17153 4939 17187
rect 4997 17153 5031 17187
rect 6285 17153 6319 17187
rect 7481 17153 7515 17187
rect 8677 17153 8711 17187
rect 1501 17085 1535 17119
rect 2421 17085 2455 17119
rect 4077 17085 4111 17119
rect 9505 17085 9539 17119
rect 9781 17085 9815 17119
rect 10517 17085 10551 17119
rect 11253 17085 11287 17119
rect 12633 17085 12667 17119
rect 13369 17085 13403 17119
rect 7389 17017 7423 17051
rect 8493 17017 8527 17051
rect 8585 17017 8619 17051
rect 3249 16949 3283 16983
rect 3341 16949 3375 16983
rect 5641 16949 5675 16983
rect 6009 16949 6043 16983
rect 6101 16949 6135 16983
rect 6929 16949 6963 16983
rect 7297 16949 7331 16983
rect 9965 16949 9999 16983
rect 10701 16949 10735 16983
rect 13553 16949 13587 16983
rect 3709 16745 3743 16779
rect 5457 16745 5491 16779
rect 6285 16745 6319 16779
rect 6653 16745 6687 16779
rect 7481 16745 7515 16779
rect 7849 16745 7883 16779
rect 12081 16745 12115 16779
rect 13553 16745 13587 16779
rect 14289 16745 14323 16779
rect 1685 16677 1719 16711
rect 3065 16677 3099 16711
rect 6745 16677 6779 16711
rect 1409 16609 1443 16643
rect 2697 16609 2731 16643
rect 2789 16609 2823 16643
rect 3893 16609 3927 16643
rect 4077 16609 4111 16643
rect 4353 16609 4387 16643
rect 5365 16609 5399 16643
rect 8677 16609 8711 16643
rect 8953 16609 8987 16643
rect 9689 16609 9723 16643
rect 10425 16609 10459 16643
rect 11161 16609 11195 16643
rect 11897 16609 11931 16643
rect 12633 16609 12667 16643
rect 13369 16609 13403 16643
rect 14105 16609 14139 16643
rect 5549 16541 5583 16575
rect 6837 16541 6871 16575
rect 7941 16541 7975 16575
rect 8033 16541 8067 16575
rect 4997 16473 5031 16507
rect 9873 16473 9907 16507
rect 10609 16473 10643 16507
rect 11345 16473 11379 16507
rect 12817 16473 12851 16507
rect 2513 16405 2547 16439
rect 4353 16201 4387 16235
rect 10609 16201 10643 16235
rect 6837 16133 6871 16167
rect 13369 16133 13403 16167
rect 1685 16065 1719 16099
rect 2605 16065 2639 16099
rect 4997 16065 5031 16099
rect 6009 16065 6043 16099
rect 6101 16065 6135 16099
rect 7389 16065 7423 16099
rect 8585 16065 8619 16099
rect 9781 16065 9815 16099
rect 1501 15997 1535 16031
rect 2410 15997 2444 16031
rect 3341 15997 3375 16031
rect 7205 15997 7239 16031
rect 7297 15997 7331 16031
rect 9689 15997 9723 16031
rect 10425 15997 10459 16031
rect 11161 15997 11195 16031
rect 12449 15997 12483 16031
rect 13185 15997 13219 16031
rect 3617 15929 3651 15963
rect 4721 15929 4755 15963
rect 5917 15929 5951 15963
rect 4813 15861 4847 15895
rect 5549 15861 5583 15895
rect 8033 15861 8067 15895
rect 8401 15861 8435 15895
rect 8493 15861 8527 15895
rect 9229 15861 9263 15895
rect 9597 15861 9631 15895
rect 11345 15861 11379 15895
rect 12633 15861 12667 15895
rect 3433 15657 3467 15691
rect 7205 15657 7239 15691
rect 8125 15657 8159 15691
rect 10057 15657 10091 15691
rect 12541 15657 12575 15691
rect 4997 15589 5031 15623
rect 1409 15521 1443 15555
rect 2329 15521 2363 15555
rect 3249 15521 3283 15555
rect 6092 15521 6126 15555
rect 8033 15521 8067 15555
rect 8861 15521 8895 15555
rect 10885 15521 10919 15555
rect 11621 15521 11655 15555
rect 12357 15521 12391 15555
rect 1685 15453 1719 15487
rect 2513 15453 2547 15487
rect 5089 15453 5123 15487
rect 5273 15453 5307 15487
rect 5825 15453 5859 15487
rect 8217 15453 8251 15487
rect 10149 15453 10183 15487
rect 10333 15453 10367 15487
rect 13093 15453 13127 15487
rect 13737 15453 13771 15487
rect 11069 15385 11103 15419
rect 11805 15385 11839 15419
rect 4629 15317 4663 15351
rect 7665 15317 7699 15351
rect 9045 15317 9079 15351
rect 9689 15317 9723 15351
rect 3709 15113 3743 15147
rect 8217 15113 8251 15147
rect 8677 15113 8711 15147
rect 9873 15113 9907 15147
rect 11069 15045 11103 15079
rect 2053 14977 2087 15011
rect 4169 14977 4203 15011
rect 4353 14977 4387 15011
rect 9229 14977 9263 15011
rect 10425 14977 10459 15011
rect 11529 14977 11563 15011
rect 11713 14977 11747 15011
rect 13737 14977 13771 15011
rect 1777 14909 1811 14943
rect 2697 14909 2731 14943
rect 4905 14909 4939 14943
rect 5172 14909 5206 14943
rect 6837 14909 6871 14943
rect 7104 14909 7138 14943
rect 9045 14909 9079 14943
rect 2973 14841 3007 14875
rect 10241 14841 10275 14875
rect 13093 14841 13127 14875
rect 4077 14773 4111 14807
rect 6285 14773 6319 14807
rect 9137 14773 9171 14807
rect 10333 14773 10367 14807
rect 11437 14773 11471 14807
rect 12449 14773 12483 14807
rect 14381 14773 14415 14807
rect 7021 14569 7055 14603
rect 8861 14569 8895 14603
rect 9689 14569 9723 14603
rect 10885 14569 10919 14603
rect 14105 14569 14139 14603
rect 2145 14501 2179 14535
rect 3157 14501 3191 14535
rect 5886 14501 5920 14535
rect 11345 14501 11379 14535
rect 1869 14433 1903 14467
rect 3249 14433 3283 14467
rect 4813 14433 4847 14467
rect 4905 14433 4939 14467
rect 7748 14433 7782 14467
rect 9505 14433 9539 14467
rect 10057 14433 10091 14467
rect 11253 14433 11287 14467
rect 12081 14433 12115 14467
rect 13369 14433 13403 14467
rect 3433 14365 3467 14399
rect 5089 14365 5123 14399
rect 5641 14365 5675 14399
rect 7481 14365 7515 14399
rect 10149 14365 10183 14399
rect 10241 14365 10275 14399
rect 11437 14365 11471 14399
rect 12265 14365 12299 14399
rect 2789 14297 2823 14331
rect 4445 14229 4479 14263
rect 9321 14229 9355 14263
rect 13553 14229 13587 14263
rect 2513 14025 2547 14059
rect 3709 14025 3743 14059
rect 6285 14025 6319 14059
rect 10517 14025 10551 14059
rect 8217 13957 8251 13991
rect 12449 13957 12483 13991
rect 14013 13957 14047 13991
rect 2973 13889 3007 13923
rect 3157 13889 3191 13923
rect 4353 13889 4387 13923
rect 6837 13889 6871 13923
rect 10977 13889 11011 13923
rect 11069 13889 11103 13923
rect 13093 13889 13127 13923
rect 1593 13821 1627 13855
rect 1869 13821 1903 13855
rect 4169 13821 4203 13855
rect 4905 13821 4939 13855
rect 7104 13821 7138 13855
rect 8677 13821 8711 13855
rect 8933 13821 8967 13855
rect 13829 13821 13863 13855
rect 5172 13753 5206 13787
rect 10885 13753 10919 13787
rect 12817 13753 12851 13787
rect 14565 13753 14599 13787
rect 2881 13685 2915 13719
rect 4077 13685 4111 13719
rect 10057 13685 10091 13719
rect 11713 13685 11747 13719
rect 12909 13685 12943 13719
rect 1593 13481 1627 13515
rect 1961 13481 1995 13515
rect 8033 13481 8067 13515
rect 8401 13481 8435 13515
rect 9505 13481 9539 13515
rect 12725 13481 12759 13515
rect 13093 13481 13127 13515
rect 13185 13481 13219 13515
rect 3157 13413 3191 13447
rect 6438 13413 6472 13447
rect 2053 13345 2087 13379
rect 4353 13345 4387 13379
rect 4620 13345 4654 13379
rect 6193 13345 6227 13379
rect 8493 13345 8527 13379
rect 9413 13345 9447 13379
rect 14197 13413 14231 13447
rect 9945 13345 9979 13379
rect 11897 13345 11931 13379
rect 11989 13345 12023 13379
rect 13921 13345 13955 13379
rect 2237 13277 2271 13311
rect 3249 13277 3283 13311
rect 3433 13277 3467 13311
rect 8677 13277 8711 13311
rect 9505 13277 9539 13311
rect 9689 13277 9723 13311
rect 12081 13277 12115 13311
rect 13277 13277 13311 13311
rect 5733 13209 5767 13243
rect 9229 13209 9263 13243
rect 11529 13209 11563 13243
rect 2789 13141 2823 13175
rect 7573 13141 7607 13175
rect 11069 13141 11103 13175
rect 6285 12937 6319 12971
rect 8217 12937 8251 12971
rect 13645 12937 13679 12971
rect 10057 12869 10091 12903
rect 2513 12801 2547 12835
rect 6837 12801 6871 12835
rect 8677 12801 8711 12835
rect 11161 12801 11195 12835
rect 11713 12801 11747 12835
rect 13001 12801 13035 12835
rect 3065 12733 3099 12767
rect 4905 12733 4939 12767
rect 7104 12733 7138 12767
rect 10885 12733 10919 12767
rect 13829 12733 13863 12767
rect 13921 12733 13955 12767
rect 14841 12733 14875 12767
rect 3332 12665 3366 12699
rect 5172 12665 5206 12699
rect 8944 12665 8978 12699
rect 10977 12665 11011 12699
rect 12817 12665 12851 12699
rect 14197 12665 14231 12699
rect 1869 12597 1903 12631
rect 2237 12597 2271 12631
rect 2329 12597 2363 12631
rect 4445 12597 4479 12631
rect 10517 12597 10551 12631
rect 12449 12597 12483 12631
rect 12909 12597 12943 12631
rect 15025 12597 15059 12631
rect 2789 12393 2823 12427
rect 3157 12393 3191 12427
rect 3249 12393 3283 12427
rect 8769 12393 8803 12427
rect 9229 12393 9263 12427
rect 12541 12393 12575 12427
rect 2053 12325 2087 12359
rect 5794 12325 5828 12359
rect 7656 12325 7690 12359
rect 10057 12325 10091 12359
rect 1961 12257 1995 12291
rect 4721 12257 4755 12291
rect 4813 12257 4847 12291
rect 9413 12257 9447 12291
rect 11253 12257 11287 12291
rect 12449 12257 12483 12291
rect 13461 12257 13495 12291
rect 13553 12257 13587 12291
rect 14473 12257 14507 12291
rect 2237 12189 2271 12223
rect 3433 12189 3467 12223
rect 4905 12189 4939 12223
rect 5549 12189 5583 12223
rect 7389 12189 7423 12223
rect 10149 12189 10183 12223
rect 10333 12189 10367 12223
rect 11345 12189 11379 12223
rect 11437 12189 11471 12223
rect 12633 12189 12667 12223
rect 13829 12189 13863 12223
rect 6929 12121 6963 12155
rect 10885 12121 10919 12155
rect 1593 12053 1627 12087
rect 4353 12053 4387 12087
rect 9689 12053 9723 12087
rect 12081 12053 12115 12087
rect 13277 12053 13311 12087
rect 14657 12053 14691 12087
rect 2513 11849 2547 11883
rect 3709 11849 3743 11883
rect 12449 11849 12483 11883
rect 3157 11713 3191 11747
rect 4169 11713 4203 11747
rect 4353 11713 4387 11747
rect 7389 11713 7423 11747
rect 9781 11713 9815 11747
rect 10977 11713 11011 11747
rect 13001 11713 13035 11747
rect 13921 11713 13955 11747
rect 1593 11645 1627 11679
rect 2881 11645 2915 11679
rect 4905 11645 4939 11679
rect 9597 11645 9631 11679
rect 11621 11645 11655 11679
rect 12909 11645 12943 11679
rect 13645 11645 13679 11679
rect 14565 11645 14599 11679
rect 1869 11577 1903 11611
rect 2973 11577 3007 11611
rect 5172 11577 5206 11611
rect 7634 11577 7668 11611
rect 10885 11577 10919 11611
rect 14841 11577 14875 11611
rect 4077 11509 4111 11543
rect 6285 11509 6319 11543
rect 8769 11509 8803 11543
rect 9229 11509 9263 11543
rect 9689 11509 9723 11543
rect 10425 11509 10459 11543
rect 10793 11509 10827 11543
rect 11805 11509 11839 11543
rect 12817 11509 12851 11543
rect 1593 11305 1627 11339
rect 4629 11305 4663 11339
rect 9689 11305 9723 11339
rect 10149 11305 10183 11339
rect 10885 11305 10919 11339
rect 11345 11305 11379 11339
rect 12449 11305 12483 11339
rect 13277 11305 13311 11339
rect 10057 11237 10091 11271
rect 12541 11237 12575 11271
rect 1961 11169 1995 11203
rect 2053 11169 2087 11203
rect 3157 11169 3191 11203
rect 4997 11169 5031 11203
rect 5825 11169 5859 11203
rect 6092 11169 6126 11203
rect 7932 11169 7966 11203
rect 11253 11169 11287 11203
rect 13645 11169 13679 11203
rect 14473 11169 14507 11203
rect 2145 11101 2179 11135
rect 3249 11101 3283 11135
rect 3433 11101 3467 11135
rect 5089 11101 5123 11135
rect 5273 11101 5307 11135
rect 7665 11101 7699 11135
rect 10333 11101 10367 11135
rect 11437 11101 11471 11135
rect 12633 11101 12667 11135
rect 13737 11101 13771 11135
rect 13829 11101 13863 11135
rect 2789 11033 2823 11067
rect 9045 11033 9079 11067
rect 12081 11033 12115 11067
rect 14657 11033 14691 11067
rect 7205 10965 7239 10999
rect 3709 10761 3743 10795
rect 6285 10761 6319 10795
rect 6837 10761 6871 10795
rect 8033 10761 8067 10795
rect 10333 10761 10367 10795
rect 11713 10693 11747 10727
rect 12265 10693 12299 10727
rect 15025 10693 15059 10727
rect 2973 10625 3007 10659
rect 3157 10625 3191 10659
rect 4353 10625 4387 10659
rect 7481 10625 7515 10659
rect 8493 10625 8527 10659
rect 10977 10625 11011 10659
rect 1593 10557 1627 10591
rect 4077 10557 4111 10591
rect 4905 10557 4939 10591
rect 7297 10557 7331 10591
rect 8217 10557 8251 10591
rect 10701 10557 10735 10591
rect 11529 10557 11563 10591
rect 13001 10625 13035 10659
rect 14197 10625 14231 10659
rect 12817 10557 12851 10591
rect 14013 10557 14047 10591
rect 14841 10557 14875 10591
rect 1869 10489 1903 10523
rect 5150 10489 5184 10523
rect 8760 10489 8794 10523
rect 12265 10489 12299 10523
rect 12909 10489 12943 10523
rect 2513 10421 2547 10455
rect 2881 10421 2915 10455
rect 4169 10421 4203 10455
rect 7205 10421 7239 10455
rect 9873 10421 9907 10455
rect 10793 10421 10827 10455
rect 12449 10421 12483 10455
rect 13645 10421 13679 10455
rect 14105 10421 14139 10455
rect 2789 10217 2823 10251
rect 4261 10217 4295 10251
rect 4721 10217 4755 10251
rect 10885 10217 10919 10251
rect 11253 10217 11287 10251
rect 13277 10217 13311 10251
rect 1961 10149 1995 10183
rect 4629 10149 4663 10183
rect 5724 10149 5758 10183
rect 10149 10149 10183 10183
rect 12449 10149 12483 10183
rect 2053 10081 2087 10115
rect 3157 10081 3191 10115
rect 3249 10081 3283 10115
rect 7297 10081 7331 10115
rect 7564 10081 7598 10115
rect 9321 10081 9355 10115
rect 10057 10081 10091 10115
rect 13645 10081 13679 10115
rect 13737 10081 13771 10115
rect 14473 10081 14507 10115
rect 2237 10013 2271 10047
rect 3433 10013 3467 10047
rect 4905 10013 4939 10047
rect 5457 10013 5491 10047
rect 10241 10013 10275 10047
rect 11345 10013 11379 10047
rect 11529 10013 11563 10047
rect 12541 10013 12575 10047
rect 12725 10013 12759 10047
rect 13829 10013 13863 10047
rect 9689 9945 9723 9979
rect 14657 9945 14691 9979
rect 1593 9877 1627 9911
rect 6837 9877 6871 9911
rect 8677 9877 8711 9911
rect 9137 9877 9171 9911
rect 12081 9877 12115 9911
rect 5181 9673 5215 9707
rect 12449 9673 12483 9707
rect 2145 9605 2179 9639
rect 9873 9605 9907 9639
rect 13645 9605 13679 9639
rect 2605 9537 2639 9571
rect 2789 9537 2823 9571
rect 3617 9537 3651 9571
rect 3801 9537 3835 9571
rect 5273 9537 5307 9571
rect 6837 9537 6871 9571
rect 9321 9537 9355 9571
rect 10425 9537 10459 9571
rect 11621 9537 11655 9571
rect 13001 9537 13035 9571
rect 14105 9537 14139 9571
rect 14197 9537 14231 9571
rect 1593 9469 1627 9503
rect 1869 9469 1903 9503
rect 9045 9469 9079 9503
rect 9137 9469 9171 9503
rect 10241 9469 10275 9503
rect 11529 9469 11563 9503
rect 14013 9469 14047 9503
rect 14841 9469 14875 9503
rect 2513 9401 2547 9435
rect 4068 9401 4102 9435
rect 5540 9401 5574 9435
rect 7082 9401 7116 9435
rect 12817 9401 12851 9435
rect 2973 9333 3007 9367
rect 3341 9333 3375 9367
rect 3433 9333 3467 9367
rect 6653 9333 6687 9367
rect 8217 9333 8251 9367
rect 8677 9333 8711 9367
rect 10333 9333 10367 9367
rect 11069 9333 11103 9367
rect 11437 9333 11471 9367
rect 12909 9333 12943 9367
rect 15025 9333 15059 9367
rect 2789 9129 2823 9163
rect 10885 9129 10919 9163
rect 11345 9129 11379 9163
rect 13277 9129 13311 9163
rect 3249 9061 3283 9095
rect 8125 9061 8159 9095
rect 8217 9061 8251 9095
rect 10149 9061 10183 9095
rect 13737 9061 13771 9095
rect 1961 8993 1995 9027
rect 3157 8993 3191 9027
rect 4629 8993 4663 9027
rect 5917 8993 5951 9027
rect 8585 8993 8619 9027
rect 10057 8993 10091 9027
rect 11253 8993 11287 9027
rect 12449 8993 12483 9027
rect 13645 8993 13679 9027
rect 14473 8993 14507 9027
rect 2053 8925 2087 8959
rect 2237 8925 2271 8959
rect 3433 8925 3467 8959
rect 4721 8925 4755 8959
rect 4905 8925 4939 8959
rect 8309 8925 8343 8959
rect 8769 8925 8803 8959
rect 10333 8925 10367 8959
rect 11529 8925 11563 8959
rect 12541 8925 12575 8959
rect 12633 8925 12667 8959
rect 13829 8925 13863 8959
rect 7757 8857 7791 8891
rect 1593 8789 1627 8823
rect 4261 8789 4295 8823
rect 7389 8789 7423 8823
rect 9689 8789 9723 8823
rect 12081 8789 12115 8823
rect 14657 8789 14691 8823
rect 11069 8585 11103 8619
rect 12449 8585 12483 8619
rect 13645 8585 13679 8619
rect 3709 8517 3743 8551
rect 6285 8517 6319 8551
rect 8217 8517 8251 8551
rect 15025 8517 15059 8551
rect 3157 8449 3191 8483
rect 4353 8449 4387 8483
rect 9321 8449 9355 8483
rect 10425 8449 10459 8483
rect 11529 8449 11563 8483
rect 11621 8449 11655 8483
rect 13001 8449 13035 8483
rect 14197 8449 14231 8483
rect 1593 8381 1627 8415
rect 2973 8381 3007 8415
rect 4077 8381 4111 8415
rect 4169 8381 4203 8415
rect 4905 8381 4939 8415
rect 6837 8381 6871 8415
rect 9137 8381 9171 8415
rect 10241 8381 10275 8415
rect 14841 8381 14875 8415
rect 1869 8313 1903 8347
rect 2881 8313 2915 8347
rect 5172 8313 5206 8347
rect 7104 8313 7138 8347
rect 9045 8313 9079 8347
rect 11437 8313 11471 8347
rect 12817 8313 12851 8347
rect 12909 8313 12943 8347
rect 14013 8313 14047 8347
rect 2513 8245 2547 8279
rect 8677 8245 8711 8279
rect 9873 8245 9907 8279
rect 10333 8245 10367 8279
rect 14105 8245 14139 8279
rect 1593 8041 1627 8075
rect 1961 8041 1995 8075
rect 9137 8041 9171 8075
rect 9689 8041 9723 8075
rect 10149 8041 10183 8075
rect 10885 8041 10919 8075
rect 11253 8041 11287 8075
rect 11345 8041 11379 8075
rect 12081 8041 12115 8075
rect 13737 8041 13771 8075
rect 2053 7973 2087 8007
rect 3157 7973 3191 8007
rect 4344 7905 4378 7939
rect 6173 7905 6207 7939
rect 8024 7905 8058 7939
rect 10057 7905 10091 7939
rect 12449 7905 12483 7939
rect 13645 7905 13679 7939
rect 14473 7905 14507 7939
rect 2237 7837 2271 7871
rect 3249 7837 3283 7871
rect 3433 7837 3467 7871
rect 4077 7837 4111 7871
rect 5917 7837 5951 7871
rect 7757 7837 7791 7871
rect 10333 7837 10367 7871
rect 11437 7837 11471 7871
rect 12541 7837 12575 7871
rect 12725 7837 12759 7871
rect 13829 7837 13863 7871
rect 7297 7769 7331 7803
rect 2789 7701 2823 7735
rect 5457 7701 5491 7735
rect 13277 7701 13311 7735
rect 14657 7701 14691 7735
rect 1869 7497 1903 7531
rect 6285 7497 6319 7531
rect 4445 7429 4479 7463
rect 8217 7429 8251 7463
rect 12449 7429 12483 7463
rect 2329 7361 2363 7395
rect 2513 7361 2547 7395
rect 11069 7361 11103 7395
rect 12909 7361 12943 7395
rect 13001 7361 13035 7395
rect 14197 7361 14231 7395
rect 2237 7293 2271 7327
rect 3065 7293 3099 7327
rect 4905 7293 4939 7327
rect 6837 7293 6871 7327
rect 7093 7293 7127 7327
rect 8677 7293 8711 7327
rect 8933 7293 8967 7327
rect 10977 7293 11011 7327
rect 14841 7293 14875 7327
rect 3332 7225 3366 7259
rect 5172 7225 5206 7259
rect 14013 7225 14047 7259
rect 10057 7157 10091 7191
rect 10517 7157 10551 7191
rect 10885 7157 10919 7191
rect 11713 7157 11747 7191
rect 12817 7157 12851 7191
rect 13645 7157 13679 7191
rect 14105 7157 14139 7191
rect 15025 7157 15059 7191
rect 3525 6953 3559 6987
rect 7113 6953 7147 6987
rect 8953 6953 8987 6987
rect 10057 6953 10091 6987
rect 10885 6953 10919 6987
rect 12081 6953 12115 6987
rect 12449 6953 12483 6987
rect 12541 6953 12575 6987
rect 10149 6885 10183 6919
rect 11253 6885 11287 6919
rect 11345 6885 11379 6919
rect 13645 6885 13679 6919
rect 1409 6817 1443 6851
rect 2412 6817 2446 6851
rect 4261 6817 4295 6851
rect 5089 6817 5123 6851
rect 6000 6817 6034 6851
rect 7840 6817 7874 6851
rect 14473 6817 14507 6851
rect 2145 6749 2179 6783
rect 5733 6749 5767 6783
rect 7573 6749 7607 6783
rect 10241 6749 10275 6783
rect 11437 6749 11471 6783
rect 12633 6749 12667 6783
rect 13737 6749 13771 6783
rect 13829 6749 13863 6783
rect 14657 6681 14691 6715
rect 1593 6613 1627 6647
rect 9689 6613 9723 6647
rect 13277 6613 13311 6647
rect 1869 6409 1903 6443
rect 4445 6409 4479 6443
rect 10057 6409 10091 6443
rect 12449 6409 12483 6443
rect 6285 6341 6319 6375
rect 10517 6341 10551 6375
rect 2421 6273 2455 6307
rect 4905 6273 4939 6307
rect 11069 6273 11103 6307
rect 11713 6273 11747 6307
rect 13001 6273 13035 6307
rect 14289 6273 14323 6307
rect 2237 6205 2271 6239
rect 3065 6205 3099 6239
rect 3332 6205 3366 6239
rect 6837 6205 6871 6239
rect 8677 6205 8711 6239
rect 8933 6205 8967 6239
rect 10885 6205 10919 6239
rect 10977 6205 11011 6239
rect 12909 6205 12943 6239
rect 14841 6205 14875 6239
rect 5150 6137 5184 6171
rect 7104 6137 7138 6171
rect 14105 6137 14139 6171
rect 2329 6069 2363 6103
rect 8217 6069 8251 6103
rect 12817 6069 12851 6103
rect 13645 6069 13679 6103
rect 14013 6069 14047 6103
rect 15025 6069 15059 6103
rect 4629 5865 4663 5899
rect 11897 5865 11931 5899
rect 12725 5865 12759 5899
rect 14381 5865 14415 5899
rect 4721 5797 4755 5831
rect 5702 5797 5736 5831
rect 1409 5729 1443 5763
rect 2145 5729 2179 5763
rect 2412 5729 2446 5763
rect 7553 5729 7587 5763
rect 9321 5729 9355 5763
rect 9956 5729 9990 5763
rect 11989 5729 12023 5763
rect 13093 5729 13127 5763
rect 13185 5729 13219 5763
rect 14289 5729 14323 5763
rect 4905 5661 4939 5695
rect 5457 5661 5491 5695
rect 7297 5661 7331 5695
rect 9689 5661 9723 5695
rect 12173 5661 12207 5695
rect 13277 5661 13311 5695
rect 14473 5661 14507 5695
rect 8677 5593 8711 5627
rect 9137 5593 9171 5627
rect 11069 5593 11103 5627
rect 1593 5525 1627 5559
rect 3525 5525 3559 5559
rect 4261 5525 4295 5559
rect 6837 5525 6871 5559
rect 11529 5525 11563 5559
rect 13921 5525 13955 5559
rect 1869 5321 1903 5355
rect 8217 5321 8251 5355
rect 12449 5321 12483 5355
rect 13645 5321 13679 5355
rect 4445 5253 4479 5287
rect 10057 5253 10091 5287
rect 15025 5253 15059 5287
rect 2513 5185 2547 5219
rect 11069 5185 11103 5219
rect 13001 5185 13035 5219
rect 13461 5185 13495 5219
rect 14197 5185 14231 5219
rect 2237 5117 2271 5151
rect 3065 5117 3099 5151
rect 4905 5117 4939 5151
rect 5172 5117 5206 5151
rect 6837 5117 6871 5151
rect 7104 5117 7138 5151
rect 8677 5117 8711 5151
rect 8944 5117 8978 5151
rect 10885 5117 10919 5151
rect 11713 5117 11747 5151
rect 14013 5117 14047 5151
rect 14841 5117 14875 5151
rect 3332 5049 3366 5083
rect 10977 5049 11011 5083
rect 12817 5049 12851 5083
rect 14105 5049 14139 5083
rect 2329 4981 2363 5015
rect 6285 4981 6319 5015
rect 10517 4981 10551 5015
rect 12909 4981 12943 5015
rect 10057 4777 10091 4811
rect 10149 4777 10183 4811
rect 12541 4777 12575 4811
rect 13277 4777 13311 4811
rect 13645 4777 13679 4811
rect 2412 4709 2446 4743
rect 4537 4709 4571 4743
rect 8953 4709 8987 4743
rect 12449 4709 12483 4743
rect 1409 4641 1443 4675
rect 2145 4641 2179 4675
rect 4445 4641 4479 4675
rect 5540 4641 5574 4675
rect 7380 4641 7414 4675
rect 11253 4641 11287 4675
rect 13737 4641 13771 4675
rect 14473 4641 14507 4675
rect 4721 4573 4755 4607
rect 5273 4573 5307 4607
rect 7113 4573 7147 4607
rect 10241 4573 10275 4607
rect 11345 4573 11379 4607
rect 11437 4573 11471 4607
rect 12633 4573 12667 4607
rect 13829 4573 13863 4607
rect 3525 4505 3559 4539
rect 8493 4505 8527 4539
rect 12081 4505 12115 4539
rect 14657 4505 14691 4539
rect 1593 4437 1627 4471
rect 4077 4437 4111 4471
rect 6653 4437 6687 4471
rect 9689 4437 9723 4471
rect 10885 4437 10919 4471
rect 11069 4233 11103 4267
rect 4445 4165 4479 4199
rect 8677 4165 8711 4199
rect 9873 4165 9907 4199
rect 2513 4097 2547 4131
rect 3065 4097 3099 4131
rect 9321 4097 9355 4131
rect 10425 4097 10459 4131
rect 11529 4097 11563 4131
rect 11621 4097 11655 4131
rect 13001 4097 13035 4131
rect 14105 4097 14139 4131
rect 14197 4097 14231 4131
rect 2237 4029 2271 4063
rect 4905 4029 4939 4063
rect 6837 4029 6871 4063
rect 10241 4029 10275 4063
rect 10333 4029 10367 4063
rect 12817 4029 12851 4063
rect 12909 4029 12943 4063
rect 14841 4029 14875 4063
rect 3332 3961 3366 3995
rect 5172 3961 5206 3995
rect 7082 3961 7116 3995
rect 14013 3961 14047 3995
rect 1869 3893 1903 3927
rect 2329 3893 2363 3927
rect 6285 3893 6319 3927
rect 8217 3893 8251 3927
rect 9045 3893 9079 3927
rect 9137 3893 9171 3927
rect 11437 3893 11471 3927
rect 12449 3893 12483 3927
rect 13645 3893 13679 3927
rect 15025 3893 15059 3927
rect 1593 3689 1627 3723
rect 1961 3689 1995 3723
rect 3157 3689 3191 3723
rect 3249 3689 3283 3723
rect 4997 3689 5031 3723
rect 8953 3689 8987 3723
rect 10885 3689 10919 3723
rect 11253 3689 11287 3723
rect 12081 3689 12115 3723
rect 12449 3689 12483 3723
rect 13645 3689 13679 3723
rect 2053 3621 2087 3655
rect 4905 3621 4939 3655
rect 10057 3621 10091 3655
rect 12541 3621 12575 3655
rect 6000 3553 6034 3587
rect 7573 3553 7607 3587
rect 7829 3553 7863 3587
rect 11345 3553 11379 3587
rect 14473 3553 14507 3587
rect 2237 3485 2271 3519
rect 3433 3485 3467 3519
rect 5181 3485 5215 3519
rect 5733 3485 5767 3519
rect 10149 3485 10183 3519
rect 10241 3485 10275 3519
rect 11437 3485 11471 3519
rect 12633 3485 12667 3519
rect 13737 3485 13771 3519
rect 13921 3485 13955 3519
rect 2789 3417 2823 3451
rect 9689 3417 9723 3451
rect 13277 3417 13311 3451
rect 4537 3349 4571 3383
rect 7113 3349 7147 3383
rect 14657 3349 14691 3383
rect 2513 3145 2547 3179
rect 3709 3145 3743 3179
rect 6285 3145 6319 3179
rect 12265 3145 12299 3179
rect 13645 3145 13679 3179
rect 8677 3077 8711 3111
rect 9781 3077 9815 3111
rect 1869 3009 1903 3043
rect 3157 3009 3191 3043
rect 4169 3009 4203 3043
rect 4353 3009 4387 3043
rect 6837 3009 6871 3043
rect 9137 3009 9171 3043
rect 9321 3009 9355 3043
rect 10517 3009 10551 3043
rect 11621 3009 11655 3043
rect 1593 2941 1627 2975
rect 4077 2941 4111 2975
rect 4905 2941 4939 2975
rect 10241 2941 10275 2975
rect 2973 2873 3007 2907
rect 5150 2873 5184 2907
rect 7082 2873 7116 2907
rect 10333 2873 10367 2907
rect 13001 3009 13035 3043
rect 14105 3009 14139 3043
rect 14289 3009 14323 3043
rect 12817 2941 12851 2975
rect 14841 2941 14875 2975
rect 2881 2805 2915 2839
rect 8217 2805 8251 2839
rect 9045 2805 9079 2839
rect 9873 2805 9907 2839
rect 11069 2805 11103 2839
rect 11437 2805 11471 2839
rect 11529 2805 11563 2839
rect 12265 2805 12299 2839
rect 12449 2805 12483 2839
rect 12909 2805 12943 2839
rect 14013 2805 14047 2839
rect 15025 2805 15059 2839
rect 6377 2601 6411 2635
rect 6929 2601 6963 2635
rect 7389 2601 7423 2635
rect 8125 2601 8159 2635
rect 10149 2601 10183 2635
rect 10241 2601 10275 2635
rect 11437 2601 11471 2635
rect 13093 2601 13127 2635
rect 14289 2601 14323 2635
rect 5242 2533 5276 2567
rect 11345 2533 11379 2567
rect 13001 2533 13035 2567
rect 1409 2465 1443 2499
rect 2412 2465 2446 2499
rect 4077 2465 4111 2499
rect 7297 2465 7331 2499
rect 8493 2465 8527 2499
rect 9505 2465 9539 2499
rect 12357 2465 12391 2499
rect 14197 2465 14231 2499
rect 15209 2465 15243 2499
rect 2145 2397 2179 2431
rect 4353 2397 4387 2431
rect 4997 2397 5031 2431
rect 7481 2397 7515 2431
rect 8585 2397 8619 2431
rect 8677 2397 8711 2431
rect 10333 2397 10367 2431
rect 11529 2397 11563 2431
rect 13277 2397 13311 2431
rect 14381 2397 14415 2431
rect 10977 2329 11011 2363
rect 12633 2329 12667 2363
rect 1593 2261 1627 2295
rect 3525 2261 3559 2295
rect 9321 2261 9355 2295
rect 9781 2261 9815 2295
rect 12173 2261 12207 2295
rect 13829 2261 13863 2295
rect 15025 2261 15059 2295
<< metal1 >>
rect 7558 18436 7564 18488
rect 7616 18476 7622 18488
rect 9398 18476 9404 18488
rect 7616 18448 9404 18476
rect 7616 18436 7622 18448
rect 9398 18436 9404 18448
rect 9456 18436 9462 18488
rect 11422 18096 11428 18148
rect 11480 18136 11486 18148
rect 12066 18136 12072 18148
rect 11480 18108 12072 18136
rect 11480 18096 11486 18108
rect 12066 18096 12072 18108
rect 12124 18096 12130 18148
rect 9674 18028 9680 18080
rect 9732 18068 9738 18080
rect 14458 18068 14464 18080
rect 9732 18040 14464 18068
rect 9732 18028 9738 18040
rect 14458 18028 14464 18040
rect 14516 18068 14522 18080
rect 16022 18068 16028 18080
rect 14516 18040 16028 18068
rect 14516 18028 14522 18040
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 4062 17960 4068 18012
rect 4120 18000 4126 18012
rect 9217 18003 9275 18009
rect 9217 18000 9229 18003
rect 4120 17972 9229 18000
rect 4120 17960 4126 17972
rect 9217 17969 9229 17972
rect 9263 17969 9275 18003
rect 9217 17963 9275 17969
rect 10137 18003 10195 18009
rect 10137 17969 10149 18003
rect 10183 18000 10195 18003
rect 13906 18000 13912 18012
rect 10183 17972 13912 18000
rect 10183 17969 10195 17972
rect 10137 17963 10195 17969
rect 13906 17960 13912 17972
rect 13964 17960 13970 18012
rect 7926 17892 7932 17944
rect 7984 17932 7990 17944
rect 8846 17932 8852 17944
rect 7984 17904 8852 17932
rect 7984 17892 7990 17904
rect 8846 17892 8852 17904
rect 8904 17892 8910 17944
rect 8938 17892 8944 17944
rect 8996 17932 9002 17944
rect 12802 17932 12808 17944
rect 8996 17904 12808 17932
rect 8996 17892 9002 17904
rect 12802 17892 12808 17904
rect 12860 17892 12866 17944
rect 5166 17824 5172 17876
rect 5224 17864 5230 17876
rect 9122 17864 9128 17876
rect 5224 17836 9128 17864
rect 5224 17824 5230 17836
rect 9122 17824 9128 17836
rect 9180 17824 9186 17876
rect 9217 17867 9275 17873
rect 9217 17833 9229 17867
rect 9263 17864 9275 17867
rect 10137 17867 10195 17873
rect 10137 17864 10149 17867
rect 9263 17836 10149 17864
rect 9263 17833 9275 17836
rect 9217 17827 9275 17833
rect 10137 17833 10149 17836
rect 10183 17833 10195 17867
rect 10137 17827 10195 17833
rect 7834 17756 7840 17808
rect 7892 17796 7898 17808
rect 13170 17796 13176 17808
rect 7892 17768 13176 17796
rect 7892 17756 7898 17768
rect 13170 17756 13176 17768
rect 13228 17756 13234 17808
rect 6914 17688 6920 17740
rect 6972 17728 6978 17740
rect 14274 17728 14280 17740
rect 6972 17700 14280 17728
rect 6972 17688 6978 17700
rect 14274 17688 14280 17700
rect 14332 17688 14338 17740
rect 5442 17620 5448 17672
rect 5500 17660 5506 17672
rect 12710 17660 12716 17672
rect 5500 17632 12716 17660
rect 5500 17620 5506 17632
rect 12710 17620 12716 17632
rect 12768 17620 12774 17672
rect 3510 17552 3516 17604
rect 3568 17592 3574 17604
rect 9858 17592 9864 17604
rect 3568 17564 9864 17592
rect 3568 17552 3574 17564
rect 9858 17552 9864 17564
rect 9916 17552 9922 17604
rect 5718 17484 5724 17536
rect 5776 17524 5782 17536
rect 9306 17524 9312 17536
rect 5776 17496 9312 17524
rect 5776 17484 5782 17496
rect 9306 17484 9312 17496
rect 9364 17484 9370 17536
rect 10226 17484 10232 17536
rect 10284 17524 10290 17536
rect 11790 17524 11796 17536
rect 10284 17496 11796 17524
rect 10284 17484 10290 17496
rect 11790 17484 11796 17496
rect 11848 17524 11854 17536
rect 14366 17524 14372 17536
rect 11848 17496 14372 17524
rect 11848 17484 11854 17496
rect 14366 17484 14372 17496
rect 14424 17484 14430 17536
rect 1104 17434 15824 17456
rect 1104 17382 3447 17434
rect 3499 17382 3511 17434
rect 3563 17382 3575 17434
rect 3627 17382 3639 17434
rect 3691 17382 8378 17434
rect 8430 17382 8442 17434
rect 8494 17382 8506 17434
rect 8558 17382 8570 17434
rect 8622 17382 13308 17434
rect 13360 17382 13372 17434
rect 13424 17382 13436 17434
rect 13488 17382 13500 17434
rect 13552 17382 15824 17434
rect 1104 17360 15824 17382
rect 6178 17280 6184 17332
rect 6236 17320 6242 17332
rect 11425 17323 11483 17329
rect 11425 17320 11437 17323
rect 6236 17292 11437 17320
rect 6236 17280 6242 17292
rect 11425 17289 11437 17292
rect 11471 17289 11483 17323
rect 11425 17283 11483 17289
rect 2406 17212 2412 17264
rect 2464 17252 2470 17264
rect 2464 17224 2636 17252
rect 2464 17212 2470 17224
rect 750 17144 756 17196
rect 808 17184 814 17196
rect 1765 17187 1823 17193
rect 808 17156 1624 17184
rect 808 17144 814 17156
rect 1486 17116 1492 17128
rect 1399 17088 1492 17116
rect 1486 17076 1492 17088
rect 1544 17076 1550 17128
rect 1596 17116 1624 17156
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 2130 17184 2136 17196
rect 1811 17156 2136 17184
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 2130 17144 2136 17156
rect 2188 17144 2194 17196
rect 2608 17193 2636 17224
rect 3786 17212 3792 17264
rect 3844 17252 3850 17264
rect 6362 17252 6368 17264
rect 3844 17224 6368 17252
rect 3844 17212 3850 17224
rect 6362 17212 6368 17224
rect 6420 17212 6426 17264
rect 7300 17224 7604 17252
rect 2593 17187 2651 17193
rect 2593 17153 2605 17187
rect 2639 17153 2651 17187
rect 2593 17147 2651 17153
rect 3142 17144 3148 17196
rect 3200 17184 3206 17196
rect 4249 17187 4307 17193
rect 4249 17184 4261 17187
rect 3200 17156 4261 17184
rect 3200 17144 3206 17156
rect 4249 17153 4261 17156
rect 4295 17153 4307 17187
rect 4249 17147 4307 17153
rect 4893 17187 4951 17193
rect 4893 17153 4905 17187
rect 4939 17184 4951 17187
rect 4982 17184 4988 17196
rect 4939 17156 4988 17184
rect 4939 17153 4951 17156
rect 4893 17147 4951 17153
rect 4982 17144 4988 17156
rect 5040 17144 5046 17196
rect 6273 17187 6331 17193
rect 6273 17153 6285 17187
rect 6319 17184 6331 17187
rect 7300 17184 7328 17224
rect 7466 17184 7472 17196
rect 6319 17156 7328 17184
rect 7427 17156 7472 17184
rect 6319 17153 6331 17156
rect 6273 17147 6331 17153
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 7576 17184 7604 17224
rect 7650 17212 7656 17264
rect 7708 17252 7714 17264
rect 8113 17255 8171 17261
rect 8113 17252 8125 17255
rect 7708 17224 8125 17252
rect 7708 17212 7714 17224
rect 8113 17221 8125 17224
rect 8159 17221 8171 17255
rect 8113 17215 8171 17221
rect 8938 17212 8944 17264
rect 8996 17252 9002 17264
rect 9309 17255 9367 17261
rect 9309 17252 9321 17255
rect 8996 17224 9321 17252
rect 8996 17212 9002 17224
rect 9309 17221 9321 17224
rect 9355 17221 9367 17255
rect 9309 17215 9367 17221
rect 9398 17212 9404 17264
rect 9456 17252 9462 17264
rect 12805 17255 12863 17261
rect 12805 17252 12817 17255
rect 9456 17224 12817 17252
rect 9456 17212 9462 17224
rect 12805 17221 12817 17224
rect 12851 17221 12863 17255
rect 12805 17215 12863 17221
rect 8018 17184 8024 17196
rect 7576 17156 8024 17184
rect 8018 17144 8024 17156
rect 8076 17184 8082 17196
rect 8665 17187 8723 17193
rect 8665 17184 8677 17187
rect 8076 17156 8677 17184
rect 8076 17144 8082 17156
rect 8665 17153 8677 17156
rect 8711 17153 8723 17187
rect 8665 17147 8723 17153
rect 2409 17119 2467 17125
rect 2409 17116 2421 17119
rect 1596 17088 2421 17116
rect 2409 17085 2421 17088
rect 2455 17116 2467 17119
rect 2682 17116 2688 17128
rect 2455 17088 2688 17116
rect 2455 17085 2467 17088
rect 2409 17079 2467 17085
rect 2682 17076 2688 17088
rect 2740 17076 2746 17128
rect 3234 17076 3240 17128
rect 3292 17116 3298 17128
rect 4062 17116 4068 17128
rect 3292 17088 4068 17116
rect 3292 17076 3298 17088
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 5534 17076 5540 17128
rect 5592 17116 5598 17128
rect 8846 17116 8852 17128
rect 5592 17088 8852 17116
rect 5592 17076 5598 17088
rect 8846 17076 8852 17088
rect 8904 17076 8910 17128
rect 9490 17076 9496 17128
rect 9548 17116 9554 17128
rect 9769 17119 9827 17125
rect 9548 17088 9593 17116
rect 9548 17076 9554 17088
rect 9769 17085 9781 17119
rect 9815 17116 9827 17119
rect 10042 17116 10048 17128
rect 9815 17088 10048 17116
rect 9815 17085 9827 17088
rect 9769 17079 9827 17085
rect 10042 17076 10048 17088
rect 10100 17076 10106 17128
rect 10410 17076 10416 17128
rect 10468 17116 10474 17128
rect 10505 17119 10563 17125
rect 10505 17116 10517 17119
rect 10468 17088 10517 17116
rect 10468 17076 10474 17088
rect 10505 17085 10517 17088
rect 10551 17085 10563 17119
rect 10505 17079 10563 17085
rect 11241 17119 11299 17125
rect 11241 17085 11253 17119
rect 11287 17116 11299 17119
rect 12526 17116 12532 17128
rect 11287 17088 12532 17116
rect 11287 17085 11299 17088
rect 11241 17079 11299 17085
rect 12526 17076 12532 17088
rect 12584 17076 12590 17128
rect 12621 17119 12679 17125
rect 12621 17085 12633 17119
rect 12667 17116 12679 17119
rect 13078 17116 13084 17128
rect 12667 17088 13084 17116
rect 12667 17085 12679 17088
rect 12621 17079 12679 17085
rect 13078 17076 13084 17088
rect 13136 17076 13142 17128
rect 13357 17119 13415 17125
rect 13357 17085 13369 17119
rect 13403 17085 13415 17119
rect 13357 17079 13415 17085
rect 1504 17048 1532 17076
rect 1854 17048 1860 17060
rect 1504 17020 1860 17048
rect 1854 17008 1860 17020
rect 1912 17008 1918 17060
rect 2958 17008 2964 17060
rect 3016 17048 3022 17060
rect 6270 17048 6276 17060
rect 3016 17020 6276 17048
rect 3016 17008 3022 17020
rect 6270 17008 6276 17020
rect 6328 17008 6334 17060
rect 7377 17051 7435 17057
rect 7377 17017 7389 17051
rect 7423 17048 7435 17051
rect 7926 17048 7932 17060
rect 7423 17020 7932 17048
rect 7423 17017 7435 17020
rect 7377 17011 7435 17017
rect 7926 17008 7932 17020
rect 7984 17008 7990 17060
rect 8478 17048 8484 17060
rect 8439 17020 8484 17048
rect 8478 17008 8484 17020
rect 8536 17008 8542 17060
rect 8573 17051 8631 17057
rect 8573 17017 8585 17051
rect 8619 17048 8631 17051
rect 8754 17048 8760 17060
rect 8619 17020 8760 17048
rect 8619 17017 8631 17020
rect 8573 17011 8631 17017
rect 8754 17008 8760 17020
rect 8812 17008 8818 17060
rect 9582 17008 9588 17060
rect 9640 17048 9646 17060
rect 11422 17048 11428 17060
rect 9640 17020 11428 17048
rect 9640 17008 9646 17020
rect 11422 17008 11428 17020
rect 11480 17008 11486 17060
rect 11698 17008 11704 17060
rect 11756 17048 11762 17060
rect 13372 17048 13400 17079
rect 11756 17020 13400 17048
rect 11756 17008 11762 17020
rect 3237 16983 3295 16989
rect 3237 16949 3249 16983
rect 3283 16980 3295 16983
rect 3326 16980 3332 16992
rect 3283 16952 3332 16980
rect 3283 16949 3295 16952
rect 3237 16943 3295 16949
rect 3326 16940 3332 16952
rect 3384 16940 3390 16992
rect 5626 16980 5632 16992
rect 5587 16952 5632 16980
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 5718 16940 5724 16992
rect 5776 16980 5782 16992
rect 5997 16983 6055 16989
rect 5997 16980 6009 16983
rect 5776 16952 6009 16980
rect 5776 16940 5782 16952
rect 5997 16949 6009 16952
rect 6043 16949 6055 16983
rect 5997 16943 6055 16949
rect 6089 16983 6147 16989
rect 6089 16949 6101 16983
rect 6135 16980 6147 16983
rect 6917 16983 6975 16989
rect 6917 16980 6929 16983
rect 6135 16952 6929 16980
rect 6135 16949 6147 16952
rect 6089 16943 6147 16949
rect 6917 16949 6929 16952
rect 6963 16949 6975 16983
rect 6917 16943 6975 16949
rect 7285 16983 7343 16989
rect 7285 16949 7297 16983
rect 7331 16980 7343 16983
rect 7742 16980 7748 16992
rect 7331 16952 7748 16980
rect 7331 16949 7343 16952
rect 7285 16943 7343 16949
rect 7742 16940 7748 16952
rect 7800 16940 7806 16992
rect 9766 16940 9772 16992
rect 9824 16980 9830 16992
rect 9953 16983 10011 16989
rect 9953 16980 9965 16983
rect 9824 16952 9965 16980
rect 9824 16940 9830 16952
rect 9953 16949 9965 16952
rect 9999 16949 10011 16983
rect 9953 16943 10011 16949
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10689 16983 10747 16989
rect 10689 16980 10701 16983
rect 10192 16952 10701 16980
rect 10192 16940 10198 16952
rect 10689 16949 10701 16952
rect 10735 16949 10747 16983
rect 10689 16943 10747 16949
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 11882 16980 11888 16992
rect 11204 16952 11888 16980
rect 11204 16940 11210 16952
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 13541 16983 13599 16989
rect 13541 16980 13553 16983
rect 12952 16952 13553 16980
rect 12952 16940 12958 16952
rect 13541 16949 13553 16952
rect 13587 16949 13599 16983
rect 13541 16943 13599 16949
rect 1104 16890 15824 16912
rect 1104 16838 5912 16890
rect 5964 16838 5976 16890
rect 6028 16838 6040 16890
rect 6092 16838 6104 16890
rect 6156 16838 10843 16890
rect 10895 16838 10907 16890
rect 10959 16838 10971 16890
rect 11023 16838 11035 16890
rect 11087 16838 15824 16890
rect 1104 16816 15824 16838
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 3697 16779 3755 16785
rect 2832 16748 3096 16776
rect 2832 16736 2838 16748
rect 1670 16708 1676 16720
rect 1631 16680 1676 16708
rect 1670 16668 1676 16680
rect 1728 16668 1734 16720
rect 3068 16717 3096 16748
rect 3697 16745 3709 16779
rect 3743 16776 3755 16779
rect 4614 16776 4620 16788
rect 3743 16748 4620 16776
rect 3743 16745 3755 16748
rect 3697 16739 3755 16745
rect 4614 16736 4620 16748
rect 4672 16736 4678 16788
rect 5442 16776 5448 16788
rect 5403 16748 5448 16776
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 6270 16776 6276 16788
rect 6231 16748 6276 16776
rect 6270 16736 6276 16748
rect 6328 16736 6334 16788
rect 6641 16779 6699 16785
rect 6641 16745 6653 16779
rect 6687 16776 6699 16779
rect 7469 16779 7527 16785
rect 7469 16776 7481 16779
rect 6687 16748 7481 16776
rect 6687 16745 6699 16748
rect 6641 16739 6699 16745
rect 7469 16745 7481 16748
rect 7515 16745 7527 16779
rect 7834 16776 7840 16788
rect 7795 16748 7840 16776
rect 7469 16739 7527 16745
rect 7834 16736 7840 16748
rect 7892 16736 7898 16788
rect 8110 16736 8116 16788
rect 8168 16776 8174 16788
rect 8294 16776 8300 16788
rect 8168 16748 8300 16776
rect 8168 16736 8174 16748
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 8846 16736 8852 16788
rect 8904 16776 8910 16788
rect 8904 16748 11376 16776
rect 8904 16736 8910 16748
rect 3053 16711 3111 16717
rect 3053 16677 3065 16711
rect 3099 16677 3111 16711
rect 3053 16671 3111 16677
rect 3326 16668 3332 16720
rect 3384 16708 3390 16720
rect 3384 16680 4108 16708
rect 3384 16668 3390 16680
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 1578 16640 1584 16652
rect 1443 16612 1584 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 2590 16600 2596 16652
rect 2648 16640 2654 16652
rect 2685 16643 2743 16649
rect 2685 16640 2697 16643
rect 2648 16612 2697 16640
rect 2648 16600 2654 16612
rect 2685 16609 2697 16612
rect 2731 16609 2743 16643
rect 2685 16603 2743 16609
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16609 2835 16643
rect 2777 16603 2835 16609
rect 3881 16643 3939 16649
rect 3881 16609 3893 16643
rect 3927 16640 3939 16643
rect 3970 16640 3976 16652
rect 3927 16612 3976 16640
rect 3927 16609 3939 16612
rect 3881 16603 3939 16609
rect 1118 16532 1124 16584
rect 1176 16572 1182 16584
rect 1486 16572 1492 16584
rect 1176 16544 1492 16572
rect 1176 16532 1182 16544
rect 1486 16532 1492 16544
rect 1544 16572 1550 16584
rect 2792 16572 2820 16603
rect 3970 16600 3976 16612
rect 4028 16600 4034 16652
rect 4080 16649 4108 16680
rect 4522 16668 4528 16720
rect 4580 16708 4586 16720
rect 6733 16711 6791 16717
rect 4580 16680 5488 16708
rect 4580 16668 4586 16680
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 4246 16600 4252 16652
rect 4304 16640 4310 16652
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 4304 16612 4353 16640
rect 4304 16600 4310 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 5350 16640 5356 16652
rect 5311 16612 5356 16640
rect 4341 16603 4399 16609
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 5460 16640 5488 16680
rect 6733 16677 6745 16711
rect 6779 16708 6791 16711
rect 7650 16708 7656 16720
rect 6779 16680 7656 16708
rect 6779 16677 6791 16680
rect 6733 16671 6791 16677
rect 7650 16668 7656 16680
rect 7708 16668 7714 16720
rect 9030 16708 9036 16720
rect 8680 16680 9036 16708
rect 8680 16649 8708 16680
rect 9030 16668 9036 16680
rect 9088 16668 9094 16720
rect 9306 16668 9312 16720
rect 9364 16708 9370 16720
rect 9364 16680 10456 16708
rect 9364 16668 9370 16680
rect 8665 16643 8723 16649
rect 5460 16612 8616 16640
rect 1544 16544 2820 16572
rect 5537 16575 5595 16581
rect 1544 16532 1550 16544
rect 5537 16541 5549 16575
rect 5583 16541 5595 16575
rect 5537 16535 5595 16541
rect 1578 16464 1584 16516
rect 1636 16504 1642 16516
rect 3234 16504 3240 16516
rect 1636 16476 3240 16504
rect 1636 16464 1642 16476
rect 3234 16464 3240 16476
rect 3292 16464 3298 16516
rect 3878 16464 3884 16516
rect 3936 16504 3942 16516
rect 4985 16507 5043 16513
rect 4985 16504 4997 16507
rect 3936 16476 4997 16504
rect 3936 16464 3942 16476
rect 4985 16473 4997 16476
rect 5031 16473 5043 16507
rect 4985 16467 5043 16473
rect 5074 16464 5080 16516
rect 5132 16504 5138 16516
rect 5552 16504 5580 16535
rect 6638 16532 6644 16584
rect 6696 16572 6702 16584
rect 6825 16575 6883 16581
rect 6825 16572 6837 16575
rect 6696 16544 6837 16572
rect 6696 16532 6702 16544
rect 6825 16541 6837 16544
rect 6871 16541 6883 16575
rect 6825 16535 6883 16541
rect 7190 16532 7196 16584
rect 7248 16572 7254 16584
rect 7650 16572 7656 16584
rect 7248 16544 7656 16572
rect 7248 16532 7254 16544
rect 7650 16532 7656 16544
rect 7708 16532 7714 16584
rect 7742 16532 7748 16584
rect 7800 16572 7806 16584
rect 7929 16575 7987 16581
rect 7929 16572 7941 16575
rect 7800 16544 7941 16572
rect 7800 16532 7806 16544
rect 7929 16541 7941 16544
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 8021 16575 8079 16581
rect 8021 16541 8033 16575
rect 8067 16541 8079 16575
rect 8588 16572 8616 16612
rect 8665 16609 8677 16643
rect 8711 16609 8723 16643
rect 8665 16603 8723 16609
rect 8846 16600 8852 16652
rect 8904 16640 8910 16652
rect 8941 16643 8999 16649
rect 8941 16640 8953 16643
rect 8904 16612 8953 16640
rect 8904 16600 8910 16612
rect 8941 16609 8953 16612
rect 8987 16609 8999 16643
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 8941 16603 8999 16609
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 10428 16649 10456 16680
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16609 10471 16643
rect 10413 16603 10471 16609
rect 11149 16643 11207 16649
rect 11149 16609 11161 16643
rect 11195 16609 11207 16643
rect 11149 16603 11207 16609
rect 8588 16544 10088 16572
rect 8021 16535 8079 16541
rect 5132 16476 5580 16504
rect 5132 16464 5138 16476
rect 8036 16448 8064 16535
rect 8202 16464 8208 16516
rect 8260 16504 8266 16516
rect 9766 16504 9772 16516
rect 8260 16476 9772 16504
rect 8260 16464 8266 16476
rect 9766 16464 9772 16476
rect 9824 16464 9830 16516
rect 9858 16464 9864 16516
rect 9916 16504 9922 16516
rect 10060 16504 10088 16544
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 11164 16572 11192 16603
rect 10192 16544 11192 16572
rect 10192 16532 10198 16544
rect 11348 16513 11376 16748
rect 11422 16736 11428 16788
rect 11480 16776 11486 16788
rect 12069 16779 12127 16785
rect 12069 16776 12081 16779
rect 11480 16748 12081 16776
rect 11480 16736 11486 16748
rect 12069 16745 12081 16748
rect 12115 16745 12127 16779
rect 12069 16739 12127 16745
rect 12250 16736 12256 16788
rect 12308 16776 12314 16788
rect 13541 16779 13599 16785
rect 13541 16776 13553 16779
rect 12308 16748 13553 16776
rect 12308 16736 12314 16748
rect 13541 16745 13553 16748
rect 13587 16745 13599 16779
rect 14274 16776 14280 16788
rect 14235 16748 14280 16776
rect 13541 16739 13599 16745
rect 14274 16736 14280 16748
rect 14332 16736 14338 16788
rect 11532 16680 12112 16708
rect 11532 16652 11560 16680
rect 12084 16652 12112 16680
rect 12158 16668 12164 16720
rect 12216 16708 12222 16720
rect 12216 16680 13400 16708
rect 12216 16668 12222 16680
rect 11514 16600 11520 16652
rect 11572 16600 11578 16652
rect 11882 16640 11888 16652
rect 11843 16612 11888 16640
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 12066 16600 12072 16652
rect 12124 16600 12130 16652
rect 12434 16600 12440 16652
rect 12492 16640 12498 16652
rect 13372 16649 13400 16680
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 12492 16612 12633 16640
rect 12492 16600 12498 16612
rect 12621 16609 12633 16612
rect 12667 16609 12679 16643
rect 12621 16603 12679 16609
rect 13357 16643 13415 16649
rect 13357 16609 13369 16643
rect 13403 16609 13415 16643
rect 14090 16640 14096 16652
rect 14051 16612 14096 16640
rect 13357 16603 13415 16609
rect 14090 16600 14096 16612
rect 14148 16600 14154 16652
rect 10597 16507 10655 16513
rect 10597 16504 10609 16507
rect 9916 16476 9961 16504
rect 10060 16476 10609 16504
rect 9916 16464 9922 16476
rect 10597 16473 10609 16476
rect 10643 16473 10655 16507
rect 10597 16467 10655 16473
rect 11333 16507 11391 16513
rect 11333 16473 11345 16507
rect 11379 16473 11391 16507
rect 12802 16504 12808 16516
rect 12763 16476 12808 16504
rect 11333 16467 11391 16473
rect 12802 16464 12808 16476
rect 12860 16464 12866 16516
rect 2501 16439 2559 16445
rect 2501 16405 2513 16439
rect 2547 16436 2559 16439
rect 3786 16436 3792 16448
rect 2547 16408 3792 16436
rect 2547 16405 2559 16408
rect 2501 16399 2559 16405
rect 3786 16396 3792 16408
rect 3844 16396 3850 16448
rect 6362 16396 6368 16448
rect 6420 16436 6426 16448
rect 7834 16436 7840 16448
rect 6420 16408 7840 16436
rect 6420 16396 6426 16408
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 8018 16396 8024 16448
rect 8076 16396 8082 16448
rect 8662 16396 8668 16448
rect 8720 16436 8726 16448
rect 11422 16436 11428 16448
rect 8720 16408 11428 16436
rect 8720 16396 8726 16408
rect 11422 16396 11428 16408
rect 11480 16396 11486 16448
rect 1104 16346 15824 16368
rect 1104 16294 3447 16346
rect 3499 16294 3511 16346
rect 3563 16294 3575 16346
rect 3627 16294 3639 16346
rect 3691 16294 8378 16346
rect 8430 16294 8442 16346
rect 8494 16294 8506 16346
rect 8558 16294 8570 16346
rect 8622 16294 13308 16346
rect 13360 16294 13372 16346
rect 13424 16294 13436 16346
rect 13488 16294 13500 16346
rect 13552 16294 15824 16346
rect 1104 16272 15824 16294
rect 1854 16192 1860 16244
rect 1912 16232 1918 16244
rect 4062 16232 4068 16244
rect 1912 16204 4068 16232
rect 1912 16192 1918 16204
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 4341 16235 4399 16241
rect 4341 16201 4353 16235
rect 4387 16232 4399 16235
rect 4706 16232 4712 16244
rect 4387 16204 4712 16232
rect 4387 16201 4399 16204
rect 4341 16195 4399 16201
rect 4706 16192 4712 16204
rect 4764 16192 4770 16244
rect 4798 16192 4804 16244
rect 4856 16232 4862 16244
rect 9858 16232 9864 16244
rect 4856 16204 9864 16232
rect 4856 16192 4862 16204
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 9950 16192 9956 16244
rect 10008 16232 10014 16244
rect 10597 16235 10655 16241
rect 10597 16232 10609 16235
rect 10008 16204 10609 16232
rect 10008 16192 10014 16204
rect 10597 16201 10609 16204
rect 10643 16201 10655 16235
rect 10597 16195 10655 16201
rect 11238 16192 11244 16244
rect 11296 16232 11302 16244
rect 12342 16232 12348 16244
rect 11296 16204 12348 16232
rect 11296 16192 11302 16204
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 5810 16124 5816 16176
rect 5868 16164 5874 16176
rect 6638 16164 6644 16176
rect 5868 16136 6644 16164
rect 5868 16124 5874 16136
rect 1394 16056 1400 16108
rect 1452 16096 1458 16108
rect 1673 16099 1731 16105
rect 1673 16096 1685 16099
rect 1452 16068 1685 16096
rect 1452 16056 1458 16068
rect 1673 16065 1685 16068
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 1762 16056 1768 16108
rect 1820 16096 1826 16108
rect 2593 16099 2651 16105
rect 2593 16096 2605 16099
rect 1820 16068 2605 16096
rect 1820 16056 1826 16068
rect 2593 16065 2605 16068
rect 2639 16065 2651 16099
rect 2593 16059 2651 16065
rect 4985 16099 5043 16105
rect 4985 16065 4997 16099
rect 5031 16096 5043 16099
rect 5534 16096 5540 16108
rect 5031 16068 5540 16096
rect 5031 16065 5043 16068
rect 4985 16059 5043 16065
rect 5534 16056 5540 16068
rect 5592 16056 5598 16108
rect 5626 16056 5632 16108
rect 5684 16096 5690 16108
rect 6104 16105 6132 16136
rect 6638 16124 6644 16136
rect 6696 16124 6702 16176
rect 6822 16164 6828 16176
rect 6783 16136 6828 16164
rect 6822 16124 6828 16136
rect 6880 16124 6886 16176
rect 6914 16124 6920 16176
rect 6972 16164 6978 16176
rect 6972 16136 9812 16164
rect 6972 16124 6978 16136
rect 5997 16099 6055 16105
rect 5997 16096 6009 16099
rect 5684 16068 6009 16096
rect 5684 16056 5690 16068
rect 5997 16065 6009 16068
rect 6043 16065 6055 16099
rect 5997 16059 6055 16065
rect 6089 16099 6147 16105
rect 6089 16065 6101 16099
rect 6135 16065 6147 16099
rect 7374 16096 7380 16108
rect 7335 16068 7380 16096
rect 6089 16059 6147 16065
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 7558 16056 7564 16108
rect 7616 16056 7622 16108
rect 7926 16056 7932 16108
rect 7984 16096 7990 16108
rect 8478 16096 8484 16108
rect 7984 16068 8484 16096
rect 7984 16056 7990 16068
rect 8478 16056 8484 16068
rect 8536 16056 8542 16108
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16065 8631 16099
rect 8573 16059 8631 16065
rect 106 15988 112 16040
rect 164 16028 170 16040
rect 1302 16028 1308 16040
rect 164 16000 1308 16028
rect 164 15988 170 16000
rect 1302 15988 1308 16000
rect 1360 16028 1366 16040
rect 2406 16037 2412 16040
rect 1489 16031 1547 16037
rect 1489 16028 1501 16031
rect 1360 16000 1501 16028
rect 1360 15988 1366 16000
rect 1489 15997 1501 16000
rect 1535 15997 1547 16031
rect 2398 16031 2412 16037
rect 2398 16028 2410 16031
rect 1489 15991 1547 15997
rect 1596 16000 2410 16028
rect 382 15920 388 15972
rect 440 15960 446 15972
rect 1596 15960 1624 16000
rect 2398 15997 2410 16000
rect 2398 15991 2412 15997
rect 2406 15988 2412 15991
rect 2464 15988 2470 16040
rect 3329 16031 3387 16037
rect 3329 15997 3341 16031
rect 3375 16028 3387 16031
rect 4430 16028 4436 16040
rect 3375 16000 4436 16028
rect 3375 15997 3387 16000
rect 3329 15991 3387 15997
rect 4430 15988 4436 16000
rect 4488 15988 4494 16040
rect 7190 16028 7196 16040
rect 7151 16000 7196 16028
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 7285 16031 7343 16037
rect 7285 15997 7297 16031
rect 7331 16028 7343 16031
rect 7576 16028 7604 16056
rect 7331 16000 7604 16028
rect 7331 15997 7343 16000
rect 7285 15991 7343 15997
rect 7742 15988 7748 16040
rect 7800 16028 7806 16040
rect 8294 16028 8300 16040
rect 7800 16000 8300 16028
rect 7800 15988 7806 16000
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 3602 15960 3608 15972
rect 440 15932 1624 15960
rect 3563 15932 3608 15960
rect 440 15920 446 15932
rect 3602 15920 3608 15932
rect 3660 15920 3666 15972
rect 4706 15960 4712 15972
rect 4667 15932 4712 15960
rect 4706 15920 4712 15932
rect 4764 15920 4770 15972
rect 5905 15963 5963 15969
rect 5905 15929 5917 15963
rect 5951 15960 5963 15963
rect 6178 15960 6184 15972
rect 5951 15932 6184 15960
rect 5951 15929 5963 15932
rect 5905 15923 5963 15929
rect 6178 15920 6184 15932
rect 6236 15920 6242 15972
rect 7558 15920 7564 15972
rect 7616 15960 7622 15972
rect 8588 15960 8616 16059
rect 9122 16056 9128 16108
rect 9180 16096 9186 16108
rect 9784 16105 9812 16136
rect 10778 16124 10784 16176
rect 10836 16164 10842 16176
rect 12894 16164 12900 16176
rect 10836 16136 12900 16164
rect 10836 16124 10842 16136
rect 12894 16124 12900 16136
rect 12952 16124 12958 16176
rect 13357 16167 13415 16173
rect 13357 16133 13369 16167
rect 13403 16133 13415 16167
rect 13357 16127 13415 16133
rect 9769 16099 9827 16105
rect 9180 16068 9352 16096
rect 9180 16056 9186 16068
rect 9122 15960 9128 15972
rect 7616 15932 8616 15960
rect 8680 15932 9128 15960
rect 7616 15920 7622 15932
rect 4798 15892 4804 15904
rect 4759 15864 4804 15892
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 5537 15895 5595 15901
rect 5537 15892 5549 15895
rect 5224 15864 5549 15892
rect 5224 15852 5230 15864
rect 5537 15861 5549 15864
rect 5583 15861 5595 15895
rect 5537 15855 5595 15861
rect 7374 15852 7380 15904
rect 7432 15892 7438 15904
rect 8021 15895 8079 15901
rect 8021 15892 8033 15895
rect 7432 15864 8033 15892
rect 7432 15852 7438 15864
rect 8021 15861 8033 15864
rect 8067 15861 8079 15895
rect 8386 15892 8392 15904
rect 8347 15864 8392 15892
rect 8021 15855 8079 15861
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 8481 15895 8539 15901
rect 8481 15861 8493 15895
rect 8527 15892 8539 15895
rect 8680 15892 8708 15932
rect 9122 15920 9128 15932
rect 9180 15920 9186 15972
rect 9324 15960 9352 16068
rect 9769 16065 9781 16099
rect 9815 16065 9827 16099
rect 9769 16059 9827 16065
rect 10686 16056 10692 16108
rect 10744 16096 10750 16108
rect 13372 16096 13400 16127
rect 10744 16068 13400 16096
rect 10744 16056 10750 16068
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 16028 9735 16031
rect 10226 16028 10232 16040
rect 9723 16000 10232 16028
rect 9723 15997 9735 16000
rect 9677 15991 9735 15997
rect 10226 15988 10232 16000
rect 10284 15988 10290 16040
rect 10413 16031 10471 16037
rect 10413 15997 10425 16031
rect 10459 15997 10471 16031
rect 10413 15991 10471 15997
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 16028 11207 16031
rect 11330 16028 11336 16040
rect 11195 16000 11336 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 10428 15960 10456 15991
rect 11330 15988 11336 16000
rect 11388 15988 11394 16040
rect 12342 15988 12348 16040
rect 12400 16028 12406 16040
rect 12437 16031 12495 16037
rect 12437 16028 12449 16031
rect 12400 16000 12449 16028
rect 12400 15988 12406 16000
rect 12437 15997 12449 16000
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 13173 16031 13231 16037
rect 13173 15997 13185 16031
rect 13219 15997 13231 16031
rect 13173 15991 13231 15997
rect 11882 15960 11888 15972
rect 9324 15932 9720 15960
rect 10428 15932 11888 15960
rect 8527 15864 8708 15892
rect 8527 15861 8539 15864
rect 8481 15855 8539 15861
rect 8754 15852 8760 15904
rect 8812 15892 8818 15904
rect 9217 15895 9275 15901
rect 9217 15892 9229 15895
rect 8812 15864 9229 15892
rect 8812 15852 8818 15864
rect 9217 15861 9229 15864
rect 9263 15861 9275 15895
rect 9217 15855 9275 15861
rect 9490 15852 9496 15904
rect 9548 15892 9554 15904
rect 9585 15895 9643 15901
rect 9585 15892 9597 15895
rect 9548 15864 9597 15892
rect 9548 15852 9554 15864
rect 9585 15861 9597 15864
rect 9631 15861 9643 15895
rect 9692 15892 9720 15932
rect 11882 15920 11888 15932
rect 11940 15920 11946 15972
rect 12066 15920 12072 15972
rect 12124 15960 12130 15972
rect 13188 15960 13216 15991
rect 12124 15932 13216 15960
rect 12124 15920 12130 15932
rect 11333 15895 11391 15901
rect 11333 15892 11345 15895
rect 9692 15864 11345 15892
rect 9585 15855 9643 15861
rect 11333 15861 11345 15864
rect 11379 15861 11391 15895
rect 11333 15855 11391 15861
rect 11422 15852 11428 15904
rect 11480 15892 11486 15904
rect 12621 15895 12679 15901
rect 12621 15892 12633 15895
rect 11480 15864 12633 15892
rect 11480 15852 11486 15864
rect 12621 15861 12633 15864
rect 12667 15861 12679 15895
rect 12621 15855 12679 15861
rect 1104 15802 15824 15824
rect 1104 15750 5912 15802
rect 5964 15750 5976 15802
rect 6028 15750 6040 15802
rect 6092 15750 6104 15802
rect 6156 15750 10843 15802
rect 10895 15750 10907 15802
rect 10959 15750 10971 15802
rect 11023 15750 11035 15802
rect 11087 15750 15824 15802
rect 1104 15728 15824 15750
rect 3050 15648 3056 15700
rect 3108 15688 3114 15700
rect 3421 15691 3479 15697
rect 3421 15688 3433 15691
rect 3108 15660 3433 15688
rect 3108 15648 3114 15660
rect 3421 15657 3433 15660
rect 3467 15657 3479 15691
rect 3421 15651 3479 15657
rect 4522 15648 4528 15700
rect 4580 15688 4586 15700
rect 7193 15691 7251 15697
rect 7193 15688 7205 15691
rect 4580 15660 7205 15688
rect 4580 15648 4586 15660
rect 7193 15657 7205 15660
rect 7239 15688 7251 15691
rect 7282 15688 7288 15700
rect 7239 15660 7288 15688
rect 7239 15657 7251 15660
rect 7193 15651 7251 15657
rect 7282 15648 7288 15660
rect 7340 15648 7346 15700
rect 8110 15688 8116 15700
rect 8071 15660 8116 15688
rect 8110 15648 8116 15660
rect 8168 15648 8174 15700
rect 10045 15691 10103 15697
rect 10045 15657 10057 15691
rect 10091 15688 10103 15691
rect 10091 15660 10272 15688
rect 10091 15657 10103 15660
rect 10045 15651 10103 15657
rect 4985 15623 5043 15629
rect 4985 15589 4997 15623
rect 5031 15620 5043 15623
rect 6822 15620 6828 15632
rect 5031 15592 6828 15620
rect 5031 15589 5043 15592
rect 4985 15583 5043 15589
rect 6822 15580 6828 15592
rect 6880 15580 6886 15632
rect 8202 15580 8208 15632
rect 8260 15620 8266 15632
rect 9766 15620 9772 15632
rect 8260 15592 9772 15620
rect 8260 15580 8266 15592
rect 9766 15580 9772 15592
rect 9824 15580 9830 15632
rect 10244 15620 10272 15660
rect 12250 15648 12256 15700
rect 12308 15688 12314 15700
rect 12529 15691 12587 15697
rect 12529 15688 12541 15691
rect 12308 15660 12541 15688
rect 12308 15648 12314 15660
rect 12529 15657 12541 15660
rect 12575 15657 12587 15691
rect 12529 15651 12587 15657
rect 11238 15620 11244 15632
rect 10244 15592 11244 15620
rect 11238 15580 11244 15592
rect 11296 15580 11302 15632
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15521 1455 15555
rect 1397 15515 1455 15521
rect 1412 15348 1440 15515
rect 1486 15512 1492 15564
rect 1544 15552 1550 15564
rect 2317 15555 2375 15561
rect 2317 15552 2329 15555
rect 1544 15524 2329 15552
rect 1544 15512 1550 15524
rect 2317 15521 2329 15524
rect 2363 15521 2375 15555
rect 3234 15552 3240 15564
rect 3195 15524 3240 15552
rect 2317 15515 2375 15521
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 6080 15555 6138 15561
rect 6080 15521 6092 15555
rect 6126 15552 6138 15555
rect 8018 15552 8024 15564
rect 6126 15524 7880 15552
rect 7979 15524 8024 15552
rect 6126 15521 6138 15524
rect 6080 15515 6138 15521
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 1688 15416 1716 15447
rect 2038 15444 2044 15496
rect 2096 15484 2102 15496
rect 2501 15487 2559 15493
rect 2501 15484 2513 15487
rect 2096 15456 2513 15484
rect 2096 15444 2102 15456
rect 2501 15453 2513 15456
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 4338 15444 4344 15496
rect 4396 15484 4402 15496
rect 5077 15487 5135 15493
rect 5077 15484 5089 15487
rect 4396 15456 5089 15484
rect 4396 15444 4402 15456
rect 5077 15453 5089 15456
rect 5123 15453 5135 15487
rect 5077 15447 5135 15453
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15484 5319 15487
rect 5718 15484 5724 15496
rect 5307 15456 5724 15484
rect 5307 15453 5319 15456
rect 5261 15447 5319 15453
rect 5718 15444 5724 15456
rect 5776 15444 5782 15496
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15453 5871 15487
rect 7852 15484 7880 15524
rect 8018 15512 8024 15524
rect 8076 15512 8082 15564
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 8849 15555 8907 15561
rect 8849 15552 8861 15555
rect 8536 15524 8861 15552
rect 8536 15512 8542 15524
rect 8849 15521 8861 15524
rect 8895 15552 8907 15555
rect 9306 15552 9312 15564
rect 8895 15524 9312 15552
rect 8895 15521 8907 15524
rect 8849 15515 8907 15521
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 10226 15512 10232 15564
rect 10284 15552 10290 15564
rect 10594 15552 10600 15564
rect 10284 15524 10600 15552
rect 10284 15512 10290 15524
rect 10594 15512 10600 15524
rect 10652 15552 10658 15564
rect 10873 15555 10931 15561
rect 10873 15552 10885 15555
rect 10652 15524 10885 15552
rect 10652 15512 10658 15524
rect 10873 15521 10885 15524
rect 10919 15521 10931 15555
rect 10873 15515 10931 15521
rect 11422 15512 11428 15564
rect 11480 15552 11486 15564
rect 11609 15555 11667 15561
rect 11609 15552 11621 15555
rect 11480 15524 11621 15552
rect 11480 15512 11486 15524
rect 11609 15521 11621 15524
rect 11655 15521 11667 15555
rect 11609 15515 11667 15521
rect 11790 15512 11796 15564
rect 11848 15552 11854 15564
rect 12250 15552 12256 15564
rect 11848 15524 12256 15552
rect 11848 15512 11854 15524
rect 12250 15512 12256 15524
rect 12308 15512 12314 15564
rect 12345 15555 12403 15561
rect 12345 15521 12357 15555
rect 12391 15521 12403 15555
rect 12345 15515 12403 15521
rect 8110 15484 8116 15496
rect 7852 15456 8116 15484
rect 5813 15447 5871 15453
rect 2682 15416 2688 15428
rect 1688 15388 2688 15416
rect 2682 15376 2688 15388
rect 2740 15376 2746 15428
rect 4982 15376 4988 15428
rect 5040 15416 5046 15428
rect 5626 15416 5632 15428
rect 5040 15388 5632 15416
rect 5040 15376 5046 15388
rect 5626 15376 5632 15388
rect 5684 15416 5690 15428
rect 5828 15416 5856 15447
rect 8110 15444 8116 15456
rect 8168 15484 8174 15496
rect 8205 15487 8263 15493
rect 8205 15484 8217 15487
rect 8168 15456 8217 15484
rect 8168 15444 8174 15456
rect 8205 15453 8217 15456
rect 8251 15453 8263 15487
rect 8205 15447 8263 15453
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 8662 15484 8668 15496
rect 8352 15456 8668 15484
rect 8352 15444 8358 15456
rect 8662 15444 8668 15456
rect 8720 15444 8726 15496
rect 10134 15484 10140 15496
rect 10095 15456 10140 15484
rect 10134 15444 10140 15456
rect 10192 15444 10198 15496
rect 10321 15487 10379 15493
rect 10321 15453 10333 15487
rect 10367 15484 10379 15487
rect 10686 15484 10692 15496
rect 10367 15456 10692 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 10686 15444 10692 15456
rect 10744 15444 10750 15496
rect 11698 15444 11704 15496
rect 11756 15484 11762 15496
rect 12360 15484 12388 15515
rect 11756 15456 12388 15484
rect 11756 15444 11762 15456
rect 12894 15444 12900 15496
rect 12952 15484 12958 15496
rect 13081 15487 13139 15493
rect 13081 15484 13093 15487
rect 12952 15456 13093 15484
rect 12952 15444 12958 15456
rect 13081 15453 13093 15456
rect 13127 15453 13139 15487
rect 13081 15447 13139 15453
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 13998 15484 14004 15496
rect 13771 15456 14004 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 13998 15444 14004 15456
rect 14056 15444 14062 15496
rect 8386 15416 8392 15428
rect 5684 15388 5856 15416
rect 6748 15388 8392 15416
rect 5684 15376 5690 15388
rect 2314 15348 2320 15360
rect 1412 15320 2320 15348
rect 2314 15308 2320 15320
rect 2372 15308 2378 15360
rect 4154 15308 4160 15360
rect 4212 15348 4218 15360
rect 4617 15351 4675 15357
rect 4617 15348 4629 15351
rect 4212 15320 4629 15348
rect 4212 15308 4218 15320
rect 4617 15317 4629 15320
rect 4663 15317 4675 15351
rect 4617 15311 4675 15317
rect 5350 15308 5356 15360
rect 5408 15348 5414 15360
rect 6748 15348 6776 15388
rect 8386 15376 8392 15388
rect 8444 15376 8450 15428
rect 9214 15376 9220 15428
rect 9272 15416 9278 15428
rect 11057 15419 11115 15425
rect 11057 15416 11069 15419
rect 9272 15388 11069 15416
rect 9272 15376 9278 15388
rect 11057 15385 11069 15388
rect 11103 15385 11115 15419
rect 11790 15416 11796 15428
rect 11751 15388 11796 15416
rect 11057 15379 11115 15385
rect 11790 15376 11796 15388
rect 11848 15376 11854 15428
rect 5408 15320 6776 15348
rect 5408 15308 5414 15320
rect 6914 15308 6920 15360
rect 6972 15348 6978 15360
rect 7190 15348 7196 15360
rect 6972 15320 7196 15348
rect 6972 15308 6978 15320
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 7650 15348 7656 15360
rect 7611 15320 7656 15348
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 7834 15308 7840 15360
rect 7892 15348 7898 15360
rect 9033 15351 9091 15357
rect 9033 15348 9045 15351
rect 7892 15320 9045 15348
rect 7892 15308 7898 15320
rect 9033 15317 9045 15320
rect 9079 15317 9091 15351
rect 9033 15311 9091 15317
rect 9677 15351 9735 15357
rect 9677 15317 9689 15351
rect 9723 15348 9735 15351
rect 9766 15348 9772 15360
rect 9723 15320 9772 15348
rect 9723 15317 9735 15320
rect 9677 15311 9735 15317
rect 9766 15308 9772 15320
rect 9824 15308 9830 15360
rect 1104 15258 15824 15280
rect 1104 15206 3447 15258
rect 3499 15206 3511 15258
rect 3563 15206 3575 15258
rect 3627 15206 3639 15258
rect 3691 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 13308 15258
rect 13360 15206 13372 15258
rect 13424 15206 13436 15258
rect 13488 15206 13500 15258
rect 13552 15206 15824 15258
rect 1104 15184 15824 15206
rect 3697 15147 3755 15153
rect 3697 15113 3709 15147
rect 3743 15144 3755 15147
rect 4798 15144 4804 15156
rect 3743 15116 4804 15144
rect 3743 15113 3755 15116
rect 3697 15107 3755 15113
rect 4798 15104 4804 15116
rect 4856 15104 4862 15156
rect 5258 15144 5264 15156
rect 4908 15116 5264 15144
rect 3418 15036 3424 15088
rect 3476 15076 3482 15088
rect 4908 15076 4936 15116
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 5920 15116 8217 15144
rect 3476 15048 4936 15076
rect 3476 15036 3482 15048
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 15008 2099 15011
rect 3050 15008 3056 15020
rect 2087 14980 3056 15008
rect 2087 14977 2099 14980
rect 2041 14971 2099 14977
rect 3050 14968 3056 14980
rect 3108 14968 3114 15020
rect 4154 15008 4160 15020
rect 4115 14980 4160 15008
rect 4154 14968 4160 14980
rect 4212 14968 4218 15020
rect 4356 15017 4384 15048
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 14977 4399 15011
rect 4341 14971 4399 14977
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 1854 14900 1860 14952
rect 1912 14940 1918 14952
rect 2685 14943 2743 14949
rect 2685 14940 2697 14943
rect 1912 14912 2697 14940
rect 1912 14900 1918 14912
rect 2685 14909 2697 14912
rect 2731 14909 2743 14943
rect 2685 14903 2743 14909
rect 3786 14900 3792 14952
rect 3844 14940 3850 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 3844 14912 4905 14940
rect 3844 14900 3850 14912
rect 4893 14909 4905 14912
rect 4939 14940 4951 14943
rect 4982 14940 4988 14952
rect 4939 14912 4988 14940
rect 4939 14909 4951 14912
rect 4893 14903 4951 14909
rect 4982 14900 4988 14912
rect 5040 14900 5046 14952
rect 5160 14943 5218 14949
rect 5160 14909 5172 14943
rect 5206 14940 5218 14943
rect 5920 14940 5948 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 8662 15144 8668 15156
rect 8623 15116 8668 15144
rect 8205 15107 8263 15113
rect 8662 15104 8668 15116
rect 8720 15104 8726 15156
rect 9122 15104 9128 15156
rect 9180 15144 9186 15156
rect 9861 15147 9919 15153
rect 9861 15144 9873 15147
rect 9180 15116 9873 15144
rect 9180 15104 9186 15116
rect 9861 15113 9873 15116
rect 9907 15113 9919 15147
rect 9861 15107 9919 15113
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10870 15144 10876 15156
rect 10008 15116 10876 15144
rect 10008 15104 10014 15116
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 10980 15116 12388 15144
rect 8018 15036 8024 15088
rect 8076 15076 8082 15088
rect 10980 15076 11008 15116
rect 8076 15048 11008 15076
rect 8076 15036 8082 15048
rect 11054 15036 11060 15088
rect 11112 15076 11118 15088
rect 11112 15048 11157 15076
rect 11112 15036 11118 15048
rect 6546 14968 6552 15020
rect 6604 15008 6610 15020
rect 6604 14980 6960 15008
rect 6604 14968 6610 14980
rect 5206 14912 5948 14940
rect 5206 14909 5218 14912
rect 5160 14903 5218 14909
rect 2961 14875 3019 14881
rect 2961 14841 2973 14875
rect 3007 14872 3019 14875
rect 3234 14872 3240 14884
rect 3007 14844 3240 14872
rect 3007 14841 3019 14844
rect 2961 14835 3019 14841
rect 3234 14832 3240 14844
rect 3292 14832 3298 14884
rect 4154 14832 4160 14884
rect 4212 14872 4218 14884
rect 5175 14872 5203 14903
rect 6730 14900 6736 14952
rect 6788 14940 6794 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6788 14912 6837 14940
rect 6788 14900 6794 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6932 14940 6960 14980
rect 8110 14968 8116 15020
rect 8168 15008 8174 15020
rect 9214 15008 9220 15020
rect 8168 14980 9220 15008
rect 8168 14968 8174 14980
rect 9214 14968 9220 14980
rect 9272 14968 9278 15020
rect 9490 14968 9496 15020
rect 9548 15008 9554 15020
rect 10413 15011 10471 15017
rect 10413 15008 10425 15011
rect 9548 14980 10425 15008
rect 9548 14968 9554 14980
rect 10413 14977 10425 14980
rect 10459 14977 10471 15011
rect 11514 15008 11520 15020
rect 11475 14980 11520 15008
rect 10413 14971 10471 14977
rect 11514 14968 11520 14980
rect 11572 14968 11578 15020
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 15008 11759 15011
rect 11790 15008 11796 15020
rect 11747 14980 11796 15008
rect 11747 14977 11759 14980
rect 11701 14971 11759 14977
rect 11790 14968 11796 14980
rect 11848 14968 11854 15020
rect 12360 15008 12388 15116
rect 13725 15011 13783 15017
rect 13725 15008 13737 15011
rect 12360 14980 13737 15008
rect 13725 14977 13737 14980
rect 13771 14977 13783 15011
rect 13725 14971 13783 14977
rect 7092 14943 7150 14949
rect 7092 14940 7104 14943
rect 6932 14912 7104 14940
rect 6825 14903 6883 14909
rect 7092 14909 7104 14912
rect 7138 14940 7150 14943
rect 7558 14940 7564 14952
rect 7138 14912 7564 14940
rect 7138 14909 7150 14912
rect 7092 14903 7150 14909
rect 7558 14900 7564 14912
rect 7616 14900 7622 14952
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14940 9091 14943
rect 12434 14940 12440 14952
rect 9079 14912 12440 14940
rect 9079 14909 9091 14912
rect 9033 14903 9091 14909
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 8294 14872 8300 14884
rect 4212 14844 5203 14872
rect 5368 14844 8300 14872
rect 4212 14832 4218 14844
rect 4065 14807 4123 14813
rect 4065 14773 4077 14807
rect 4111 14804 4123 14807
rect 5368 14804 5396 14844
rect 8294 14832 8300 14844
rect 8352 14832 8358 14884
rect 8386 14832 8392 14884
rect 8444 14872 8450 14884
rect 9950 14872 9956 14884
rect 8444 14844 9956 14872
rect 8444 14832 8450 14844
rect 9950 14832 9956 14844
rect 10008 14832 10014 14884
rect 10229 14875 10287 14881
rect 10229 14841 10241 14875
rect 10275 14872 10287 14875
rect 10502 14872 10508 14884
rect 10275 14844 10508 14872
rect 10275 14841 10287 14844
rect 10229 14835 10287 14841
rect 10502 14832 10508 14844
rect 10560 14832 10566 14884
rect 13081 14875 13139 14881
rect 13081 14872 13093 14875
rect 11072 14844 13093 14872
rect 4111 14776 5396 14804
rect 4111 14773 4123 14776
rect 4065 14767 4123 14773
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 6273 14807 6331 14813
rect 6273 14804 6285 14807
rect 5500 14776 6285 14804
rect 5500 14764 5506 14776
rect 6273 14773 6285 14776
rect 6319 14804 6331 14807
rect 8110 14804 8116 14816
rect 6319 14776 8116 14804
rect 6319 14773 6331 14776
rect 6273 14767 6331 14773
rect 8110 14764 8116 14776
rect 8168 14764 8174 14816
rect 8662 14764 8668 14816
rect 8720 14804 8726 14816
rect 9125 14807 9183 14813
rect 9125 14804 9137 14807
rect 8720 14776 9137 14804
rect 8720 14764 8726 14776
rect 9125 14773 9137 14776
rect 9171 14773 9183 14807
rect 9125 14767 9183 14773
rect 9306 14764 9312 14816
rect 9364 14804 9370 14816
rect 10134 14804 10140 14816
rect 9364 14776 10140 14804
rect 9364 14764 9370 14776
rect 10134 14764 10140 14776
rect 10192 14804 10198 14816
rect 10321 14807 10379 14813
rect 10321 14804 10333 14807
rect 10192 14776 10333 14804
rect 10192 14764 10198 14776
rect 10321 14773 10333 14776
rect 10367 14773 10379 14807
rect 10321 14767 10379 14773
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 11072 14804 11100 14844
rect 13081 14841 13093 14844
rect 13127 14841 13139 14875
rect 13081 14835 13139 14841
rect 10652 14776 11100 14804
rect 11425 14807 11483 14813
rect 10652 14764 10658 14776
rect 11425 14773 11437 14807
rect 11471 14804 11483 14807
rect 11698 14804 11704 14816
rect 11471 14776 11704 14804
rect 11471 14773 11483 14776
rect 11425 14767 11483 14773
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 14366 14804 14372 14816
rect 12492 14776 12537 14804
rect 14327 14776 14372 14804
rect 12492 14764 12498 14776
rect 14366 14764 14372 14776
rect 14424 14764 14430 14816
rect 1104 14714 15824 14736
rect 1104 14662 5912 14714
rect 5964 14662 5976 14714
rect 6028 14662 6040 14714
rect 6092 14662 6104 14714
rect 6156 14662 10843 14714
rect 10895 14662 10907 14714
rect 10959 14662 10971 14714
rect 11023 14662 11035 14714
rect 11087 14662 15824 14714
rect 1104 14640 15824 14662
rect 6638 14600 6644 14612
rect 3068 14572 6644 14600
rect 2133 14535 2191 14541
rect 2133 14501 2145 14535
rect 2179 14532 2191 14535
rect 2774 14532 2780 14544
rect 2179 14504 2780 14532
rect 2179 14501 2191 14504
rect 2133 14495 2191 14501
rect 2774 14492 2780 14504
rect 2832 14492 2838 14544
rect 1857 14467 1915 14473
rect 1857 14433 1869 14467
rect 1903 14464 1915 14467
rect 3068 14464 3096 14572
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 7009 14603 7067 14609
rect 7009 14569 7021 14603
rect 7055 14600 7067 14603
rect 7466 14600 7472 14612
rect 7055 14572 7472 14600
rect 7055 14569 7067 14572
rect 7009 14563 7067 14569
rect 7466 14560 7472 14572
rect 7524 14560 7530 14612
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 8849 14603 8907 14609
rect 8849 14600 8861 14603
rect 7616 14572 8861 14600
rect 7616 14560 7622 14572
rect 8849 14569 8861 14572
rect 8895 14569 8907 14603
rect 8849 14563 8907 14569
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 9677 14603 9735 14609
rect 9677 14600 9689 14603
rect 9640 14572 9689 14600
rect 9640 14560 9646 14572
rect 9677 14569 9689 14572
rect 9723 14569 9735 14603
rect 10873 14603 10931 14609
rect 10873 14600 10885 14603
rect 9677 14563 9735 14569
rect 10244 14572 10885 14600
rect 3145 14535 3203 14541
rect 3145 14501 3157 14535
rect 3191 14532 3203 14535
rect 3191 14504 5488 14532
rect 3191 14501 3203 14504
rect 3145 14495 3203 14501
rect 1903 14436 3096 14464
rect 3237 14467 3295 14473
rect 1903 14433 1915 14436
rect 1857 14427 1915 14433
rect 3237 14433 3249 14467
rect 3283 14464 3295 14467
rect 4798 14464 4804 14476
rect 3283 14436 4016 14464
rect 4759 14436 4804 14464
rect 3283 14433 3295 14436
rect 3237 14427 3295 14433
rect 3418 14396 3424 14408
rect 3379 14368 3424 14396
rect 3418 14356 3424 14368
rect 3476 14356 3482 14408
rect 3988 14396 4016 14436
rect 4798 14424 4804 14436
rect 4856 14424 4862 14476
rect 4890 14424 4896 14476
rect 4948 14464 4954 14476
rect 5460 14464 5488 14504
rect 5534 14492 5540 14544
rect 5592 14532 5598 14544
rect 5874 14535 5932 14541
rect 5874 14532 5886 14535
rect 5592 14504 5886 14532
rect 5592 14492 5598 14504
rect 5874 14501 5886 14504
rect 5920 14532 5932 14535
rect 6270 14532 6276 14544
rect 5920 14504 6276 14532
rect 5920 14501 5932 14504
rect 5874 14495 5932 14501
rect 6270 14492 6276 14504
rect 6328 14492 6334 14544
rect 6822 14492 6828 14544
rect 6880 14532 6886 14544
rect 10244 14532 10272 14572
rect 10873 14569 10885 14572
rect 10919 14569 10931 14603
rect 10873 14563 10931 14569
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13320 14572 14105 14600
rect 13320 14560 13326 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 14093 14563 14151 14569
rect 11333 14535 11391 14541
rect 11333 14532 11345 14535
rect 6880 14504 10272 14532
rect 10612 14504 11345 14532
rect 6880 14492 6886 14504
rect 7558 14464 7564 14476
rect 4948 14436 4993 14464
rect 5460 14436 7564 14464
rect 4948 14424 4954 14436
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 7742 14473 7748 14476
rect 7736 14464 7748 14473
rect 7703 14436 7748 14464
rect 7736 14427 7748 14436
rect 7742 14424 7748 14427
rect 7800 14424 7806 14476
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 9493 14467 9551 14473
rect 8352 14436 8524 14464
rect 8352 14424 8358 14436
rect 5077 14399 5135 14405
rect 3988 14368 5028 14396
rect 2777 14331 2835 14337
rect 2777 14297 2789 14331
rect 2823 14328 2835 14331
rect 4706 14328 4712 14340
rect 2823 14300 4712 14328
rect 2823 14297 2835 14300
rect 2777 14291 2835 14297
rect 4706 14288 4712 14300
rect 4764 14288 4770 14340
rect 5000 14328 5028 14368
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5534 14396 5540 14408
rect 5123 14368 5540 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 5626 14356 5632 14408
rect 5684 14396 5690 14408
rect 5684 14368 5729 14396
rect 5684 14356 5690 14368
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 7469 14399 7527 14405
rect 7469 14396 7481 14399
rect 6880 14368 7481 14396
rect 6880 14356 6886 14368
rect 7469 14365 7481 14368
rect 7515 14365 7527 14399
rect 8496 14396 8524 14436
rect 9493 14433 9505 14467
rect 9539 14464 9551 14467
rect 9582 14464 9588 14476
rect 9539 14436 9588 14464
rect 9539 14433 9551 14436
rect 9493 14427 9551 14433
rect 9582 14424 9588 14436
rect 9640 14424 9646 14476
rect 10042 14464 10048 14476
rect 10003 14436 10048 14464
rect 10042 14424 10048 14436
rect 10100 14464 10106 14476
rect 10612 14464 10640 14504
rect 11333 14501 11345 14504
rect 11379 14501 11391 14535
rect 11333 14495 11391 14501
rect 10100 14436 10640 14464
rect 10100 14424 10106 14436
rect 11146 14424 11152 14476
rect 11204 14464 11210 14476
rect 11241 14467 11299 14473
rect 11241 14464 11253 14467
rect 11204 14436 11253 14464
rect 11204 14424 11210 14436
rect 11241 14433 11253 14436
rect 11287 14433 11299 14467
rect 11241 14427 11299 14433
rect 11790 14424 11796 14476
rect 11848 14464 11854 14476
rect 12069 14467 12127 14473
rect 12069 14464 12081 14467
rect 11848 14436 12081 14464
rect 11848 14424 11854 14436
rect 12069 14433 12081 14436
rect 12115 14433 12127 14467
rect 12069 14427 12127 14433
rect 12710 14424 12716 14476
rect 12768 14464 12774 14476
rect 13357 14467 13415 14473
rect 13357 14464 13369 14467
rect 12768 14436 13369 14464
rect 12768 14424 12774 14436
rect 13357 14433 13369 14436
rect 13403 14464 13415 14467
rect 13630 14464 13636 14476
rect 13403 14436 13636 14464
rect 13403 14433 13415 14436
rect 13357 14427 13415 14433
rect 13630 14424 13636 14436
rect 13688 14424 13694 14476
rect 9858 14396 9864 14408
rect 8496 14368 9864 14396
rect 7469 14359 7527 14365
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 10134 14396 10140 14408
rect 10095 14368 10140 14396
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 5000 14300 5672 14328
rect 1670 14220 1676 14272
rect 1728 14260 1734 14272
rect 4246 14260 4252 14272
rect 1728 14232 4252 14260
rect 1728 14220 1734 14232
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 4430 14260 4436 14272
rect 4391 14232 4436 14260
rect 4430 14220 4436 14232
rect 4488 14220 4494 14272
rect 5644 14260 5672 14300
rect 8662 14288 8668 14340
rect 8720 14328 8726 14340
rect 8938 14328 8944 14340
rect 8720 14300 8944 14328
rect 8720 14288 8726 14300
rect 8938 14288 8944 14300
rect 8996 14288 9002 14340
rect 9214 14288 9220 14340
rect 9272 14328 9278 14340
rect 10244 14328 10272 14359
rect 10962 14356 10968 14408
rect 11020 14396 11026 14408
rect 11425 14399 11483 14405
rect 11425 14396 11437 14399
rect 11020 14368 11437 14396
rect 11020 14356 11026 14368
rect 11425 14365 11437 14368
rect 11471 14365 11483 14399
rect 11425 14359 11483 14365
rect 12253 14399 12311 14405
rect 12253 14365 12265 14399
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 9272 14300 10272 14328
rect 9272 14288 9278 14300
rect 10686 14288 10692 14340
rect 10744 14328 10750 14340
rect 12268 14328 12296 14359
rect 10744 14300 12296 14328
rect 10744 14288 10750 14300
rect 8754 14260 8760 14272
rect 5644 14232 8760 14260
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 9309 14263 9367 14269
rect 9309 14229 9321 14263
rect 9355 14260 9367 14263
rect 9398 14260 9404 14272
rect 9355 14232 9404 14260
rect 9355 14229 9367 14232
rect 9309 14223 9367 14229
rect 9398 14220 9404 14232
rect 9456 14220 9462 14272
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 11698 14260 11704 14272
rect 9916 14232 11704 14260
rect 9916 14220 9922 14232
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 13541 14263 13599 14269
rect 13541 14229 13553 14263
rect 13587 14260 13599 14263
rect 15010 14260 15016 14272
rect 13587 14232 15016 14260
rect 13587 14229 13599 14232
rect 13541 14223 13599 14229
rect 15010 14220 15016 14232
rect 15068 14220 15074 14272
rect 1104 14170 15824 14192
rect 1104 14118 3447 14170
rect 3499 14118 3511 14170
rect 3563 14118 3575 14170
rect 3627 14118 3639 14170
rect 3691 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 13308 14170
rect 13360 14118 13372 14170
rect 13424 14118 13436 14170
rect 13488 14118 13500 14170
rect 13552 14118 15824 14170
rect 1104 14096 15824 14118
rect 2501 14059 2559 14065
rect 2501 14025 2513 14059
rect 2547 14056 2559 14059
rect 3326 14056 3332 14068
rect 2547 14028 3332 14056
rect 2547 14025 2559 14028
rect 2501 14019 2559 14025
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 3697 14059 3755 14065
rect 3697 14025 3709 14059
rect 3743 14056 3755 14059
rect 4798 14056 4804 14068
rect 3743 14028 4804 14056
rect 3743 14025 3755 14028
rect 3697 14019 3755 14025
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 5166 14056 5172 14068
rect 4908 14028 5172 14056
rect 4908 13988 4936 14028
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 6270 14056 6276 14068
rect 6231 14028 6276 14056
rect 6270 14016 6276 14028
rect 6328 14016 6334 14068
rect 7558 14016 7564 14068
rect 7616 14056 7622 14068
rect 7616 14028 9628 14056
rect 7616 14016 7622 14028
rect 2976 13960 4936 13988
rect 2976 13929 3004 13960
rect 7926 13948 7932 14000
rect 7984 13988 7990 14000
rect 8205 13991 8263 13997
rect 8205 13988 8217 13991
rect 7984 13960 8217 13988
rect 7984 13948 7990 13960
rect 8205 13957 8217 13960
rect 8251 13957 8263 13991
rect 9600 13988 9628 14028
rect 10134 14016 10140 14068
rect 10192 14056 10198 14068
rect 10505 14059 10563 14065
rect 10505 14056 10517 14059
rect 10192 14028 10517 14056
rect 10192 14016 10198 14028
rect 10505 14025 10517 14028
rect 10551 14025 10563 14059
rect 10505 14019 10563 14025
rect 10686 14016 10692 14068
rect 10744 14056 10750 14068
rect 11054 14056 11060 14068
rect 10744 14028 11060 14056
rect 10744 14016 10750 14028
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 12437 13991 12495 13997
rect 9600 13960 11192 13988
rect 8205 13951 8263 13957
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13889 3019 13923
rect 2961 13883 3019 13889
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 4246 13920 4252 13932
rect 3191 13892 4252 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4522 13920 4528 13932
rect 4387 13892 4528 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 6822 13920 6828 13932
rect 6783 13892 6828 13920
rect 6822 13880 6828 13892
rect 6880 13880 6886 13932
rect 8110 13880 8116 13932
rect 8168 13920 8174 13932
rect 8168 13892 8800 13920
rect 8168 13880 8174 13892
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13852 1915 13855
rect 2498 13852 2504 13864
rect 1903 13824 2504 13852
rect 1903 13821 1915 13824
rect 1857 13815 1915 13821
rect 2498 13812 2504 13824
rect 2556 13812 2562 13864
rect 4157 13855 4215 13861
rect 4157 13821 4169 13855
rect 4203 13852 4215 13855
rect 4893 13855 4951 13861
rect 4203 13824 4844 13852
rect 4203 13821 4215 13824
rect 4157 13815 4215 13821
rect 4816 13784 4844 13824
rect 4893 13821 4905 13855
rect 4939 13852 4951 13855
rect 4982 13852 4988 13864
rect 4939 13824 4988 13852
rect 4939 13821 4951 13824
rect 4893 13815 4951 13821
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 6730 13852 6736 13864
rect 5092 13824 6736 13852
rect 5092 13784 5120 13824
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 7092 13855 7150 13861
rect 7092 13821 7104 13855
rect 7138 13852 7150 13855
rect 7466 13852 7472 13864
rect 7138 13824 7472 13852
rect 7138 13821 7150 13824
rect 7092 13815 7150 13821
rect 7466 13812 7472 13824
rect 7524 13812 7530 13864
rect 8662 13852 8668 13864
rect 7567 13824 8668 13852
rect 4816 13756 5120 13784
rect 5160 13787 5218 13793
rect 5160 13753 5172 13787
rect 5206 13784 5218 13787
rect 5258 13784 5264 13796
rect 5206 13756 5264 13784
rect 5206 13753 5218 13756
rect 5160 13747 5218 13753
rect 5258 13744 5264 13756
rect 5316 13784 5322 13796
rect 6362 13784 6368 13796
rect 5316 13756 6368 13784
rect 5316 13744 5322 13756
rect 6362 13744 6368 13756
rect 6420 13744 6426 13796
rect 6822 13744 6828 13796
rect 6880 13784 6886 13796
rect 7567 13784 7595 13824
rect 8662 13812 8668 13824
rect 8720 13812 8726 13864
rect 8772 13852 8800 13892
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 9950 13920 9956 13932
rect 9732 13892 9956 13920
rect 9732 13880 9738 13892
rect 9950 13880 9956 13892
rect 10008 13920 10014 13932
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 10008 13892 10977 13920
rect 10008 13880 10014 13892
rect 10965 13889 10977 13892
rect 11011 13889 11023 13923
rect 10965 13883 11023 13889
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13889 11115 13923
rect 11164 13920 11192 13960
rect 12437 13957 12449 13991
rect 12483 13957 12495 13991
rect 12437 13951 12495 13957
rect 14001 13991 14059 13997
rect 14001 13957 14013 13991
rect 14047 13988 14059 13991
rect 14918 13988 14924 14000
rect 14047 13960 14924 13988
rect 14047 13957 14059 13960
rect 14001 13951 14059 13957
rect 12452 13920 12480 13951
rect 14918 13948 14924 13960
rect 14976 13948 14982 14000
rect 11164 13892 12480 13920
rect 13081 13923 13139 13929
rect 11057 13883 11115 13889
rect 13081 13889 13093 13923
rect 13127 13920 13139 13923
rect 13262 13920 13268 13932
rect 13127 13892 13268 13920
rect 13127 13889 13139 13892
rect 13081 13883 13139 13889
rect 8921 13855 8979 13861
rect 8921 13852 8933 13855
rect 8772 13824 8933 13852
rect 8921 13821 8933 13824
rect 8967 13821 8979 13855
rect 11072 13852 11100 13883
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 8921 13815 8979 13821
rect 9692 13824 11100 13852
rect 6880 13756 7595 13784
rect 6880 13744 6886 13756
rect 8110 13744 8116 13796
rect 8168 13784 8174 13796
rect 9692 13784 9720 13824
rect 12342 13812 12348 13864
rect 12400 13852 12406 13864
rect 12710 13852 12716 13864
rect 12400 13824 12716 13852
rect 12400 13812 12406 13824
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 13814 13852 13820 13864
rect 13775 13824 13820 13852
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 14182 13812 14188 13864
rect 14240 13852 14246 13864
rect 14458 13852 14464 13864
rect 14240 13824 14464 13852
rect 14240 13812 14246 13824
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 8168 13756 9720 13784
rect 8168 13744 8174 13756
rect 10318 13744 10324 13796
rect 10376 13784 10382 13796
rect 10870 13784 10876 13796
rect 10376 13756 10876 13784
rect 10376 13744 10382 13756
rect 10870 13744 10876 13756
rect 10928 13744 10934 13796
rect 10962 13744 10968 13796
rect 11020 13744 11026 13796
rect 12805 13787 12863 13793
rect 12805 13753 12817 13787
rect 12851 13784 12863 13787
rect 14553 13787 14611 13793
rect 14553 13784 14565 13787
rect 12851 13756 14565 13784
rect 12851 13753 12863 13756
rect 12805 13747 12863 13753
rect 14553 13753 14565 13756
rect 14599 13753 14611 13787
rect 14553 13747 14611 13753
rect 2869 13719 2927 13725
rect 2869 13685 2881 13719
rect 2915 13716 2927 13719
rect 2958 13716 2964 13728
rect 2915 13688 2964 13716
rect 2915 13685 2927 13688
rect 2869 13679 2927 13685
rect 2958 13676 2964 13688
rect 3016 13676 3022 13728
rect 4065 13719 4123 13725
rect 4065 13685 4077 13719
rect 4111 13716 4123 13719
rect 7650 13716 7656 13728
rect 4111 13688 7656 13716
rect 4111 13685 4123 13688
rect 4065 13679 4123 13685
rect 7650 13676 7656 13688
rect 7708 13676 7714 13728
rect 8386 13676 8392 13728
rect 8444 13716 8450 13728
rect 9582 13716 9588 13728
rect 8444 13688 9588 13716
rect 8444 13676 8450 13688
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 10045 13719 10103 13725
rect 10045 13716 10057 13719
rect 9824 13688 10057 13716
rect 9824 13676 9830 13688
rect 10045 13685 10057 13688
rect 10091 13716 10103 13719
rect 10980 13716 11008 13744
rect 10091 13688 11008 13716
rect 10091 13685 10103 13688
rect 10045 13679 10103 13685
rect 11146 13676 11152 13728
rect 11204 13716 11210 13728
rect 11701 13719 11759 13725
rect 11701 13716 11713 13719
rect 11204 13688 11713 13716
rect 11204 13676 11210 13688
rect 11701 13685 11713 13688
rect 11747 13685 11759 13719
rect 12894 13716 12900 13728
rect 12807 13688 12900 13716
rect 11701 13679 11759 13685
rect 12894 13676 12900 13688
rect 12952 13716 12958 13728
rect 15286 13716 15292 13728
rect 12952 13688 15292 13716
rect 12952 13676 12958 13688
rect 15286 13676 15292 13688
rect 15344 13716 15350 13728
rect 15746 13716 15752 13728
rect 15344 13688 15752 13716
rect 15344 13676 15350 13688
rect 15746 13676 15752 13688
rect 15804 13676 15810 13728
rect 1104 13626 15824 13648
rect 1104 13574 5912 13626
rect 5964 13574 5976 13626
rect 6028 13574 6040 13626
rect 6092 13574 6104 13626
rect 6156 13574 10843 13626
rect 10895 13574 10907 13626
rect 10959 13574 10971 13626
rect 11023 13574 11035 13626
rect 11087 13574 15824 13626
rect 1104 13552 15824 13574
rect 1581 13515 1639 13521
rect 1581 13481 1593 13515
rect 1627 13512 1639 13515
rect 1670 13512 1676 13524
rect 1627 13484 1676 13512
rect 1627 13481 1639 13484
rect 1581 13475 1639 13481
rect 1670 13472 1676 13484
rect 1728 13472 1734 13524
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 1995 13484 2912 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 2041 13379 2099 13385
rect 2041 13345 2053 13379
rect 2087 13376 2099 13379
rect 2682 13376 2688 13388
rect 2087 13348 2688 13376
rect 2087 13345 2099 13348
rect 2041 13339 2099 13345
rect 2682 13336 2688 13348
rect 2740 13336 2746 13388
rect 2884 13376 2912 13484
rect 2958 13472 2964 13524
rect 3016 13512 3022 13524
rect 4798 13512 4804 13524
rect 3016 13484 4804 13512
rect 3016 13472 3022 13484
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 6730 13472 6736 13524
rect 6788 13512 6794 13524
rect 8021 13515 8079 13521
rect 8021 13512 8033 13515
rect 6788 13484 8033 13512
rect 6788 13472 6794 13484
rect 8021 13481 8033 13484
rect 8067 13481 8079 13515
rect 8386 13512 8392 13524
rect 8347 13484 8392 13512
rect 8021 13475 8079 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8662 13472 8668 13524
rect 8720 13512 8726 13524
rect 9493 13515 9551 13521
rect 9493 13512 9505 13515
rect 8720 13484 9505 13512
rect 8720 13472 8726 13484
rect 9493 13481 9505 13484
rect 9539 13481 9551 13515
rect 9493 13475 9551 13481
rect 9582 13472 9588 13524
rect 9640 13512 9646 13524
rect 10686 13512 10692 13524
rect 9640 13484 10692 13512
rect 9640 13472 9646 13484
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 11698 13472 11704 13524
rect 11756 13512 11762 13524
rect 12713 13515 12771 13521
rect 12713 13512 12725 13515
rect 11756 13484 12725 13512
rect 11756 13472 11762 13484
rect 12713 13481 12725 13484
rect 12759 13481 12771 13515
rect 13078 13512 13084 13524
rect 13039 13484 13084 13512
rect 12713 13475 12771 13481
rect 13078 13472 13084 13484
rect 13136 13472 13142 13524
rect 13170 13472 13176 13524
rect 13228 13512 13234 13524
rect 13228 13484 13273 13512
rect 13228 13472 13234 13484
rect 3145 13447 3203 13453
rect 3145 13413 3157 13447
rect 3191 13444 3203 13447
rect 3326 13444 3332 13456
rect 3191 13416 3332 13444
rect 3191 13413 3203 13416
rect 3145 13407 3203 13413
rect 3326 13404 3332 13416
rect 3384 13404 3390 13456
rect 5442 13444 5448 13456
rect 3436 13416 5448 13444
rect 2884 13348 3372 13376
rect 2222 13308 2228 13320
rect 2183 13280 2228 13308
rect 2222 13268 2228 13280
rect 2280 13268 2286 13320
rect 2774 13268 2780 13320
rect 2832 13308 2838 13320
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 2832 13280 3249 13308
rect 2832 13268 2838 13280
rect 3237 13277 3249 13280
rect 3283 13277 3295 13311
rect 3237 13271 3295 13277
rect 2777 13175 2835 13181
rect 2777 13141 2789 13175
rect 2823 13172 2835 13175
rect 3142 13172 3148 13184
rect 2823 13144 3148 13172
rect 2823 13141 2835 13144
rect 2777 13135 2835 13141
rect 3142 13132 3148 13144
rect 3200 13132 3206 13184
rect 3344 13172 3372 13348
rect 3436 13317 3464 13416
rect 5442 13404 5448 13416
rect 5500 13404 5506 13456
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 6270 13444 6276 13456
rect 5592 13416 6276 13444
rect 5592 13404 5598 13416
rect 6270 13404 6276 13416
rect 6328 13444 6334 13456
rect 6426 13447 6484 13453
rect 6426 13444 6438 13447
rect 6328 13416 6438 13444
rect 6328 13404 6334 13416
rect 6426 13413 6438 13416
rect 6472 13413 6484 13447
rect 6426 13407 6484 13413
rect 6914 13404 6920 13456
rect 6972 13444 6978 13456
rect 6972 13416 9536 13444
rect 6972 13404 6978 13416
rect 3786 13336 3792 13388
rect 3844 13376 3850 13388
rect 4341 13379 4399 13385
rect 4341 13376 4353 13379
rect 3844 13348 4353 13376
rect 3844 13336 3850 13348
rect 4341 13345 4353 13348
rect 4387 13345 4399 13379
rect 4341 13339 4399 13345
rect 4608 13379 4666 13385
rect 4608 13345 4620 13379
rect 4654 13376 4666 13379
rect 5810 13376 5816 13388
rect 4654 13348 5816 13376
rect 4654 13345 4666 13348
rect 4608 13339 4666 13345
rect 5810 13336 5816 13348
rect 5868 13336 5874 13388
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13376 6239 13379
rect 6822 13376 6828 13388
rect 6227 13348 6828 13376
rect 6227 13345 6239 13348
rect 6181 13339 6239 13345
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 7282 13336 7288 13388
rect 7340 13376 7346 13388
rect 7650 13376 7656 13388
rect 7340 13348 7656 13376
rect 7340 13336 7346 13348
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 8481 13379 8539 13385
rect 8481 13345 8493 13379
rect 8527 13376 8539 13379
rect 9398 13376 9404 13388
rect 8527 13348 9260 13376
rect 9359 13348 9404 13376
rect 8527 13345 8539 13348
rect 8481 13339 8539 13345
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 8018 13268 8024 13320
rect 8076 13308 8082 13320
rect 8665 13311 8723 13317
rect 8665 13308 8677 13311
rect 8076 13280 8677 13308
rect 8076 13268 8082 13280
rect 8665 13277 8677 13280
rect 8711 13308 8723 13311
rect 9122 13308 9128 13320
rect 8711 13280 9128 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 9232 13308 9260 13348
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 9508 13376 9536 13416
rect 9674 13404 9680 13456
rect 9732 13444 9738 13456
rect 9732 13416 10088 13444
rect 9732 13404 9738 13416
rect 9766 13376 9772 13388
rect 9508 13348 9772 13376
rect 9766 13336 9772 13348
rect 9824 13376 9830 13388
rect 9933 13379 9991 13385
rect 9933 13376 9945 13379
rect 9824 13348 9945 13376
rect 9824 13336 9830 13348
rect 9933 13345 9945 13348
rect 9979 13345 9991 13379
rect 10060 13376 10088 13416
rect 10134 13404 10140 13456
rect 10192 13444 10198 13456
rect 14185 13447 14243 13453
rect 14185 13444 14197 13447
rect 10192 13416 14197 13444
rect 10192 13404 10198 13416
rect 14185 13413 14197 13416
rect 14231 13413 14243 13447
rect 14185 13407 14243 13413
rect 10060 13348 10732 13376
rect 9933 13339 9991 13345
rect 9493 13311 9551 13317
rect 9232 13280 9444 13308
rect 5626 13200 5632 13252
rect 5684 13240 5690 13252
rect 5721 13243 5779 13249
rect 5721 13240 5733 13243
rect 5684 13212 5733 13240
rect 5684 13200 5690 13212
rect 5721 13209 5733 13212
rect 5767 13209 5779 13243
rect 5721 13203 5779 13209
rect 7466 13200 7472 13252
rect 7524 13240 7530 13252
rect 9217 13243 9275 13249
rect 7524 13212 8892 13240
rect 7524 13200 7530 13212
rect 7098 13172 7104 13184
rect 3344 13144 7104 13172
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 7558 13172 7564 13184
rect 7519 13144 7564 13172
rect 7558 13132 7564 13144
rect 7616 13132 7622 13184
rect 8864 13172 8892 13212
rect 9217 13209 9229 13243
rect 9263 13240 9275 13243
rect 9306 13240 9312 13252
rect 9263 13212 9312 13240
rect 9263 13209 9275 13212
rect 9217 13203 9275 13209
rect 9306 13200 9312 13212
rect 9364 13200 9370 13252
rect 9416 13240 9444 13280
rect 9493 13277 9505 13311
rect 9539 13308 9551 13311
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9539 13280 9689 13308
rect 9539 13277 9551 13280
rect 9493 13271 9551 13277
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 10704 13308 10732 13348
rect 10962 13336 10968 13388
rect 11020 13376 11026 13388
rect 11020 13348 11652 13376
rect 11020 13336 11026 13348
rect 10704 13280 11192 13308
rect 9677 13271 9735 13277
rect 9416 13212 9720 13240
rect 9692 13184 9720 13212
rect 10962 13200 10968 13252
rect 11020 13200 11026 13252
rect 11164 13240 11192 13280
rect 11517 13243 11575 13249
rect 11517 13240 11529 13243
rect 11164 13212 11529 13240
rect 11517 13209 11529 13212
rect 11563 13209 11575 13243
rect 11624 13240 11652 13348
rect 11698 13336 11704 13388
rect 11756 13376 11762 13388
rect 11885 13379 11943 13385
rect 11885 13376 11897 13379
rect 11756 13348 11897 13376
rect 11756 13336 11762 13348
rect 11885 13345 11897 13348
rect 11931 13345 11943 13379
rect 11885 13339 11943 13345
rect 11977 13379 12035 13385
rect 11977 13345 11989 13379
rect 12023 13376 12035 13379
rect 12526 13376 12532 13388
rect 12023 13348 12532 13376
rect 12023 13345 12035 13348
rect 11977 13339 12035 13345
rect 12526 13336 12532 13348
rect 12584 13376 12590 13388
rect 13906 13376 13912 13388
rect 12584 13348 13584 13376
rect 13867 13348 13912 13376
rect 12584 13336 12590 13348
rect 11790 13268 11796 13320
rect 11848 13308 11854 13320
rect 12069 13311 12127 13317
rect 12069 13308 12081 13311
rect 11848 13280 12081 13308
rect 11848 13268 11854 13280
rect 12069 13277 12081 13280
rect 12115 13308 12127 13311
rect 12250 13308 12256 13320
rect 12115 13280 12256 13308
rect 12115 13277 12127 13280
rect 12069 13271 12127 13277
rect 12250 13268 12256 13280
rect 12308 13268 12314 13320
rect 13262 13308 13268 13320
rect 13175 13280 13268 13308
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 13556 13308 13584 13348
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 14458 13308 14464 13320
rect 13556 13280 14464 13308
rect 14458 13268 14464 13280
rect 14516 13308 14522 13320
rect 15378 13308 15384 13320
rect 14516 13280 15384 13308
rect 14516 13268 14522 13280
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 13280 13240 13308 13268
rect 11624 13212 13308 13240
rect 11517 13203 11575 13209
rect 9398 13172 9404 13184
rect 8864 13144 9404 13172
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 9674 13132 9680 13184
rect 9732 13132 9738 13184
rect 10980 13172 11008 13200
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 10980 13144 11069 13172
rect 11057 13141 11069 13144
rect 11103 13141 11115 13175
rect 11057 13135 11115 13141
rect 1104 13082 15824 13104
rect 1104 13030 3447 13082
rect 3499 13030 3511 13082
rect 3563 13030 3575 13082
rect 3627 13030 3639 13082
rect 3691 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 13308 13082
rect 13360 13030 13372 13082
rect 13424 13030 13436 13082
rect 13488 13030 13500 13082
rect 13552 13030 15824 13082
rect 1104 13008 15824 13030
rect 6270 12968 6276 12980
rect 2516 12940 4476 12968
rect 2516 12841 2544 12940
rect 4448 12900 4476 12940
rect 4908 12940 6132 12968
rect 6231 12940 6276 12968
rect 4908 12900 4936 12940
rect 4448 12872 4936 12900
rect 6104 12900 6132 12940
rect 6270 12928 6276 12940
rect 6328 12928 6334 12980
rect 6840 12940 7972 12968
rect 6546 12900 6552 12912
rect 6104 12872 6552 12900
rect 6546 12860 6552 12872
rect 6604 12860 6610 12912
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12801 2559 12835
rect 2501 12795 2559 12801
rect 6638 12792 6644 12844
rect 6696 12832 6702 12844
rect 6840 12841 6868 12940
rect 7944 12900 7972 12940
rect 8018 12928 8024 12980
rect 8076 12968 8082 12980
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 8076 12940 8217 12968
rect 8076 12928 8082 12940
rect 8205 12937 8217 12940
rect 8251 12937 8263 12971
rect 13633 12971 13691 12977
rect 13633 12968 13645 12971
rect 8205 12931 8263 12937
rect 8312 12940 13645 12968
rect 8312 12900 8340 12940
rect 13633 12937 13645 12940
rect 13679 12937 13691 12971
rect 13633 12931 13691 12937
rect 7944 12872 8340 12900
rect 9858 12860 9864 12912
rect 9916 12900 9922 12912
rect 10045 12903 10103 12909
rect 10045 12900 10057 12903
rect 9916 12872 10057 12900
rect 9916 12860 9922 12872
rect 10045 12869 10057 12872
rect 10091 12869 10103 12903
rect 10045 12863 10103 12869
rect 10134 12860 10140 12912
rect 10192 12900 10198 12912
rect 10962 12900 10968 12912
rect 10192 12872 10968 12900
rect 10192 12860 10198 12872
rect 10962 12860 10968 12872
rect 11020 12860 11026 12912
rect 13262 12900 13268 12912
rect 11072 12872 13268 12900
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6696 12804 6837 12832
rect 6696 12792 6702 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 8662 12832 8668 12844
rect 8623 12804 8668 12832
rect 6825 12795 6883 12801
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 9674 12792 9680 12844
rect 9732 12832 9738 12844
rect 11072 12832 11100 12872
rect 13262 12860 13268 12872
rect 13320 12860 13326 12912
rect 9732 12804 11100 12832
rect 11149 12835 11207 12841
rect 9732 12792 9738 12804
rect 11149 12801 11161 12835
rect 11195 12801 11207 12835
rect 11698 12832 11704 12844
rect 11659 12804 11704 12832
rect 11149 12795 11207 12801
rect 3053 12767 3111 12773
rect 3053 12733 3065 12767
rect 3099 12764 3111 12767
rect 3694 12764 3700 12776
rect 3099 12736 3700 12764
rect 3099 12733 3111 12736
rect 3053 12727 3111 12733
rect 3694 12724 3700 12736
rect 3752 12764 3758 12776
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 3752 12736 4905 12764
rect 3752 12724 3758 12736
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 4893 12727 4951 12733
rect 5000 12736 5396 12764
rect 3142 12696 3148 12708
rect 1872 12668 3148 12696
rect 1872 12637 1900 12668
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 3320 12699 3378 12705
rect 3320 12665 3332 12699
rect 3366 12696 3378 12699
rect 3786 12696 3792 12708
rect 3366 12668 3792 12696
rect 3366 12665 3378 12668
rect 3320 12659 3378 12665
rect 3786 12656 3792 12668
rect 3844 12656 3850 12708
rect 5000 12696 5028 12736
rect 5166 12705 5172 12708
rect 5160 12696 5172 12705
rect 4356 12668 5028 12696
rect 5127 12668 5172 12696
rect 1857 12631 1915 12637
rect 1857 12597 1869 12631
rect 1903 12597 1915 12631
rect 2222 12628 2228 12640
rect 2183 12600 2228 12628
rect 1857 12591 1915 12597
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 2317 12631 2375 12637
rect 2317 12597 2329 12631
rect 2363 12628 2375 12631
rect 4356 12628 4384 12668
rect 5160 12659 5172 12668
rect 5166 12656 5172 12659
rect 5224 12656 5230 12708
rect 2363 12600 4384 12628
rect 4433 12631 4491 12637
rect 2363 12597 2375 12600
rect 2317 12591 2375 12597
rect 4433 12597 4445 12631
rect 4479 12628 4491 12631
rect 5258 12628 5264 12640
rect 4479 12600 5264 12628
rect 4479 12597 4491 12600
rect 4433 12591 4491 12597
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5368 12628 5396 12736
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 7092 12767 7150 12773
rect 7092 12764 7104 12767
rect 6972 12736 7104 12764
rect 6972 12724 6978 12736
rect 7092 12733 7104 12736
rect 7138 12764 7150 12767
rect 8110 12764 8116 12776
rect 7138 12736 8116 12764
rect 7138 12733 7150 12736
rect 7092 12727 7150 12733
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 8570 12724 8576 12776
rect 8628 12764 8634 12776
rect 10042 12764 10048 12776
rect 8628 12736 10048 12764
rect 8628 12724 8634 12736
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10873 12767 10931 12773
rect 10873 12764 10885 12767
rect 10152 12736 10885 12764
rect 7650 12656 7656 12708
rect 7708 12696 7714 12708
rect 7708 12668 7880 12696
rect 7708 12656 7714 12668
rect 7742 12628 7748 12640
rect 5368 12600 7748 12628
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 7852 12628 7880 12668
rect 7926 12656 7932 12708
rect 7984 12696 7990 12708
rect 8932 12699 8990 12705
rect 8932 12696 8944 12699
rect 7984 12668 8944 12696
rect 7984 12656 7990 12668
rect 8932 12665 8944 12668
rect 8978 12696 8990 12699
rect 9490 12696 9496 12708
rect 8978 12668 9496 12696
rect 8978 12665 8990 12668
rect 8932 12659 8990 12665
rect 9490 12656 9496 12668
rect 9548 12656 9554 12708
rect 9674 12656 9680 12708
rect 9732 12696 9738 12708
rect 10152 12696 10180 12736
rect 10873 12733 10885 12736
rect 10919 12733 10931 12767
rect 10873 12727 10931 12733
rect 9732 12668 10180 12696
rect 9732 12656 9738 12668
rect 10778 12656 10784 12708
rect 10836 12696 10842 12708
rect 10965 12699 11023 12705
rect 10965 12696 10977 12699
rect 10836 12668 10977 12696
rect 10836 12656 10842 12668
rect 10965 12665 10977 12668
rect 11011 12665 11023 12699
rect 10965 12659 11023 12665
rect 10134 12628 10140 12640
rect 7852 12600 10140 12628
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 10505 12631 10563 12637
rect 10505 12597 10517 12631
rect 10551 12628 10563 12631
rect 10594 12628 10600 12640
rect 10551 12600 10600 12628
rect 10551 12597 10563 12600
rect 10505 12591 10563 12597
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 11164 12628 11192 12795
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 12250 12792 12256 12844
rect 12308 12832 12314 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12308 12804 13001 12832
rect 12308 12792 12314 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13630 12792 13636 12844
rect 13688 12832 13694 12844
rect 13688 12804 13952 12832
rect 13688 12792 13694 12804
rect 11790 12724 11796 12776
rect 11848 12764 11854 12776
rect 13924 12773 13952 12804
rect 13817 12767 13875 12773
rect 13817 12764 13829 12767
rect 11848 12736 13829 12764
rect 11848 12724 11854 12736
rect 13817 12733 13829 12736
rect 13863 12733 13875 12767
rect 13817 12727 13875 12733
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12733 13967 12767
rect 14826 12764 14832 12776
rect 14787 12736 14832 12764
rect 13909 12727 13967 12733
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 12710 12656 12716 12708
rect 12768 12696 12774 12708
rect 12805 12699 12863 12705
rect 12805 12696 12817 12699
rect 12768 12668 12817 12696
rect 12768 12656 12774 12668
rect 12805 12665 12817 12668
rect 12851 12696 12863 12699
rect 13170 12696 13176 12708
rect 12851 12668 13176 12696
rect 12851 12665 12863 12668
rect 12805 12659 12863 12665
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 14185 12699 14243 12705
rect 14185 12665 14197 12699
rect 14231 12696 14243 12699
rect 15746 12696 15752 12708
rect 14231 12668 15752 12696
rect 14231 12665 14243 12668
rect 14185 12659 14243 12665
rect 15746 12656 15752 12668
rect 15804 12656 15810 12708
rect 10744 12600 11192 12628
rect 12437 12631 12495 12637
rect 10744 12588 10750 12600
rect 12437 12597 12449 12631
rect 12483 12628 12495 12631
rect 12618 12628 12624 12640
rect 12483 12600 12624 12628
rect 12483 12597 12495 12600
rect 12437 12591 12495 12597
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 14274 12628 14280 12640
rect 12943 12600 14280 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 14274 12588 14280 12600
rect 14332 12588 14338 12640
rect 15010 12628 15016 12640
rect 14971 12600 15016 12628
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 1104 12538 15824 12560
rect 1104 12486 5912 12538
rect 5964 12486 5976 12538
rect 6028 12486 6040 12538
rect 6092 12486 6104 12538
rect 6156 12486 10843 12538
rect 10895 12486 10907 12538
rect 10959 12486 10971 12538
rect 11023 12486 11035 12538
rect 11087 12486 15824 12538
rect 1104 12464 15824 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3142 12424 3148 12436
rect 2832 12396 2877 12424
rect 3103 12396 3148 12424
rect 2832 12384 2838 12396
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 3237 12427 3295 12433
rect 3237 12393 3249 12427
rect 3283 12424 3295 12427
rect 3283 12396 5948 12424
rect 3283 12393 3295 12396
rect 3237 12387 3295 12393
rect 2041 12359 2099 12365
rect 2041 12325 2053 12359
rect 2087 12356 2099 12359
rect 5534 12356 5540 12368
rect 2087 12328 5540 12356
rect 2087 12325 2099 12328
rect 2041 12319 2099 12325
rect 5534 12316 5540 12328
rect 5592 12316 5598 12368
rect 5626 12316 5632 12368
rect 5684 12356 5690 12368
rect 5782 12359 5840 12365
rect 5782 12356 5794 12359
rect 5684 12328 5794 12356
rect 5684 12316 5690 12328
rect 5782 12325 5794 12328
rect 5828 12325 5840 12359
rect 5920 12356 5948 12396
rect 6362 12384 6368 12436
rect 6420 12424 6426 12436
rect 8757 12427 8815 12433
rect 8757 12424 8769 12427
rect 6420 12396 8769 12424
rect 6420 12384 6426 12396
rect 8757 12393 8769 12396
rect 8803 12393 8815 12427
rect 8757 12387 8815 12393
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 9122 12424 9128 12436
rect 8904 12396 9128 12424
rect 8904 12384 8910 12396
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 9217 12427 9275 12433
rect 9217 12393 9229 12427
rect 9263 12424 9275 12427
rect 9306 12424 9312 12436
rect 9263 12396 9312 12424
rect 9263 12393 9275 12396
rect 9217 12387 9275 12393
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 9582 12384 9588 12436
rect 9640 12424 9646 12436
rect 11514 12424 11520 12436
rect 9640 12396 11520 12424
rect 9640 12384 9646 12396
rect 11514 12384 11520 12396
rect 11572 12424 11578 12436
rect 12342 12424 12348 12436
rect 11572 12396 12348 12424
rect 11572 12384 11578 12396
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 12526 12424 12532 12436
rect 12487 12396 12532 12424
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 7374 12356 7380 12368
rect 5920 12328 7380 12356
rect 5782 12319 5840 12325
rect 7374 12316 7380 12328
rect 7432 12316 7438 12368
rect 7650 12365 7656 12368
rect 7644 12356 7656 12365
rect 7611 12328 7656 12356
rect 7644 12319 7656 12328
rect 7650 12316 7656 12319
rect 7708 12316 7714 12368
rect 9766 12356 9772 12368
rect 7852 12328 9772 12356
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 4706 12288 4712 12300
rect 1995 12260 3280 12288
rect 4667 12260 4712 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 3252 12232 3280 12260
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 4801 12291 4859 12297
rect 4801 12257 4813 12291
rect 4847 12288 4859 12291
rect 6362 12288 6368 12300
rect 4847 12260 6368 12288
rect 4847 12257 4859 12260
rect 4801 12251 4859 12257
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 7852 12288 7880 12328
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 10045 12359 10103 12365
rect 10045 12325 10057 12359
rect 10091 12356 10103 12359
rect 10870 12356 10876 12368
rect 10091 12328 10876 12356
rect 10091 12325 10103 12328
rect 10045 12319 10103 12325
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 11054 12316 11060 12368
rect 11112 12356 11118 12368
rect 11112 12328 13584 12356
rect 11112 12316 11118 12328
rect 7248 12260 7880 12288
rect 7248 12248 7254 12260
rect 7926 12248 7932 12300
rect 7984 12288 7990 12300
rect 8570 12288 8576 12300
rect 7984 12260 8576 12288
rect 7984 12248 7990 12260
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 9398 12288 9404 12300
rect 9359 12260 9404 12288
rect 9398 12248 9404 12260
rect 9456 12248 9462 12300
rect 11241 12291 11299 12297
rect 9876 12260 10364 12288
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 2240 12152 2268 12183
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12220 3479 12223
rect 4154 12220 4160 12232
rect 3467 12192 4160 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 4154 12180 4160 12192
rect 4212 12180 4218 12232
rect 4890 12220 4896 12232
rect 4851 12192 4896 12220
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 5074 12152 5080 12164
rect 2240 12124 5080 12152
rect 5074 12112 5080 12124
rect 5132 12112 5138 12164
rect 1581 12087 1639 12093
rect 1581 12053 1593 12087
rect 1627 12084 1639 12087
rect 2866 12084 2872 12096
rect 1627 12056 2872 12084
rect 1627 12053 1639 12056
rect 1581 12047 1639 12053
rect 2866 12044 2872 12056
rect 2924 12044 2930 12096
rect 4338 12084 4344 12096
rect 4299 12056 4344 12084
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 5166 12084 5172 12096
rect 4764 12056 5172 12084
rect 4764 12044 4770 12056
rect 5166 12044 5172 12056
rect 5224 12044 5230 12096
rect 5552 12084 5580 12183
rect 6546 12180 6552 12232
rect 6604 12220 6610 12232
rect 6730 12220 6736 12232
rect 6604 12192 6736 12220
rect 6604 12180 6610 12192
rect 6730 12180 6736 12192
rect 6788 12180 6794 12232
rect 7377 12223 7435 12229
rect 7377 12220 7389 12223
rect 7024 12192 7389 12220
rect 6914 12152 6920 12164
rect 6875 12124 6920 12152
rect 6914 12112 6920 12124
rect 6972 12112 6978 12164
rect 6638 12084 6644 12096
rect 5552 12056 6644 12084
rect 6638 12044 6644 12056
rect 6696 12084 6702 12096
rect 6822 12084 6828 12096
rect 6696 12056 6828 12084
rect 6696 12044 6702 12056
rect 6822 12044 6828 12056
rect 6880 12084 6886 12096
rect 7024 12084 7052 12192
rect 7377 12189 7389 12192
rect 7423 12189 7435 12223
rect 7377 12183 7435 12189
rect 9490 12180 9496 12232
rect 9548 12220 9554 12232
rect 9876 12220 9904 12260
rect 9548 12192 9904 12220
rect 9548 12180 9554 12192
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10336 12229 10364 12260
rect 11241 12257 11253 12291
rect 11287 12288 11299 12291
rect 11698 12288 11704 12300
rect 11287 12260 11704 12288
rect 11287 12257 11299 12260
rect 11241 12251 11299 12257
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 11882 12248 11888 12300
rect 11940 12288 11946 12300
rect 13556 12297 13584 12328
rect 12437 12291 12495 12297
rect 12437 12288 12449 12291
rect 11940 12260 12449 12288
rect 11940 12248 11946 12260
rect 12437 12257 12449 12260
rect 12483 12257 12495 12291
rect 13449 12291 13507 12297
rect 13449 12288 13461 12291
rect 12437 12251 12495 12257
rect 12544 12260 13461 12288
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 10008 12192 10149 12220
rect 10008 12180 10014 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 8662 12112 8668 12164
rect 8720 12152 8726 12164
rect 9858 12152 9864 12164
rect 8720 12124 9864 12152
rect 8720 12112 8726 12124
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 6880 12056 7052 12084
rect 6880 12044 6886 12056
rect 9122 12044 9128 12096
rect 9180 12084 9186 12096
rect 9677 12087 9735 12093
rect 9677 12084 9689 12087
rect 9180 12056 9689 12084
rect 9180 12044 9186 12056
rect 9677 12053 9689 12056
rect 9723 12053 9735 12087
rect 9677 12047 9735 12053
rect 9766 12044 9772 12096
rect 9824 12084 9830 12096
rect 10226 12084 10232 12096
rect 9824 12056 10232 12084
rect 9824 12044 9830 12056
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 10336 12084 10364 12183
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 10468 12192 10916 12220
rect 10468 12180 10474 12192
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 10778 12152 10784 12164
rect 10560 12124 10784 12152
rect 10560 12112 10566 12124
rect 10778 12112 10784 12124
rect 10836 12112 10842 12164
rect 10888 12161 10916 12192
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 11020 12192 11345 12220
rect 11020 12180 11026 12192
rect 11333 12189 11345 12192
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 11425 12223 11483 12229
rect 11425 12189 11437 12223
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 10873 12155 10931 12161
rect 10873 12121 10885 12155
rect 10919 12121 10931 12155
rect 11440 12152 11468 12183
rect 11514 12180 11520 12232
rect 11572 12220 11578 12232
rect 12544 12220 12572 12260
rect 13449 12257 13461 12260
rect 13495 12257 13507 12291
rect 13449 12251 13507 12257
rect 13541 12291 13599 12297
rect 13541 12257 13553 12291
rect 13587 12288 13599 12291
rect 14461 12291 14519 12297
rect 14461 12288 14473 12291
rect 13587 12260 14473 12288
rect 13587 12257 13599 12260
rect 13541 12251 13599 12257
rect 14461 12257 14473 12260
rect 14507 12257 14519 12291
rect 14461 12251 14519 12257
rect 11572 12192 12572 12220
rect 12621 12223 12679 12229
rect 11572 12180 11578 12192
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 13817 12223 13875 12229
rect 13817 12189 13829 12223
rect 13863 12220 13875 12223
rect 15378 12220 15384 12232
rect 13863 12192 15384 12220
rect 13863 12189 13875 12192
rect 13817 12183 13875 12189
rect 10873 12115 10931 12121
rect 11348 12124 11468 12152
rect 11348 12084 11376 12124
rect 11606 12112 11612 12164
rect 11664 12152 11670 12164
rect 12636 12152 12664 12183
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 13078 12152 13084 12164
rect 11664 12124 12664 12152
rect 12728 12124 13084 12152
rect 11664 12112 11670 12124
rect 10336 12056 11376 12084
rect 11514 12044 11520 12096
rect 11572 12084 11578 12096
rect 12069 12087 12127 12093
rect 12069 12084 12081 12087
rect 11572 12056 12081 12084
rect 11572 12044 11578 12056
rect 12069 12053 12081 12056
rect 12115 12053 12127 12087
rect 12069 12047 12127 12053
rect 12434 12044 12440 12096
rect 12492 12084 12498 12096
rect 12728 12084 12756 12124
rect 13078 12112 13084 12124
rect 13136 12112 13142 12164
rect 12492 12056 12756 12084
rect 12492 12044 12498 12056
rect 12802 12044 12808 12096
rect 12860 12084 12866 12096
rect 13265 12087 13323 12093
rect 13265 12084 13277 12087
rect 12860 12056 13277 12084
rect 12860 12044 12866 12056
rect 13265 12053 13277 12056
rect 13311 12053 13323 12087
rect 13265 12047 13323 12053
rect 14090 12044 14096 12096
rect 14148 12084 14154 12096
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 14148 12056 14657 12084
rect 14148 12044 14154 12056
rect 14645 12053 14657 12056
rect 14691 12053 14703 12087
rect 14645 12047 14703 12053
rect 1104 11994 15824 12016
rect 1104 11942 3447 11994
rect 3499 11942 3511 11994
rect 3563 11942 3575 11994
rect 3627 11942 3639 11994
rect 3691 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 13308 11994
rect 13360 11942 13372 11994
rect 13424 11942 13436 11994
rect 13488 11942 13500 11994
rect 13552 11942 15824 11994
rect 1104 11920 15824 11942
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 2501 11883 2559 11889
rect 2501 11880 2513 11883
rect 1820 11852 2513 11880
rect 1820 11840 1826 11852
rect 2501 11849 2513 11852
rect 2547 11849 2559 11883
rect 2501 11843 2559 11849
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3142 11880 3148 11892
rect 3016 11852 3148 11880
rect 3016 11840 3022 11852
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 3326 11840 3332 11892
rect 3384 11880 3390 11892
rect 3697 11883 3755 11889
rect 3697 11880 3709 11883
rect 3384 11852 3709 11880
rect 3384 11840 3390 11852
rect 3697 11849 3709 11852
rect 3743 11849 3755 11883
rect 5626 11880 5632 11892
rect 3697 11843 3755 11849
rect 4080 11852 5632 11880
rect 3145 11747 3203 11753
rect 3145 11713 3157 11747
rect 3191 11744 3203 11747
rect 3786 11744 3792 11756
rect 3191 11716 3792 11744
rect 3191 11713 3203 11716
rect 3145 11707 3203 11713
rect 3786 11704 3792 11716
rect 3844 11744 3850 11756
rect 4080 11744 4108 11852
rect 5626 11840 5632 11852
rect 5684 11840 5690 11892
rect 6546 11840 6552 11892
rect 6604 11880 6610 11892
rect 10226 11880 10232 11892
rect 6604 11852 10232 11880
rect 6604 11840 6610 11852
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 11698 11880 11704 11892
rect 10796 11852 11704 11880
rect 4430 11812 4436 11824
rect 4172 11784 4436 11812
rect 4172 11753 4200 11784
rect 4430 11772 4436 11784
rect 4488 11772 4494 11824
rect 8570 11772 8576 11824
rect 8628 11812 8634 11824
rect 9030 11812 9036 11824
rect 8628 11784 9036 11812
rect 8628 11772 8634 11784
rect 9030 11772 9036 11784
rect 9088 11772 9094 11824
rect 10796 11812 10824 11852
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 12437 11883 12495 11889
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 12894 11880 12900 11892
rect 12483 11852 12900 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 10520 11784 10824 11812
rect 3844 11716 4108 11744
rect 4157 11747 4215 11753
rect 3844 11704 3850 11716
rect 4157 11713 4169 11747
rect 4203 11713 4215 11747
rect 4157 11707 4215 11713
rect 4338 11704 4344 11756
rect 4396 11744 4402 11756
rect 4396 11716 4441 11744
rect 4396 11704 4402 11716
rect 6822 11704 6828 11756
rect 6880 11744 6886 11756
rect 7374 11744 7380 11756
rect 6880 11716 7380 11744
rect 6880 11704 6886 11716
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8846 11744 8852 11756
rect 8536 11716 8852 11744
rect 8536 11704 8542 11716
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11676 1639 11679
rect 1670 11676 1676 11688
rect 1627 11648 1676 11676
rect 1627 11645 1639 11648
rect 1581 11639 1639 11645
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 2866 11676 2872 11688
rect 2827 11648 2872 11676
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 4890 11676 4896 11688
rect 4851 11648 4896 11676
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 8938 11676 8944 11688
rect 5592 11648 8944 11676
rect 5592 11636 5598 11648
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 9582 11676 9588 11688
rect 9543 11648 9588 11676
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 1857 11611 1915 11617
rect 1857 11577 1869 11611
rect 1903 11577 1915 11611
rect 1857 11571 1915 11577
rect 2961 11611 3019 11617
rect 2961 11577 2973 11611
rect 3007 11608 3019 11611
rect 4246 11608 4252 11620
rect 3007 11580 4252 11608
rect 3007 11577 3019 11580
rect 2961 11571 3019 11577
rect 1872 11540 1900 11571
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 5166 11617 5172 11620
rect 5160 11608 5172 11617
rect 5127 11580 5172 11608
rect 5160 11571 5172 11580
rect 5166 11568 5172 11571
rect 5224 11568 5230 11620
rect 7282 11608 7288 11620
rect 6196 11580 7288 11608
rect 3142 11540 3148 11552
rect 1872 11512 3148 11540
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 4065 11543 4123 11549
rect 4065 11509 4077 11543
rect 4111 11540 4123 11543
rect 6196 11540 6224 11580
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 7558 11568 7564 11620
rect 7616 11617 7622 11620
rect 7616 11611 7680 11617
rect 7616 11577 7634 11611
rect 7668 11608 7680 11611
rect 9490 11608 9496 11620
rect 7668 11580 9496 11608
rect 7668 11577 7680 11580
rect 7616 11571 7680 11577
rect 7616 11568 7622 11571
rect 9490 11568 9496 11580
rect 9548 11608 9554 11620
rect 9784 11608 9812 11707
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10520 11744 10548 11784
rect 10870 11772 10876 11824
rect 10928 11812 10934 11824
rect 10928 11784 11192 11812
rect 10928 11772 10934 11784
rect 10100 11716 10548 11744
rect 10100 11704 10106 11716
rect 10594 11704 10600 11756
rect 10652 11704 10658 11756
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 9548 11580 9812 11608
rect 10612 11608 10640 11704
rect 10980 11620 11008 11707
rect 10873 11611 10931 11617
rect 10873 11608 10885 11611
rect 10612 11580 10885 11608
rect 9548 11568 9554 11580
rect 10873 11577 10885 11580
rect 10919 11577 10931 11611
rect 10873 11571 10931 11577
rect 10962 11568 10968 11620
rect 11020 11568 11026 11620
rect 11164 11608 11192 11784
rect 11330 11772 11336 11824
rect 11388 11812 11394 11824
rect 11514 11812 11520 11824
rect 11388 11784 11520 11812
rect 11388 11772 11394 11784
rect 11514 11772 11520 11784
rect 11572 11772 11578 11824
rect 12986 11744 12992 11756
rect 12947 11716 12992 11744
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 13909 11747 13967 11753
rect 13909 11713 13921 11747
rect 13955 11744 13967 11747
rect 15102 11744 15108 11756
rect 13955 11716 15108 11744
rect 13955 11713 13967 11716
rect 13909 11707 13967 11713
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 11238 11636 11244 11688
rect 11296 11676 11302 11688
rect 11514 11676 11520 11688
rect 11296 11648 11520 11676
rect 11296 11636 11302 11648
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11676 11667 11679
rect 12526 11676 12532 11688
rect 11655 11648 12532 11676
rect 11655 11645 11667 11648
rect 11609 11639 11667 11645
rect 12526 11636 12532 11648
rect 12584 11636 12590 11688
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11676 12955 11679
rect 13262 11676 13268 11688
rect 12943 11648 13268 11676
rect 12943 11645 12955 11648
rect 12897 11639 12955 11645
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 13633 11679 13691 11685
rect 13633 11645 13645 11679
rect 13679 11676 13691 11679
rect 13722 11676 13728 11688
rect 13679 11648 13728 11676
rect 13679 11645 13691 11648
rect 13633 11639 13691 11645
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 13814 11636 13820 11688
rect 13872 11676 13878 11688
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 13872 11648 14565 11676
rect 13872 11636 13878 11648
rect 14553 11645 14565 11648
rect 14599 11645 14611 11679
rect 14553 11639 14611 11645
rect 13906 11608 13912 11620
rect 11164 11580 13912 11608
rect 13906 11568 13912 11580
rect 13964 11568 13970 11620
rect 14829 11611 14887 11617
rect 14829 11577 14841 11611
rect 14875 11608 14887 11611
rect 16390 11608 16396 11620
rect 14875 11580 16396 11608
rect 14875 11577 14887 11580
rect 14829 11571 14887 11577
rect 16390 11568 16396 11580
rect 16448 11568 16454 11620
rect 4111 11512 6224 11540
rect 6273 11543 6331 11549
rect 4111 11509 4123 11512
rect 4065 11503 4123 11509
rect 6273 11509 6285 11543
rect 6319 11540 6331 11543
rect 6914 11540 6920 11552
rect 6319 11512 6920 11540
rect 6319 11509 6331 11512
rect 6273 11503 6331 11509
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 8757 11543 8815 11549
rect 8757 11509 8769 11543
rect 8803 11540 8815 11543
rect 8846 11540 8852 11552
rect 8803 11512 8852 11540
rect 8803 11509 8815 11512
rect 8757 11503 8815 11509
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 9214 11540 9220 11552
rect 9175 11512 9220 11540
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 9677 11543 9735 11549
rect 9677 11509 9689 11543
rect 9723 11540 9735 11543
rect 9766 11540 9772 11552
rect 9723 11512 9772 11540
rect 9723 11509 9735 11512
rect 9677 11503 9735 11509
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10226 11500 10232 11552
rect 10284 11540 10290 11552
rect 10413 11543 10471 11549
rect 10413 11540 10425 11543
rect 10284 11512 10425 11540
rect 10284 11500 10290 11512
rect 10413 11509 10425 11512
rect 10459 11509 10471 11543
rect 10413 11503 10471 11509
rect 10502 11500 10508 11552
rect 10560 11540 10566 11552
rect 10781 11543 10839 11549
rect 10781 11540 10793 11543
rect 10560 11512 10793 11540
rect 10560 11500 10566 11512
rect 10781 11509 10793 11512
rect 10827 11509 10839 11543
rect 10781 11503 10839 11509
rect 11238 11500 11244 11552
rect 11296 11540 11302 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11296 11512 11805 11540
rect 11296 11500 11302 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 12710 11500 12716 11552
rect 12768 11540 12774 11552
rect 12805 11543 12863 11549
rect 12805 11540 12817 11543
rect 12768 11512 12817 11540
rect 12768 11500 12774 11512
rect 12805 11509 12817 11512
rect 12851 11509 12863 11543
rect 12805 11503 12863 11509
rect 1104 11450 15824 11472
rect 1104 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 6104 11450
rect 6156 11398 10843 11450
rect 10895 11398 10907 11450
rect 10959 11398 10971 11450
rect 11023 11398 11035 11450
rect 11087 11398 15824 11450
rect 1104 11376 15824 11398
rect 1394 11296 1400 11348
rect 1452 11296 1458 11348
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 4617 11339 4675 11345
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 5350 11336 5356 11348
rect 4663 11308 5356 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 7834 11336 7840 11348
rect 5500 11308 7840 11336
rect 5500 11296 5506 11308
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 9490 11336 9496 11348
rect 8260 11308 9496 11336
rect 8260 11296 8266 11308
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 9677 11339 9735 11345
rect 9677 11305 9689 11339
rect 9723 11336 9735 11339
rect 9950 11336 9956 11348
rect 9723 11308 9956 11336
rect 9723 11305 9735 11308
rect 9677 11299 9735 11305
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10137 11339 10195 11345
rect 10137 11305 10149 11339
rect 10183 11336 10195 11339
rect 10410 11336 10416 11348
rect 10183 11308 10416 11336
rect 10183 11305 10195 11308
rect 10137 11299 10195 11305
rect 10410 11296 10416 11308
rect 10468 11296 10474 11348
rect 10502 11296 10508 11348
rect 10560 11336 10566 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10560 11308 10885 11336
rect 10560 11296 10566 11308
rect 10873 11305 10885 11308
rect 10919 11305 10931 11339
rect 11330 11336 11336 11348
rect 11291 11308 11336 11336
rect 10873 11299 10931 11305
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 11790 11296 11796 11348
rect 11848 11336 11854 11348
rect 12437 11339 12495 11345
rect 12437 11336 12449 11339
rect 11848 11308 12449 11336
rect 11848 11296 11854 11308
rect 12437 11305 12449 11308
rect 12483 11305 12495 11339
rect 12437 11299 12495 11305
rect 13265 11339 13323 11345
rect 13265 11305 13277 11339
rect 13311 11336 13323 11339
rect 13630 11336 13636 11348
rect 13311 11308 13636 11336
rect 13311 11305 13323 11308
rect 13265 11299 13323 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 1412 11268 1440 11296
rect 1412 11240 1624 11268
rect 1596 11212 1624 11240
rect 4430 11228 4436 11280
rect 4488 11268 4494 11280
rect 4488 11240 8964 11268
rect 4488 11228 4494 11240
rect 1578 11160 1584 11212
rect 1636 11160 1642 11212
rect 1946 11200 1952 11212
rect 1907 11172 1952 11200
rect 1946 11160 1952 11172
rect 2004 11160 2010 11212
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11200 2099 11203
rect 2406 11200 2412 11212
rect 2087 11172 2412 11200
rect 2087 11169 2099 11172
rect 2041 11163 2099 11169
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 3145 11203 3203 11209
rect 3145 11169 3157 11203
rect 3191 11200 3203 11203
rect 4614 11200 4620 11212
rect 3191 11172 4620 11200
rect 3191 11169 3203 11172
rect 3145 11163 3203 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11200 5043 11203
rect 5810 11200 5816 11212
rect 5031 11172 5672 11200
rect 5771 11172 5816 11200
rect 5031 11169 5043 11172
rect 4985 11163 5043 11169
rect 1486 11092 1492 11144
rect 1544 11132 1550 11144
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 1544 11104 2145 11132
rect 1544 11092 1550 11104
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 3237 11135 3295 11141
rect 3237 11132 3249 11135
rect 2924 11104 3249 11132
rect 2924 11092 2930 11104
rect 3237 11101 3249 11104
rect 3283 11101 3295 11135
rect 3237 11095 3295 11101
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 4798 11132 4804 11144
rect 3467 11104 4804 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 4798 11092 4804 11104
rect 4856 11092 4862 11144
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5258 11132 5264 11144
rect 5171 11104 5264 11132
rect 5077 11095 5135 11101
rect 2590 11024 2596 11076
rect 2648 11064 2654 11076
rect 2777 11067 2835 11073
rect 2777 11064 2789 11067
rect 2648 11036 2789 11064
rect 2648 11024 2654 11036
rect 2777 11033 2789 11036
rect 2823 11033 2835 11067
rect 2777 11027 2835 11033
rect 4430 11024 4436 11076
rect 4488 11064 4494 11076
rect 5092 11064 5120 11095
rect 5258 11092 5264 11104
rect 5316 11132 5322 11144
rect 5442 11132 5448 11144
rect 5316 11104 5448 11132
rect 5316 11092 5322 11104
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 5644 11132 5672 11172
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 5902 11160 5908 11212
rect 5960 11160 5966 11212
rect 6080 11203 6138 11209
rect 6080 11169 6092 11203
rect 6126 11200 6138 11203
rect 6914 11200 6920 11212
rect 6126 11172 6920 11200
rect 6126 11169 6138 11172
rect 6080 11163 6138 11169
rect 6914 11160 6920 11172
rect 6972 11200 6978 11212
rect 7466 11200 7472 11212
rect 6972 11172 7472 11200
rect 6972 11160 6978 11172
rect 7466 11160 7472 11172
rect 7524 11160 7530 11212
rect 7920 11203 7978 11209
rect 7920 11169 7932 11203
rect 7966 11200 7978 11203
rect 8936 11200 8964 11240
rect 9214 11228 9220 11280
rect 9272 11268 9278 11280
rect 10045 11271 10103 11277
rect 10045 11268 10057 11271
rect 9272 11240 10057 11268
rect 9272 11228 9278 11240
rect 10045 11237 10057 11240
rect 10091 11237 10103 11271
rect 10045 11231 10103 11237
rect 10244 11240 11376 11268
rect 10244 11200 10272 11240
rect 10962 11200 10968 11212
rect 7966 11172 8892 11200
rect 8936 11172 10272 11200
rect 10336 11172 10968 11200
rect 7966 11169 7978 11172
rect 7920 11163 7978 11169
rect 5920 11132 5948 11160
rect 8864 11144 8892 11172
rect 5644 11104 5948 11132
rect 7374 11092 7380 11144
rect 7432 11132 7438 11144
rect 7653 11135 7711 11141
rect 7653 11132 7665 11135
rect 7432 11104 7665 11132
rect 7432 11092 7438 11104
rect 7653 11101 7665 11104
rect 7699 11101 7711 11135
rect 7653 11095 7711 11101
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 9214 11132 9220 11144
rect 8904 11104 9220 11132
rect 8904 11092 8910 11104
rect 9214 11092 9220 11104
rect 9272 11132 9278 11144
rect 10336 11141 10364 11172
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 11054 11160 11060 11212
rect 11112 11200 11118 11212
rect 11241 11203 11299 11209
rect 11241 11200 11253 11203
rect 11112 11172 11253 11200
rect 11112 11160 11118 11172
rect 11241 11169 11253 11172
rect 11287 11169 11299 11203
rect 11348 11200 11376 11240
rect 11698 11228 11704 11280
rect 11756 11268 11762 11280
rect 12529 11271 12587 11277
rect 12529 11268 12541 11271
rect 11756 11240 12541 11268
rect 11756 11228 11762 11240
rect 12529 11237 12541 11240
rect 12575 11237 12587 11271
rect 12529 11231 12587 11237
rect 12618 11228 12624 11280
rect 12676 11228 12682 11280
rect 12710 11228 12716 11280
rect 12768 11268 12774 11280
rect 13170 11268 13176 11280
rect 12768 11240 13176 11268
rect 12768 11228 12774 11240
rect 13170 11228 13176 11240
rect 13228 11228 13234 11280
rect 13722 11228 13728 11280
rect 13780 11228 13786 11280
rect 12636 11200 12664 11228
rect 11348 11172 12664 11200
rect 11241 11163 11299 11169
rect 13078 11160 13084 11212
rect 13136 11200 13142 11212
rect 13633 11203 13691 11209
rect 13633 11200 13645 11203
rect 13136 11172 13645 11200
rect 13136 11160 13142 11172
rect 13633 11169 13645 11172
rect 13679 11169 13691 11203
rect 13740 11200 13768 11228
rect 14461 11203 14519 11209
rect 14461 11200 14473 11203
rect 13740 11172 14473 11200
rect 13633 11163 13691 11169
rect 14461 11169 14473 11172
rect 14507 11169 14519 11203
rect 14461 11163 14519 11169
rect 10321 11135 10379 11141
rect 10321 11132 10333 11135
rect 9272 11104 10333 11132
rect 9272 11092 9278 11104
rect 10321 11101 10333 11104
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 10594 11092 10600 11144
rect 10652 11132 10658 11144
rect 11425 11135 11483 11141
rect 11425 11132 11437 11135
rect 10652 11104 11437 11132
rect 10652 11092 10658 11104
rect 11425 11101 11437 11104
rect 11471 11101 11483 11135
rect 11425 11095 11483 11101
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 12621 11135 12679 11141
rect 12621 11132 12633 11135
rect 11848 11104 12633 11132
rect 11848 11092 11854 11104
rect 12621 11101 12633 11104
rect 12667 11101 12679 11135
rect 13722 11132 13728 11144
rect 13683 11104 13728 11132
rect 12621 11095 12679 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13817 11135 13875 11141
rect 13817 11101 13829 11135
rect 13863 11101 13875 11135
rect 13817 11095 13875 11101
rect 5810 11064 5816 11076
rect 4488 11036 5816 11064
rect 4488 11024 4494 11036
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 9033 11067 9091 11073
rect 9033 11033 9045 11067
rect 9079 11064 9091 11067
rect 9306 11064 9312 11076
rect 9079 11036 9312 11064
rect 9079 11033 9091 11036
rect 9033 11027 9091 11033
rect 9306 11024 9312 11036
rect 9364 11064 9370 11076
rect 10612 11064 10640 11092
rect 9364 11036 10640 11064
rect 9364 11024 9370 11036
rect 10962 11024 10968 11076
rect 11020 11064 11026 11076
rect 11606 11064 11612 11076
rect 11020 11036 11612 11064
rect 11020 11024 11026 11036
rect 11606 11024 11612 11036
rect 11664 11024 11670 11076
rect 12069 11067 12127 11073
rect 12069 11033 12081 11067
rect 12115 11064 12127 11067
rect 12894 11064 12900 11076
rect 12115 11036 12900 11064
rect 12115 11033 12127 11036
rect 12069 11027 12127 11033
rect 12894 11024 12900 11036
rect 12952 11024 12958 11076
rect 13538 11024 13544 11076
rect 13596 11064 13602 11076
rect 13832 11064 13860 11095
rect 13596 11036 13860 11064
rect 13596 11024 13602 11036
rect 14366 11024 14372 11076
rect 14424 11064 14430 11076
rect 14645 11067 14703 11073
rect 14645 11064 14657 11067
rect 14424 11036 14657 11064
rect 14424 11024 14430 11036
rect 14645 11033 14657 11036
rect 14691 11033 14703 11067
rect 14645 11027 14703 11033
rect 2682 10956 2688 11008
rect 2740 10996 2746 11008
rect 7006 10996 7012 11008
rect 2740 10968 7012 10996
rect 2740 10956 2746 10968
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 7190 10996 7196 11008
rect 7151 10968 7196 10996
rect 7190 10956 7196 10968
rect 7248 10956 7254 11008
rect 7282 10956 7288 11008
rect 7340 10996 7346 11008
rect 11698 10996 11704 11008
rect 7340 10968 11704 10996
rect 7340 10956 7346 10968
rect 11698 10956 11704 10968
rect 11756 10956 11762 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 12618 10996 12624 11008
rect 12492 10968 12624 10996
rect 12492 10956 12498 10968
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 1104 10906 15824 10928
rect 1104 10854 3447 10906
rect 3499 10854 3511 10906
rect 3563 10854 3575 10906
rect 3627 10854 3639 10906
rect 3691 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 13308 10906
rect 13360 10854 13372 10906
rect 13424 10854 13436 10906
rect 13488 10854 13500 10906
rect 13552 10854 15824 10906
rect 1104 10832 15824 10854
rect 3234 10752 3240 10804
rect 3292 10792 3298 10804
rect 3697 10795 3755 10801
rect 3697 10792 3709 10795
rect 3292 10764 3709 10792
rect 3292 10752 3298 10764
rect 3697 10761 3709 10764
rect 3743 10761 3755 10795
rect 5166 10792 5172 10804
rect 3697 10755 3755 10761
rect 4172 10764 5172 10792
rect 2498 10684 2504 10736
rect 2556 10724 2562 10736
rect 3050 10724 3056 10736
rect 2556 10696 3056 10724
rect 2556 10684 2562 10696
rect 3050 10684 3056 10696
rect 3108 10684 3114 10736
rect 2130 10616 2136 10668
rect 2188 10656 2194 10668
rect 2961 10659 3019 10665
rect 2961 10656 2973 10659
rect 2188 10628 2973 10656
rect 2188 10616 2194 10628
rect 2961 10625 2973 10628
rect 3007 10625 3019 10659
rect 2961 10619 3019 10625
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10656 3203 10659
rect 4172 10656 4200 10764
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 6273 10795 6331 10801
rect 6273 10792 6285 10795
rect 5684 10764 6285 10792
rect 5684 10752 5690 10764
rect 6273 10761 6285 10764
rect 6319 10761 6331 10795
rect 6273 10755 6331 10761
rect 6454 10752 6460 10804
rect 6512 10792 6518 10804
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 6512 10764 6837 10792
rect 6512 10752 6518 10764
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 6825 10755 6883 10761
rect 7282 10752 7288 10804
rect 7340 10752 7346 10804
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 8021 10795 8079 10801
rect 8021 10792 8033 10795
rect 7616 10764 8033 10792
rect 7616 10752 7622 10764
rect 8021 10761 8033 10764
rect 8067 10792 8079 10795
rect 9398 10792 9404 10804
rect 8067 10764 9404 10792
rect 8067 10761 8079 10764
rect 8021 10755 8079 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 10321 10795 10379 10801
rect 10321 10761 10333 10795
rect 10367 10792 10379 10795
rect 11054 10792 11060 10804
rect 10367 10764 11060 10792
rect 10367 10761 10379 10764
rect 10321 10755 10379 10761
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 15194 10792 15200 10804
rect 11532 10764 15200 10792
rect 3191 10628 4200 10656
rect 4341 10659 4399 10665
rect 3191 10625 3203 10628
rect 3145 10619 3203 10625
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4798 10656 4804 10668
rect 4387 10628 4804 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4798 10616 4804 10628
rect 4856 10616 4862 10668
rect 7300 10656 7328 10752
rect 11532 10724 11560 10764
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 11698 10724 11704 10736
rect 9508 10696 11560 10724
rect 11659 10696 11704 10724
rect 7466 10656 7472 10668
rect 6380 10628 7328 10656
rect 7427 10628 7472 10656
rect 1581 10591 1639 10597
rect 1581 10557 1593 10591
rect 1627 10588 1639 10591
rect 4065 10591 4123 10597
rect 1627 10560 2544 10588
rect 1627 10557 1639 10560
rect 1581 10551 1639 10557
rect 1854 10520 1860 10532
rect 1815 10492 1860 10520
rect 1854 10480 1860 10492
rect 1912 10480 1918 10532
rect 2516 10461 2544 10560
rect 4065 10557 4077 10591
rect 4111 10588 4123 10591
rect 4890 10588 4896 10600
rect 4111 10560 4752 10588
rect 4851 10560 4896 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 2590 10480 2596 10532
rect 2648 10520 2654 10532
rect 4614 10520 4620 10532
rect 2648 10492 4620 10520
rect 2648 10480 2654 10492
rect 4614 10480 4620 10492
rect 4672 10480 4678 10532
rect 4724 10520 4752 10560
rect 4890 10548 4896 10560
rect 4948 10548 4954 10600
rect 5534 10588 5540 10600
rect 5000 10560 5540 10588
rect 5000 10520 5028 10560
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 4724 10492 5028 10520
rect 5074 10480 5080 10532
rect 5132 10529 5138 10532
rect 5132 10523 5196 10529
rect 5132 10489 5150 10523
rect 5184 10489 5196 10523
rect 5132 10483 5196 10489
rect 5132 10480 5138 10483
rect 5442 10480 5448 10532
rect 5500 10520 5506 10532
rect 6380 10520 6408 10628
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 8481 10659 8539 10665
rect 8481 10656 8493 10659
rect 7567 10628 8493 10656
rect 7006 10548 7012 10600
rect 7064 10588 7070 10600
rect 7285 10591 7343 10597
rect 7285 10588 7297 10591
rect 7064 10560 7297 10588
rect 7064 10548 7070 10560
rect 7285 10557 7297 10560
rect 7331 10557 7343 10591
rect 7285 10551 7343 10557
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 7567 10588 7595 10628
rect 8481 10625 8493 10628
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 8202 10588 8208 10600
rect 7432 10560 7595 10588
rect 8163 10560 8208 10588
rect 7432 10548 7438 10560
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 9508 10588 9536 10696
rect 10778 10656 10784 10668
rect 10704 10628 10784 10656
rect 10704 10597 10732 10628
rect 10778 10616 10784 10628
rect 10836 10616 10842 10668
rect 10962 10656 10968 10668
rect 10923 10628 10968 10656
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 11532 10597 11560 10696
rect 11698 10684 11704 10696
rect 11756 10684 11762 10736
rect 12253 10727 12311 10733
rect 12253 10693 12265 10727
rect 12299 10724 12311 10727
rect 12299 10696 13584 10724
rect 12299 10693 12311 10696
rect 12253 10687 12311 10693
rect 11606 10616 11612 10668
rect 11664 10656 11670 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 11664 10628 13001 10656
rect 11664 10616 11670 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13078 10616 13084 10668
rect 13136 10616 13142 10668
rect 8680 10560 9536 10588
rect 10689 10591 10747 10597
rect 8680 10520 8708 10560
rect 10689 10557 10701 10591
rect 10735 10557 10747 10591
rect 10689 10551 10747 10557
rect 11517 10591 11575 10597
rect 11517 10557 11529 10591
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 11698 10548 11704 10600
rect 11756 10588 11762 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 11756 10560 12817 10588
rect 11756 10548 11762 10560
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 13096 10588 13124 10616
rect 13096 10560 13492 10588
rect 12805 10551 12863 10557
rect 5500 10492 6408 10520
rect 7024 10492 8708 10520
rect 8748 10523 8806 10529
rect 5500 10480 5506 10492
rect 2501 10455 2559 10461
rect 2501 10421 2513 10455
rect 2547 10421 2559 10455
rect 2501 10415 2559 10421
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 2869 10455 2927 10461
rect 2869 10452 2881 10455
rect 2832 10424 2881 10452
rect 2832 10412 2838 10424
rect 2869 10421 2881 10424
rect 2915 10421 2927 10455
rect 2869 10415 2927 10421
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10452 4215 10455
rect 7024 10452 7052 10492
rect 8748 10489 8760 10523
rect 8794 10520 8806 10523
rect 9306 10520 9312 10532
rect 8794 10492 9312 10520
rect 8794 10489 8806 10492
rect 8748 10483 8806 10489
rect 9306 10480 9312 10492
rect 9364 10480 9370 10532
rect 12253 10523 12311 10529
rect 12253 10520 12265 10523
rect 11624 10492 12265 10520
rect 4203 10424 7052 10452
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7193 10455 7251 10461
rect 7193 10452 7205 10455
rect 7156 10424 7205 10452
rect 7156 10412 7162 10424
rect 7193 10421 7205 10424
rect 7239 10452 7251 10455
rect 8846 10452 8852 10464
rect 7239 10424 8852 10452
rect 7239 10421 7251 10424
rect 7193 10415 7251 10421
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 9861 10455 9919 10461
rect 9861 10421 9873 10455
rect 9907 10452 9919 10455
rect 10410 10452 10416 10464
rect 9907 10424 10416 10452
rect 9907 10421 9919 10424
rect 9861 10415 9919 10421
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10560 10424 10793 10452
rect 10560 10412 10566 10424
rect 10781 10421 10793 10424
rect 10827 10452 10839 10455
rect 11624 10452 11652 10492
rect 12253 10489 12265 10492
rect 12299 10489 12311 10523
rect 12253 10483 12311 10489
rect 12342 10480 12348 10532
rect 12400 10520 12406 10532
rect 12897 10523 12955 10529
rect 12897 10520 12909 10523
rect 12400 10492 12909 10520
rect 12400 10480 12406 10492
rect 12897 10489 12909 10492
rect 12943 10520 12955 10523
rect 13078 10520 13084 10532
rect 12943 10492 13084 10520
rect 12943 10489 12955 10492
rect 12897 10483 12955 10489
rect 13078 10480 13084 10492
rect 13136 10480 13142 10532
rect 10827 10424 11652 10452
rect 10827 10421 10839 10424
rect 10781 10415 10839 10421
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 13464 10452 13492 10560
rect 13556 10520 13584 10696
rect 13814 10684 13820 10736
rect 13872 10724 13878 10736
rect 15013 10727 15071 10733
rect 15013 10724 15025 10727
rect 13872 10696 15025 10724
rect 13872 10684 13878 10696
rect 15013 10693 15025 10696
rect 15059 10693 15071 10727
rect 15013 10687 15071 10693
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 13832 10628 14197 10656
rect 13832 10600 13860 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 13814 10548 13820 10600
rect 13872 10548 13878 10600
rect 13998 10588 14004 10600
rect 13959 10560 14004 10588
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 16758 10588 16764 10600
rect 14875 10560 16764 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 14844 10520 14872 10551
rect 16758 10548 16764 10560
rect 16816 10548 16822 10600
rect 13556 10492 14872 10520
rect 13633 10455 13691 10461
rect 13633 10452 13645 10455
rect 12492 10424 12537 10452
rect 13464 10424 13645 10452
rect 12492 10412 12498 10424
rect 13633 10421 13645 10424
rect 13679 10421 13691 10455
rect 13633 10415 13691 10421
rect 14093 10455 14151 10461
rect 14093 10421 14105 10455
rect 14139 10452 14151 10455
rect 14182 10452 14188 10464
rect 14139 10424 14188 10452
rect 14139 10421 14151 10424
rect 14093 10415 14151 10421
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 1104 10362 15824 10384
rect 1104 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 6104 10362
rect 6156 10310 10843 10362
rect 10895 10310 10907 10362
rect 10959 10310 10971 10362
rect 11023 10310 11035 10362
rect 11087 10310 15824 10362
rect 1104 10288 15824 10310
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 2832 10220 2877 10248
rect 2832 10208 2838 10220
rect 3234 10208 3240 10260
rect 3292 10248 3298 10260
rect 3970 10248 3976 10260
rect 3292 10220 3976 10248
rect 3292 10208 3298 10220
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 4246 10248 4252 10260
rect 4207 10220 4252 10248
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 4338 10208 4344 10260
rect 4396 10248 4402 10260
rect 4709 10251 4767 10257
rect 4709 10248 4721 10251
rect 4396 10220 4721 10248
rect 4396 10208 4402 10220
rect 4709 10217 4721 10220
rect 4755 10217 4767 10251
rect 4709 10211 4767 10217
rect 4890 10208 4896 10260
rect 4948 10248 4954 10260
rect 5442 10248 5448 10260
rect 4948 10220 5448 10248
rect 4948 10208 4954 10220
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 7190 10248 7196 10260
rect 5727 10220 7196 10248
rect 1949 10183 2007 10189
rect 1949 10149 1961 10183
rect 1995 10180 2007 10183
rect 4430 10180 4436 10192
rect 1995 10152 4436 10180
rect 1995 10149 2007 10152
rect 1949 10143 2007 10149
rect 4430 10140 4436 10152
rect 4488 10140 4494 10192
rect 4614 10180 4620 10192
rect 4575 10152 4620 10180
rect 4614 10140 4620 10152
rect 4672 10140 4678 10192
rect 4798 10140 4804 10192
rect 4856 10180 4862 10192
rect 5727 10189 5755 10220
rect 7190 10208 7196 10220
rect 7248 10248 7254 10260
rect 7248 10220 7788 10248
rect 7248 10208 7254 10220
rect 5712 10183 5770 10189
rect 5712 10180 5724 10183
rect 4856 10152 5724 10180
rect 4856 10140 4862 10152
rect 5712 10149 5724 10152
rect 5758 10149 5770 10183
rect 7760 10180 7788 10220
rect 8018 10208 8024 10260
rect 8076 10248 8082 10260
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 8076 10220 10885 10248
rect 8076 10208 8082 10220
rect 10873 10217 10885 10220
rect 10919 10217 10931 10251
rect 10873 10211 10931 10217
rect 11241 10251 11299 10257
rect 11241 10217 11253 10251
rect 11287 10248 11299 10251
rect 11422 10248 11428 10260
rect 11287 10220 11428 10248
rect 11287 10217 11299 10220
rect 11241 10211 11299 10217
rect 11422 10208 11428 10220
rect 11480 10248 11486 10260
rect 12066 10248 12072 10260
rect 11480 10220 12072 10248
rect 11480 10208 11486 10220
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 13265 10251 13323 10257
rect 12176 10220 13032 10248
rect 5712 10143 5770 10149
rect 5828 10152 7687 10180
rect 7760 10152 9444 10180
rect 2041 10115 2099 10121
rect 2041 10081 2053 10115
rect 2087 10112 2099 10115
rect 2774 10112 2780 10124
rect 2087 10084 2780 10112
rect 2087 10081 2099 10084
rect 2041 10075 2099 10081
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 3145 10115 3203 10121
rect 3145 10081 3157 10115
rect 3191 10081 3203 10115
rect 3145 10075 3203 10081
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 5828 10112 5856 10152
rect 3283 10084 5856 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10013 2283 10047
rect 2225 10007 2283 10013
rect 2240 9976 2268 10007
rect 3160 9976 3188 10075
rect 6822 10072 6828 10124
rect 6880 10112 6886 10124
rect 7285 10115 7343 10121
rect 7285 10112 7297 10115
rect 6880 10084 7297 10112
rect 6880 10072 6886 10084
rect 7285 10081 7297 10084
rect 7331 10112 7343 10115
rect 7374 10112 7380 10124
rect 7331 10084 7380 10112
rect 7331 10081 7343 10084
rect 7285 10075 7343 10081
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 7558 10121 7564 10124
rect 7552 10112 7564 10121
rect 7519 10084 7564 10112
rect 7552 10075 7564 10084
rect 7558 10072 7564 10075
rect 7616 10072 7622 10124
rect 7659 10112 7687 10152
rect 8018 10112 8024 10124
rect 7659 10084 8024 10112
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 9306 10112 9312 10124
rect 9267 10084 9312 10112
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 9416 10112 9444 10152
rect 9766 10140 9772 10192
rect 9824 10180 9830 10192
rect 10137 10183 10195 10189
rect 10137 10180 10149 10183
rect 9824 10152 10149 10180
rect 9824 10140 9830 10152
rect 10137 10149 10149 10152
rect 10183 10180 10195 10183
rect 10226 10180 10232 10192
rect 10183 10152 10232 10180
rect 10183 10149 10195 10152
rect 10137 10143 10195 10149
rect 10226 10140 10232 10152
rect 10284 10140 10290 10192
rect 10410 10140 10416 10192
rect 10468 10180 10474 10192
rect 10686 10180 10692 10192
rect 10468 10152 10692 10180
rect 10468 10140 10474 10152
rect 10686 10140 10692 10152
rect 10744 10180 10750 10192
rect 12176 10180 12204 10220
rect 10744 10152 12204 10180
rect 12437 10183 12495 10189
rect 10744 10140 10750 10152
rect 12437 10149 12449 10183
rect 12483 10180 12495 10183
rect 12894 10180 12900 10192
rect 12483 10152 12900 10180
rect 12483 10149 12495 10152
rect 12437 10143 12495 10149
rect 12894 10140 12900 10152
rect 12952 10140 12958 10192
rect 13004 10180 13032 10220
rect 13265 10217 13277 10251
rect 13311 10248 13323 10251
rect 13722 10248 13728 10260
rect 13311 10220 13728 10248
rect 13311 10217 13323 10220
rect 13265 10211 13323 10217
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 15562 10180 15568 10192
rect 13004 10152 15568 10180
rect 15562 10140 15568 10152
rect 15620 10140 15626 10192
rect 10045 10115 10103 10121
rect 9416 10084 9904 10112
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10044 3479 10047
rect 3878 10044 3884 10056
rect 3467 10016 3884 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10044 4951 10047
rect 5074 10044 5080 10056
rect 4939 10016 5080 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 5074 10004 5080 10016
rect 5132 10044 5138 10056
rect 5132 10016 5396 10044
rect 5132 10004 5138 10016
rect 5258 9976 5264 9988
rect 2240 9948 3096 9976
rect 3160 9948 5264 9976
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 2590 9908 2596 9920
rect 1627 9880 2596 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 3068 9908 3096 9948
rect 5258 9936 5264 9948
rect 5316 9936 5322 9988
rect 5074 9908 5080 9920
rect 3068 9880 5080 9908
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 5368 9908 5396 10016
rect 5442 10004 5448 10056
rect 5500 10044 5506 10056
rect 9876 10044 9904 10084
rect 10045 10081 10057 10115
rect 10091 10112 10103 10115
rect 11238 10112 11244 10124
rect 10091 10084 11244 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 11698 10112 11704 10124
rect 11348 10084 11704 10112
rect 10229 10047 10287 10053
rect 10229 10044 10241 10047
rect 5500 10016 5545 10044
rect 9416 10016 9812 10044
rect 9876 10016 10241 10044
rect 5500 10004 5506 10016
rect 9416 9976 9444 10016
rect 9048 9948 9444 9976
rect 6825 9911 6883 9917
rect 6825 9908 6837 9911
rect 5368 9880 6837 9908
rect 6825 9877 6837 9880
rect 6871 9877 6883 9911
rect 6825 9871 6883 9877
rect 7650 9868 7656 9920
rect 7708 9908 7714 9920
rect 8665 9911 8723 9917
rect 8665 9908 8677 9911
rect 7708 9880 8677 9908
rect 7708 9868 7714 9880
rect 8665 9877 8677 9880
rect 8711 9908 8723 9911
rect 9048 9908 9076 9948
rect 9490 9936 9496 9988
rect 9548 9976 9554 9988
rect 9677 9979 9735 9985
rect 9677 9976 9689 9979
rect 9548 9948 9689 9976
rect 9548 9936 9554 9948
rect 9677 9945 9689 9948
rect 9723 9945 9735 9979
rect 9784 9976 9812 10016
rect 10229 10013 10241 10016
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11348 10053 11376 10084
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 12636 10084 13645 10112
rect 12636 10056 12664 10084
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 13725 10115 13783 10121
rect 13725 10081 13737 10115
rect 13771 10112 13783 10115
rect 13906 10112 13912 10124
rect 13771 10084 13912 10112
rect 13771 10081 13783 10084
rect 13725 10075 13783 10081
rect 13906 10072 13912 10084
rect 13964 10072 13970 10124
rect 14461 10115 14519 10121
rect 14461 10081 14473 10115
rect 14507 10112 14519 10115
rect 14550 10112 14556 10124
rect 14507 10084 14556 10112
rect 14507 10081 14519 10084
rect 14461 10075 14519 10081
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 14642 10072 14648 10124
rect 14700 10112 14706 10124
rect 14918 10112 14924 10124
rect 14700 10084 14924 10112
rect 14700 10072 14706 10084
rect 14918 10072 14924 10084
rect 14976 10072 14982 10124
rect 11333 10047 11391 10053
rect 11333 10044 11345 10047
rect 11112 10016 11345 10044
rect 11112 10004 11118 10016
rect 11333 10013 11345 10016
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10044 11575 10047
rect 11606 10044 11612 10056
rect 11563 10016 11612 10044
rect 11563 10013 11575 10016
rect 11517 10007 11575 10013
rect 10410 9976 10416 9988
rect 9784 9948 10416 9976
rect 9677 9939 9735 9945
rect 10410 9936 10416 9948
rect 10468 9976 10474 9988
rect 11532 9976 11560 10007
rect 11606 10004 11612 10016
rect 11664 10004 11670 10056
rect 12066 10004 12072 10056
rect 12124 10044 12130 10056
rect 12529 10047 12587 10053
rect 12529 10044 12541 10047
rect 12124 10016 12541 10044
rect 12124 10004 12130 10016
rect 12529 10013 12541 10016
rect 12575 10013 12587 10047
rect 12529 10007 12587 10013
rect 12618 10004 12624 10056
rect 12676 10004 12682 10056
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10044 12771 10047
rect 12894 10044 12900 10056
rect 12759 10016 12900 10044
rect 12759 10013 12771 10016
rect 12713 10007 12771 10013
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 13814 10044 13820 10056
rect 13775 10016 13820 10044
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 13924 10044 13952 10072
rect 15470 10044 15476 10056
rect 13924 10016 15476 10044
rect 15470 10004 15476 10016
rect 15528 10004 15534 10056
rect 14642 9976 14648 9988
rect 10468 9948 11560 9976
rect 11624 9948 12204 9976
rect 14603 9948 14648 9976
rect 10468 9936 10474 9948
rect 8711 9880 9076 9908
rect 9125 9911 9183 9917
rect 8711 9877 8723 9880
rect 8665 9871 8723 9877
rect 9125 9877 9137 9911
rect 9171 9908 9183 9911
rect 9398 9908 9404 9920
rect 9171 9880 9404 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9398 9868 9404 9880
rect 9456 9908 9462 9920
rect 11624 9908 11652 9948
rect 9456 9880 11652 9908
rect 9456 9868 9462 9880
rect 11698 9868 11704 9920
rect 11756 9908 11762 9920
rect 12069 9911 12127 9917
rect 12069 9908 12081 9911
rect 11756 9880 12081 9908
rect 11756 9868 11762 9880
rect 12069 9877 12081 9880
rect 12115 9877 12127 9911
rect 12176 9908 12204 9948
rect 14642 9936 14648 9948
rect 14700 9936 14706 9988
rect 15286 9908 15292 9920
rect 12176 9880 15292 9908
rect 12069 9871 12127 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 1104 9818 15824 9840
rect 1104 9766 3447 9818
rect 3499 9766 3511 9818
rect 3563 9766 3575 9818
rect 3627 9766 3639 9818
rect 3691 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 13308 9818
rect 13360 9766 13372 9818
rect 13424 9766 13436 9818
rect 13488 9766 13500 9818
rect 13552 9766 15824 9818
rect 1104 9744 15824 9766
rect 4890 9704 4896 9716
rect 3804 9676 4896 9704
rect 2130 9636 2136 9648
rect 2091 9608 2136 9636
rect 2130 9596 2136 9608
rect 2188 9596 2194 9648
rect 3694 9636 3700 9648
rect 2424 9608 3700 9636
rect 2424 9568 2452 9608
rect 3694 9596 3700 9608
rect 3752 9596 3758 9648
rect 2590 9568 2596 9580
rect 1596 9540 2452 9568
rect 2551 9540 2596 9568
rect 1596 9509 1624 9540
rect 2590 9528 2596 9540
rect 2648 9528 2654 9580
rect 3804 9577 3832 9676
rect 4890 9664 4896 9676
rect 4948 9664 4954 9716
rect 5166 9704 5172 9716
rect 5127 9676 5172 9704
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 5316 9676 8800 9704
rect 5316 9664 5322 9676
rect 8772 9636 8800 9676
rect 9214 9664 9220 9716
rect 9272 9704 9278 9716
rect 9398 9704 9404 9716
rect 9272 9676 9404 9704
rect 9272 9664 9278 9676
rect 9398 9664 9404 9676
rect 9456 9664 9462 9716
rect 10226 9664 10232 9716
rect 10284 9704 10290 9716
rect 11330 9704 11336 9716
rect 10284 9676 11336 9704
rect 10284 9664 10290 9676
rect 11330 9664 11336 9676
rect 11388 9664 11394 9716
rect 11606 9664 11612 9716
rect 11664 9704 11670 9716
rect 12158 9704 12164 9716
rect 11664 9676 12164 9704
rect 11664 9664 11670 9676
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12437 9707 12495 9713
rect 12437 9673 12449 9707
rect 12483 9704 12495 9707
rect 13814 9704 13820 9716
rect 12483 9676 13820 9704
rect 12483 9673 12495 9676
rect 12437 9667 12495 9673
rect 13814 9664 13820 9676
rect 13872 9664 13878 9716
rect 13998 9664 14004 9716
rect 14056 9704 14062 9716
rect 14182 9704 14188 9716
rect 14056 9676 14188 9704
rect 14056 9664 14062 9676
rect 14182 9664 14188 9676
rect 14240 9704 14246 9716
rect 14240 9676 14872 9704
rect 14240 9664 14246 9676
rect 9861 9639 9919 9645
rect 9861 9636 9873 9639
rect 8772 9608 9873 9636
rect 9861 9605 9873 9608
rect 9907 9605 9919 9639
rect 12342 9636 12348 9648
rect 9861 9599 9919 9605
rect 10152 9608 12348 9636
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9568 2835 9571
rect 3605 9571 3663 9577
rect 2823 9540 3464 9568
rect 2823 9537 2835 9540
rect 2777 9531 2835 9537
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9469 1639 9503
rect 1581 9463 1639 9469
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9500 1915 9503
rect 2866 9500 2872 9512
rect 1903 9472 2872 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 3326 9500 3332 9512
rect 3016 9472 3332 9500
rect 3016 9460 3022 9472
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 2498 9432 2504 9444
rect 2459 9404 2504 9432
rect 2498 9392 2504 9404
rect 2556 9392 2562 9444
rect 3436 9432 3464 9540
rect 3605 9537 3617 9571
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 3620 9500 3648 9531
rect 4890 9528 4896 9580
rect 4948 9568 4954 9580
rect 5261 9571 5319 9577
rect 5261 9568 5273 9571
rect 4948 9540 5273 9568
rect 4948 9528 4954 9540
rect 5261 9537 5273 9540
rect 5307 9537 5319 9571
rect 6822 9568 6828 9580
rect 6783 9540 6828 9568
rect 5261 9531 5319 9537
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 8110 9528 8116 9580
rect 8168 9568 8174 9580
rect 9214 9568 9220 9580
rect 8168 9540 9220 9568
rect 8168 9528 8174 9540
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9568 9367 9571
rect 9398 9568 9404 9580
rect 9355 9540 9404 9568
rect 9355 9537 9367 9540
rect 9309 9531 9367 9537
rect 9398 9528 9404 9540
rect 9456 9528 9462 9580
rect 3620 9472 5672 9500
rect 3878 9432 3884 9444
rect 3436 9404 3884 9432
rect 3878 9392 3884 9404
rect 3936 9432 3942 9444
rect 5534 9441 5540 9444
rect 4056 9435 4114 9441
rect 4056 9432 4068 9435
rect 3936 9404 4068 9432
rect 3936 9392 3942 9404
rect 4056 9401 4068 9404
rect 4102 9432 4114 9435
rect 5528 9432 5540 9441
rect 4102 9404 5304 9432
rect 5495 9404 5540 9432
rect 4102 9401 4114 9404
rect 4056 9395 4114 9401
rect 2958 9364 2964 9376
rect 2919 9336 2964 9364
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3326 9364 3332 9376
rect 3287 9336 3332 9364
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 3421 9367 3479 9373
rect 3421 9333 3433 9367
rect 3467 9364 3479 9367
rect 5166 9364 5172 9376
rect 3467 9336 5172 9364
rect 3467 9333 3479 9336
rect 3421 9327 3479 9333
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5276 9364 5304 9404
rect 5528 9395 5540 9404
rect 5534 9392 5540 9395
rect 5592 9392 5598 9444
rect 5644 9432 5672 9472
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 8202 9500 8208 9512
rect 5868 9472 8208 9500
rect 5868 9460 5874 9472
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9469 9091 9503
rect 9033 9463 9091 9469
rect 6270 9432 6276 9444
rect 5644 9404 6276 9432
rect 6270 9392 6276 9404
rect 6328 9432 6334 9444
rect 7070 9435 7128 9441
rect 7070 9432 7082 9435
rect 6328 9404 7082 9432
rect 6328 9392 6334 9404
rect 7070 9401 7082 9404
rect 7116 9401 7128 9435
rect 7070 9395 7128 9401
rect 7834 9392 7840 9444
rect 7892 9432 7898 9444
rect 8294 9432 8300 9444
rect 7892 9404 8300 9432
rect 7892 9392 7898 9404
rect 8294 9392 8300 9404
rect 8352 9392 8358 9444
rect 9048 9432 9076 9463
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 10152 9500 10180 9608
rect 12342 9596 12348 9608
rect 12400 9636 12406 9648
rect 12710 9636 12716 9648
rect 12400 9608 12716 9636
rect 12400 9596 12406 9608
rect 12710 9596 12716 9608
rect 12768 9596 12774 9648
rect 12802 9596 12808 9648
rect 12860 9636 12866 9648
rect 13633 9639 13691 9645
rect 13633 9636 13645 9639
rect 12860 9608 13645 9636
rect 12860 9596 12866 9608
rect 13633 9605 13645 9608
rect 13679 9605 13691 9639
rect 13633 9599 13691 9605
rect 13722 9596 13728 9648
rect 13780 9636 13786 9648
rect 13780 9608 14228 9636
rect 13780 9596 13786 9608
rect 10410 9568 10416 9580
rect 10371 9540 10416 9568
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 10594 9528 10600 9580
rect 10652 9568 10658 9580
rect 11609 9571 11667 9577
rect 11609 9568 11621 9571
rect 10652 9540 11621 9568
rect 10652 9528 10658 9540
rect 11609 9537 11621 9540
rect 11655 9568 11667 9571
rect 12618 9568 12624 9580
rect 11655 9540 12624 9568
rect 11655 9537 11667 9540
rect 11609 9531 11667 9537
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 9180 9472 9225 9500
rect 9324 9472 10180 9500
rect 10229 9503 10287 9509
rect 9180 9460 9186 9472
rect 9324 9432 9352 9472
rect 10229 9469 10241 9503
rect 10275 9500 10287 9503
rect 11146 9500 11152 9512
rect 10275 9472 11152 9500
rect 10275 9469 10287 9472
rect 10229 9463 10287 9469
rect 11146 9460 11152 9472
rect 11204 9460 11210 9512
rect 11422 9460 11428 9512
rect 11480 9460 11486 9512
rect 11517 9503 11575 9509
rect 11517 9469 11529 9503
rect 11563 9500 11575 9503
rect 12250 9500 12256 9512
rect 11563 9472 12256 9500
rect 11563 9469 11575 9472
rect 11517 9463 11575 9469
rect 12250 9460 12256 9472
rect 12308 9500 12314 9512
rect 12710 9500 12716 9512
rect 12308 9472 12716 9500
rect 12308 9460 12314 9472
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 9048 9404 9352 9432
rect 10686 9392 10692 9444
rect 10744 9432 10750 9444
rect 11440 9432 11468 9460
rect 12802 9432 12808 9444
rect 10744 9404 11468 9432
rect 12763 9404 12808 9432
rect 10744 9392 10750 9404
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 13004 9432 13032 9531
rect 13078 9528 13084 9580
rect 13136 9568 13142 9580
rect 14200 9577 14228 9608
rect 14093 9571 14151 9577
rect 14093 9568 14105 9571
rect 13136 9540 14105 9568
rect 13136 9528 13142 9540
rect 14093 9537 14105 9540
rect 14139 9537 14151 9571
rect 14093 9531 14151 9537
rect 14185 9571 14243 9577
rect 14185 9537 14197 9571
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 14844 9509 14872 9676
rect 14001 9503 14059 9509
rect 14001 9500 14013 9503
rect 13964 9472 14013 9500
rect 13964 9460 13970 9472
rect 14001 9469 14013 9472
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 13078 9432 13084 9444
rect 13004 9404 13084 9432
rect 13078 9392 13084 9404
rect 13136 9392 13142 9444
rect 6641 9367 6699 9373
rect 6641 9364 6653 9367
rect 5276 9336 6653 9364
rect 6641 9333 6653 9336
rect 6687 9333 6699 9367
rect 6641 9327 6699 9333
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7558 9364 7564 9376
rect 6972 9336 7564 9364
rect 6972 9324 6978 9336
rect 7558 9324 7564 9336
rect 7616 9364 7622 9376
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 7616 9336 8217 9364
rect 7616 9324 7622 9336
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 8205 9327 8263 9333
rect 8665 9367 8723 9373
rect 8665 9333 8677 9367
rect 8711 9364 8723 9367
rect 9674 9364 9680 9376
rect 8711 9336 9680 9364
rect 8711 9333 8723 9336
rect 8665 9327 8723 9333
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 10318 9364 10324 9376
rect 10279 9336 10324 9364
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 11057 9367 11115 9373
rect 11057 9333 11069 9367
rect 11103 9364 11115 9367
rect 11330 9364 11336 9376
rect 11103 9336 11336 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 11425 9367 11483 9373
rect 11425 9333 11437 9367
rect 11471 9364 11483 9367
rect 11514 9364 11520 9376
rect 11471 9336 11520 9364
rect 11471 9333 11483 9336
rect 11425 9327 11483 9333
rect 11514 9324 11520 9336
rect 11572 9364 11578 9376
rect 11790 9364 11796 9376
rect 11572 9336 11796 9364
rect 11572 9324 11578 9336
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 12250 9324 12256 9376
rect 12308 9364 12314 9376
rect 12897 9367 12955 9373
rect 12897 9364 12909 9367
rect 12308 9336 12909 9364
rect 12308 9324 12314 9336
rect 12897 9333 12909 9336
rect 12943 9333 12955 9367
rect 12897 9327 12955 9333
rect 14182 9324 14188 9376
rect 14240 9364 14246 9376
rect 15013 9367 15071 9373
rect 15013 9364 15025 9367
rect 14240 9336 15025 9364
rect 14240 9324 14246 9336
rect 15013 9333 15025 9336
rect 15059 9333 15071 9367
rect 15013 9327 15071 9333
rect 1104 9274 15824 9296
rect 1104 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 6104 9274
rect 6156 9222 10843 9274
rect 10895 9222 10907 9274
rect 10959 9222 10971 9274
rect 11023 9222 11035 9274
rect 11087 9222 15824 9274
rect 1104 9200 15824 9222
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 2832 9132 2877 9160
rect 2832 9120 2838 9132
rect 3326 9120 3332 9172
rect 3384 9160 3390 9172
rect 10873 9163 10931 9169
rect 10873 9160 10885 9163
rect 3384 9132 10885 9160
rect 3384 9120 3390 9132
rect 10873 9129 10885 9132
rect 10919 9129 10931 9163
rect 11330 9160 11336 9172
rect 11291 9132 11336 9160
rect 10873 9123 10931 9129
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 13170 9120 13176 9172
rect 13228 9160 13234 9172
rect 13265 9163 13323 9169
rect 13265 9160 13277 9163
rect 13228 9132 13277 9160
rect 13228 9120 13234 9132
rect 13265 9129 13277 9132
rect 13311 9129 13323 9163
rect 14918 9160 14924 9172
rect 13265 9123 13323 9129
rect 13648 9132 14924 9160
rect 1302 9052 1308 9104
rect 1360 9092 1366 9104
rect 3237 9095 3295 9101
rect 3237 9092 3249 9095
rect 1360 9064 3249 9092
rect 1360 9052 1366 9064
rect 3237 9061 3249 9064
rect 3283 9061 3295 9095
rect 3237 9055 3295 9061
rect 5626 9052 5632 9104
rect 5684 9092 5690 9104
rect 7558 9092 7564 9104
rect 5684 9064 7564 9092
rect 5684 9052 5690 9064
rect 7558 9052 7564 9064
rect 7616 9052 7622 9104
rect 7650 9052 7656 9104
rect 7708 9092 7714 9104
rect 7834 9092 7840 9104
rect 7708 9064 7840 9092
rect 7708 9052 7714 9064
rect 7834 9052 7840 9064
rect 7892 9052 7898 9104
rect 8018 9052 8024 9104
rect 8076 9092 8082 9104
rect 8113 9095 8171 9101
rect 8113 9092 8125 9095
rect 8076 9064 8125 9092
rect 8076 9052 8082 9064
rect 8113 9061 8125 9064
rect 8159 9061 8171 9095
rect 8113 9055 8171 9061
rect 8205 9095 8263 9101
rect 8205 9061 8217 9095
rect 8251 9092 8263 9095
rect 8386 9092 8392 9104
rect 8251 9064 8392 9092
rect 8251 9061 8263 9064
rect 8205 9055 8263 9061
rect 8386 9052 8392 9064
rect 8444 9052 8450 9104
rect 8662 9092 8668 9104
rect 8588 9064 8668 9092
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 9024 2007 9027
rect 2590 9024 2596 9036
rect 1995 8996 2596 9024
rect 1995 8993 2007 8996
rect 1949 8987 2007 8993
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 8993 3203 9027
rect 4614 9024 4620 9036
rect 4527 8996 4620 9024
rect 3145 8987 3203 8993
rect 1762 8916 1768 8968
rect 1820 8956 1826 8968
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 1820 8928 2053 8956
rect 1820 8916 1826 8928
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2682 8956 2688 8968
rect 2271 8928 2688 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 3160 8888 3188 8987
rect 4614 8984 4620 8996
rect 4672 9024 4678 9036
rect 4798 9024 4804 9036
rect 4672 8996 4804 9024
rect 4672 8984 4678 8996
rect 4798 8984 4804 8996
rect 4856 8984 4862 9036
rect 5074 8984 5080 9036
rect 5132 9024 5138 9036
rect 8588 9033 8616 9064
rect 8662 9052 8668 9064
rect 8720 9052 8726 9104
rect 8846 9052 8852 9104
rect 8904 9092 8910 9104
rect 9122 9092 9128 9104
rect 8904 9064 9128 9092
rect 8904 9052 8910 9064
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 10134 9092 10140 9104
rect 10095 9064 10140 9092
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 10318 9052 10324 9104
rect 10376 9092 10382 9104
rect 13648 9092 13676 9132
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 10376 9064 13676 9092
rect 13725 9095 13783 9101
rect 10376 9052 10382 9064
rect 13725 9061 13737 9095
rect 13771 9092 13783 9095
rect 13814 9092 13820 9104
rect 13771 9064 13820 9092
rect 13771 9061 13783 9064
rect 13725 9055 13783 9061
rect 13814 9052 13820 9064
rect 13872 9052 13878 9104
rect 5905 9027 5963 9033
rect 5905 9024 5917 9027
rect 5132 8996 5917 9024
rect 5132 8984 5138 8996
rect 5905 8993 5917 8996
rect 5951 8993 5963 9027
rect 8573 9027 8631 9033
rect 5905 8987 5963 8993
rect 6564 8996 8524 9024
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 4430 8956 4436 8968
rect 3467 8928 4436 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 4522 8916 4528 8968
rect 4580 8956 4586 8968
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 4580 8928 4721 8956
rect 4580 8916 4586 8928
rect 4709 8925 4721 8928
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8956 4951 8959
rect 4982 8956 4988 8968
rect 4939 8928 4988 8956
rect 4939 8925 4951 8928
rect 4893 8919 4951 8925
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 5166 8916 5172 8968
rect 5224 8956 5230 8968
rect 6564 8956 6592 8996
rect 8294 8956 8300 8968
rect 5224 8928 6592 8956
rect 8255 8928 8300 8956
rect 5224 8916 5230 8928
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 8496 8956 8524 8996
rect 8573 8993 8585 9027
rect 8619 8993 8631 9027
rect 9398 9024 9404 9036
rect 8573 8987 8631 8993
rect 8680 8996 9404 9024
rect 8680 8956 8708 8996
rect 9398 8984 9404 8996
rect 9456 8984 9462 9036
rect 9858 8984 9864 9036
rect 9916 9024 9922 9036
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 9916 8996 10057 9024
rect 9916 8984 9922 8996
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 11238 9024 11244 9036
rect 10045 8987 10103 8993
rect 10152 8996 10548 9024
rect 11199 8996 11244 9024
rect 8496 8928 8708 8956
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8925 8815 8959
rect 8757 8919 8815 8925
rect 3326 8888 3332 8900
rect 3160 8860 3332 8888
rect 3326 8848 3332 8860
rect 3384 8888 3390 8900
rect 7466 8888 7472 8900
rect 3384 8860 7472 8888
rect 3384 8848 3390 8860
rect 7466 8848 7472 8860
rect 7524 8848 7530 8900
rect 7742 8888 7748 8900
rect 7703 8860 7748 8888
rect 7742 8848 7748 8860
rect 7800 8848 7806 8900
rect 7834 8848 7840 8900
rect 7892 8888 7898 8900
rect 8772 8888 8800 8919
rect 9214 8916 9220 8968
rect 9272 8956 9278 8968
rect 10152 8956 10180 8996
rect 9272 8928 10180 8956
rect 10321 8959 10379 8965
rect 9272 8916 9278 8928
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 10410 8956 10416 8968
rect 10367 8928 10416 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10520 8956 10548 8996
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 12434 9024 12440 9036
rect 12395 8996 12440 9024
rect 12434 8984 12440 8996
rect 12492 8984 12498 9036
rect 13170 8984 13176 9036
rect 13228 9024 13234 9036
rect 13633 9027 13691 9033
rect 13633 9024 13645 9027
rect 13228 8996 13645 9024
rect 13228 8984 13234 8996
rect 13633 8993 13645 8996
rect 13679 8993 13691 9027
rect 14458 9024 14464 9036
rect 14419 8996 14464 9024
rect 13633 8987 13691 8993
rect 14458 8984 14464 8996
rect 14516 8984 14522 9036
rect 11514 8956 11520 8968
rect 10520 8928 11520 8956
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 12216 8928 12541 8956
rect 12216 8916 12222 8928
rect 12529 8925 12541 8928
rect 12575 8925 12587 8959
rect 12529 8919 12587 8925
rect 12621 8959 12679 8965
rect 12621 8925 12633 8959
rect 12667 8925 12679 8959
rect 12621 8919 12679 8925
rect 7892 8860 8800 8888
rect 7892 8848 7898 8860
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 9548 8860 10088 8888
rect 9548 8848 9554 8860
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 1946 8820 1952 8832
rect 1627 8792 1952 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 2314 8780 2320 8832
rect 2372 8820 2378 8832
rect 2958 8820 2964 8832
rect 2372 8792 2964 8820
rect 2372 8780 2378 8792
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 4246 8820 4252 8832
rect 4207 8792 4252 8820
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 6914 8820 6920 8832
rect 4488 8792 6920 8820
rect 4488 8780 4494 8792
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 7374 8820 7380 8832
rect 7335 8792 7380 8820
rect 7374 8780 7380 8792
rect 7432 8820 7438 8832
rect 8846 8820 8852 8832
rect 7432 8792 8852 8820
rect 7432 8780 7438 8792
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 9674 8820 9680 8832
rect 9635 8792 9680 8820
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 10060 8820 10088 8860
rect 10778 8848 10784 8900
rect 10836 8888 10842 8900
rect 12636 8888 12664 8919
rect 12802 8916 12808 8968
rect 12860 8956 12866 8968
rect 12986 8956 12992 8968
rect 12860 8928 12992 8956
rect 12860 8916 12866 8928
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 13817 8959 13875 8965
rect 13817 8956 13829 8959
rect 13780 8928 13829 8956
rect 13780 8916 13786 8928
rect 13817 8925 13829 8928
rect 13863 8925 13875 8959
rect 13817 8919 13875 8925
rect 10836 8860 12664 8888
rect 10836 8848 10842 8860
rect 10594 8820 10600 8832
rect 10060 8792 10600 8820
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 10962 8780 10968 8832
rect 11020 8820 11026 8832
rect 11698 8820 11704 8832
rect 11020 8792 11704 8820
rect 11020 8780 11026 8792
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 12069 8823 12127 8829
rect 12069 8789 12081 8823
rect 12115 8820 12127 8823
rect 12434 8820 12440 8832
rect 12115 8792 12440 8820
rect 12115 8789 12127 8792
rect 12069 8783 12127 8789
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 14645 8823 14703 8829
rect 14645 8820 14657 8823
rect 13872 8792 14657 8820
rect 13872 8780 13878 8792
rect 14645 8789 14657 8792
rect 14691 8789 14703 8823
rect 14645 8783 14703 8789
rect 1104 8730 15824 8752
rect 1104 8678 3447 8730
rect 3499 8678 3511 8730
rect 3563 8678 3575 8730
rect 3627 8678 3639 8730
rect 3691 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 13308 8730
rect 13360 8678 13372 8730
rect 13424 8678 13436 8730
rect 13488 8678 13500 8730
rect 13552 8678 15824 8730
rect 1104 8656 15824 8678
rect 2406 8576 2412 8628
rect 2464 8616 2470 8628
rect 2464 8588 4016 8616
rect 2464 8576 2470 8588
rect 3697 8551 3755 8557
rect 3697 8548 3709 8551
rect 1596 8520 3709 8548
rect 1596 8421 1624 8520
rect 3697 8517 3709 8520
rect 3743 8517 3755 8551
rect 3988 8548 4016 8588
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 9582 8616 9588 8628
rect 4120 8588 9588 8616
rect 4120 8576 4126 8588
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 9858 8576 9864 8628
rect 9916 8616 9922 8628
rect 11057 8619 11115 8625
rect 11057 8616 11069 8619
rect 9916 8588 11069 8616
rect 9916 8576 9922 8588
rect 11057 8585 11069 8588
rect 11103 8585 11115 8619
rect 11057 8579 11115 8585
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 12437 8619 12495 8625
rect 12437 8616 12449 8619
rect 11296 8588 12449 8616
rect 11296 8576 11302 8588
rect 12437 8585 12449 8588
rect 12483 8585 12495 8619
rect 13630 8616 13636 8628
rect 13591 8588 13636 8616
rect 12437 8579 12495 8585
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 4614 8548 4620 8560
rect 3988 8520 4620 8548
rect 3697 8511 3755 8517
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 6270 8548 6276 8560
rect 6231 8520 6276 8548
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 7834 8508 7840 8560
rect 7892 8548 7898 8560
rect 8205 8551 8263 8557
rect 8205 8548 8217 8551
rect 7892 8520 8217 8548
rect 7892 8508 7898 8520
rect 8205 8517 8217 8520
rect 8251 8548 8263 8551
rect 9490 8548 9496 8560
rect 8251 8520 9496 8548
rect 8251 8517 8263 8520
rect 8205 8511 8263 8517
rect 9490 8508 9496 8520
rect 9548 8508 9554 8560
rect 11422 8508 11428 8560
rect 11480 8548 11486 8560
rect 11480 8520 11652 8548
rect 11480 8508 11486 8520
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 3602 8480 3608 8492
rect 3191 8452 3608 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 3602 8440 3608 8452
rect 3660 8440 3666 8492
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4387 8452 5028 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8381 1639 8415
rect 1581 8375 1639 8381
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8412 3019 8415
rect 3878 8412 3884 8424
rect 3007 8384 3884 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 3878 8372 3884 8384
rect 3936 8372 3942 8424
rect 4062 8412 4068 8424
rect 4023 8384 4068 8412
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4157 8415 4215 8421
rect 4157 8381 4169 8415
rect 4203 8412 4215 8415
rect 4614 8412 4620 8424
rect 4203 8384 4620 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 4798 8372 4804 8424
rect 4856 8412 4862 8424
rect 4893 8415 4951 8421
rect 4893 8412 4905 8415
rect 4856 8384 4905 8412
rect 4856 8372 4862 8384
rect 4893 8381 4905 8384
rect 4939 8381 4951 8415
rect 5000 8412 5028 8452
rect 8110 8440 8116 8492
rect 8168 8480 8174 8492
rect 9309 8483 9367 8489
rect 9309 8480 9321 8483
rect 8168 8452 9321 8480
rect 8168 8440 8174 8452
rect 9309 8449 9321 8452
rect 9355 8480 9367 8483
rect 9398 8480 9404 8492
rect 9355 8452 9404 8480
rect 9355 8449 9367 8452
rect 9309 8443 9367 8449
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 10410 8480 10416 8492
rect 10100 8452 10416 8480
rect 10100 8440 10106 8452
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 11624 8489 11652 8520
rect 12158 8508 12164 8560
rect 12216 8548 12222 8560
rect 12216 8520 13308 8548
rect 12216 8508 12222 8520
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11296 8452 11529 8480
rect 11296 8440 11302 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11609 8483 11667 8489
rect 11609 8449 11621 8483
rect 11655 8449 11667 8483
rect 11609 8443 11667 8449
rect 12618 8440 12624 8492
rect 12676 8480 12682 8492
rect 12802 8480 12808 8492
rect 12676 8452 12808 8480
rect 12676 8440 12682 8452
rect 12802 8440 12808 8452
rect 12860 8480 12866 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12860 8452 13001 8480
rect 12860 8440 12866 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 13280 8480 13308 8520
rect 13354 8508 13360 8560
rect 13412 8548 13418 8560
rect 15013 8551 15071 8557
rect 15013 8548 15025 8551
rect 13412 8520 15025 8548
rect 13412 8508 13418 8520
rect 15013 8517 15025 8520
rect 15059 8517 15071 8551
rect 15013 8511 15071 8517
rect 13722 8480 13728 8492
rect 13280 8452 13728 8480
rect 12989 8443 13047 8449
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 14182 8480 14188 8492
rect 14143 8452 14188 8480
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 6270 8412 6276 8424
rect 5000 8384 6276 8412
rect 4893 8375 4951 8381
rect 6270 8372 6276 8384
rect 6328 8372 6334 8424
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 6972 8384 9137 8412
rect 6972 8372 6978 8384
rect 9125 8381 9137 8384
rect 9171 8412 9183 8415
rect 9214 8412 9220 8424
rect 9171 8384 9220 8412
rect 9171 8381 9183 8384
rect 9125 8375 9183 8381
rect 9214 8372 9220 8384
rect 9272 8372 9278 8424
rect 10226 8412 10232 8424
rect 10187 8384 10232 8412
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 10778 8412 10784 8424
rect 10336 8384 10784 8412
rect 1210 8304 1216 8356
rect 1268 8344 1274 8356
rect 1857 8347 1915 8353
rect 1857 8344 1869 8347
rect 1268 8316 1869 8344
rect 1268 8304 1274 8316
rect 1857 8313 1869 8316
rect 1903 8313 1915 8347
rect 1857 8307 1915 8313
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8344 2927 8347
rect 4338 8344 4344 8356
rect 2915 8316 4344 8344
rect 2915 8313 2927 8316
rect 2869 8307 2927 8313
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 5160 8347 5218 8353
rect 5160 8313 5172 8347
rect 5206 8313 5218 8347
rect 5160 8307 5218 8313
rect 7092 8347 7150 8353
rect 7092 8313 7104 8347
rect 7138 8344 7150 8347
rect 7190 8344 7196 8356
rect 7138 8316 7196 8344
rect 7138 8313 7150 8316
rect 7092 8307 7150 8313
rect 1118 8236 1124 8288
rect 1176 8276 1182 8288
rect 1578 8276 1584 8288
rect 1176 8248 1584 8276
rect 1176 8236 1182 8248
rect 1578 8236 1584 8248
rect 1636 8236 1642 8288
rect 2314 8236 2320 8288
rect 2372 8276 2378 8288
rect 2501 8279 2559 8285
rect 2501 8276 2513 8279
rect 2372 8248 2513 8276
rect 2372 8236 2378 8248
rect 2501 8245 2513 8248
rect 2547 8245 2559 8279
rect 2501 8239 2559 8245
rect 2682 8236 2688 8288
rect 2740 8276 2746 8288
rect 3694 8276 3700 8288
rect 2740 8248 3700 8276
rect 2740 8236 2746 8248
rect 3694 8236 3700 8248
rect 3752 8236 3758 8288
rect 3878 8236 3884 8288
rect 3936 8276 3942 8288
rect 4890 8276 4896 8288
rect 3936 8248 4896 8276
rect 3936 8236 3942 8248
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 5184 8276 5212 8307
rect 7190 8304 7196 8316
rect 7248 8304 7254 8356
rect 9033 8347 9091 8353
rect 9033 8313 9045 8347
rect 9079 8344 9091 8347
rect 9079 8316 9352 8344
rect 9079 8313 9091 8316
rect 9033 8307 9091 8313
rect 7006 8276 7012 8288
rect 5184 8248 7012 8276
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 7374 8236 7380 8288
rect 7432 8276 7438 8288
rect 8110 8276 8116 8288
rect 7432 8248 8116 8276
rect 7432 8236 7438 8248
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 8294 8236 8300 8288
rect 8352 8276 8358 8288
rect 8665 8279 8723 8285
rect 8665 8276 8677 8279
rect 8352 8248 8677 8276
rect 8352 8236 8358 8248
rect 8665 8245 8677 8248
rect 8711 8245 8723 8279
rect 9324 8276 9352 8316
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 10336 8344 10364 8384
rect 10778 8372 10784 8384
rect 10836 8372 10842 8424
rect 13446 8412 13452 8424
rect 11624 8384 13452 8412
rect 9548 8316 10364 8344
rect 9548 8304 9554 8316
rect 10410 8304 10416 8356
rect 10468 8344 10474 8356
rect 10962 8344 10968 8356
rect 10468 8316 10968 8344
rect 10468 8304 10474 8316
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 11425 8347 11483 8353
rect 11425 8313 11437 8347
rect 11471 8344 11483 8347
rect 11514 8344 11520 8356
rect 11471 8316 11520 8344
rect 11471 8313 11483 8316
rect 11425 8307 11483 8313
rect 11514 8304 11520 8316
rect 11572 8304 11578 8356
rect 9398 8276 9404 8288
rect 9324 8248 9404 8276
rect 8665 8239 8723 8245
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 9858 8276 9864 8288
rect 9819 8248 9864 8276
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 10321 8279 10379 8285
rect 10321 8245 10333 8279
rect 10367 8276 10379 8279
rect 11624 8276 11652 8384
rect 13446 8372 13452 8384
rect 13504 8372 13510 8424
rect 13906 8412 13912 8424
rect 13556 8384 13912 8412
rect 12618 8304 12624 8356
rect 12676 8344 12682 8356
rect 12805 8347 12863 8353
rect 12805 8344 12817 8347
rect 12676 8316 12817 8344
rect 12676 8304 12682 8316
rect 12805 8313 12817 8316
rect 12851 8313 12863 8347
rect 12805 8307 12863 8313
rect 12897 8347 12955 8353
rect 12897 8313 12909 8347
rect 12943 8344 12955 8347
rect 13556 8344 13584 8384
rect 13906 8372 13912 8384
rect 13964 8412 13970 8424
rect 14550 8412 14556 8424
rect 13964 8384 14556 8412
rect 13964 8372 13970 8384
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 14829 8415 14887 8421
rect 14829 8381 14841 8415
rect 14875 8412 14887 8415
rect 14918 8412 14924 8424
rect 14875 8384 14924 8412
rect 14875 8381 14887 8384
rect 14829 8375 14887 8381
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 12943 8316 13584 8344
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 14001 8347 14059 8353
rect 14001 8344 14013 8347
rect 13780 8316 14013 8344
rect 13780 8304 13786 8316
rect 14001 8313 14013 8316
rect 14047 8313 14059 8347
rect 14001 8307 14059 8313
rect 10367 8248 11652 8276
rect 14093 8279 14151 8285
rect 10367 8245 10379 8248
rect 10321 8239 10379 8245
rect 14093 8245 14105 8279
rect 14139 8276 14151 8279
rect 14274 8276 14280 8288
rect 14139 8248 14280 8276
rect 14139 8245 14151 8248
rect 14093 8239 14151 8245
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 1104 8186 15824 8208
rect 1104 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 6104 8186
rect 6156 8134 10843 8186
rect 10895 8134 10907 8186
rect 10959 8134 10971 8186
rect 11023 8134 11035 8186
rect 11087 8134 15824 8186
rect 1104 8112 15824 8134
rect 1210 8032 1216 8084
rect 1268 8072 1274 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 1268 8044 1593 8072
rect 1268 8032 1274 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 1581 8035 1639 8041
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 4246 8072 4252 8084
rect 1995 8044 4252 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4430 8032 4436 8084
rect 4488 8072 4494 8084
rect 8294 8072 8300 8084
rect 4488 8044 8300 8072
rect 4488 8032 4494 8044
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 8938 8032 8944 8084
rect 8996 8072 9002 8084
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 8996 8044 9137 8072
rect 8996 8032 9002 8044
rect 9125 8041 9137 8044
rect 9171 8041 9183 8075
rect 9125 8035 9183 8041
rect 9582 8032 9588 8084
rect 9640 8072 9646 8084
rect 9677 8075 9735 8081
rect 9677 8072 9689 8075
rect 9640 8044 9689 8072
rect 9640 8032 9646 8044
rect 9677 8041 9689 8044
rect 9723 8041 9735 8075
rect 9677 8035 9735 8041
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 9916 8044 10149 8072
rect 9916 8032 9922 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8041 10931 8075
rect 10873 8035 10931 8041
rect 11241 8075 11299 8081
rect 11241 8041 11253 8075
rect 11287 8041 11299 8075
rect 11241 8035 11299 8041
rect 11333 8075 11391 8081
rect 11333 8041 11345 8075
rect 11379 8072 11391 8075
rect 11422 8072 11428 8084
rect 11379 8044 11428 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 2041 8007 2099 8013
rect 2041 7973 2053 8007
rect 2087 8004 2099 8007
rect 2682 8004 2688 8016
rect 2087 7976 2688 8004
rect 2087 7973 2099 7976
rect 2041 7967 2099 7973
rect 2682 7964 2688 7976
rect 2740 7964 2746 8016
rect 3145 8007 3203 8013
rect 3145 7973 3157 8007
rect 3191 8004 3203 8007
rect 10888 8004 10916 8035
rect 3191 7976 10916 8004
rect 11256 8004 11284 8035
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 12069 8075 12127 8081
rect 12069 8072 12081 8075
rect 11572 8044 12081 8072
rect 11572 8032 11578 8044
rect 12069 8041 12081 8044
rect 12115 8041 12127 8075
rect 12069 8035 12127 8041
rect 13078 8032 13084 8084
rect 13136 8072 13142 8084
rect 13354 8072 13360 8084
rect 13136 8044 13360 8072
rect 13136 8032 13142 8044
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 13725 8075 13783 8081
rect 13725 8072 13737 8075
rect 13504 8044 13737 8072
rect 13504 8032 13510 8044
rect 13725 8041 13737 8044
rect 13771 8041 13783 8075
rect 13725 8035 13783 8041
rect 11256 7976 11652 8004
rect 3191 7973 3203 7976
rect 3145 7967 3203 7973
rect 3878 7936 3884 7948
rect 2240 7908 3884 7936
rect 2240 7877 2268 7908
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 4338 7945 4344 7948
rect 4332 7936 4344 7945
rect 4299 7908 4344 7936
rect 4332 7899 4344 7908
rect 4338 7896 4344 7899
rect 4396 7896 4402 7948
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 6161 7939 6219 7945
rect 6161 7936 6173 7939
rect 4948 7908 6173 7936
rect 4948 7896 4954 7908
rect 6161 7905 6173 7908
rect 6207 7936 6219 7939
rect 7834 7936 7840 7948
rect 6207 7908 7840 7936
rect 6207 7905 6219 7908
rect 6161 7899 6219 7905
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 8012 7939 8070 7945
rect 8012 7905 8024 7939
rect 8058 7936 8070 7939
rect 8058 7908 8892 7936
rect 8058 7905 8070 7908
rect 8012 7899 8070 7905
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7837 2283 7871
rect 3234 7868 3240 7880
rect 3195 7840 3240 7868
rect 2225 7831 2283 7837
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7868 3479 7871
rect 4062 7868 4068 7880
rect 3467 7840 3924 7868
rect 4023 7840 4068 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 3896 7812 3924 7840
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 3510 7800 3516 7812
rect 2240 7772 3516 7800
rect 2240 7744 2268 7772
rect 3510 7760 3516 7772
rect 3568 7760 3574 7812
rect 3878 7760 3884 7812
rect 3936 7760 3942 7812
rect 5368 7772 5948 7800
rect 2222 7692 2228 7744
rect 2280 7692 2286 7744
rect 2777 7735 2835 7741
rect 2777 7701 2789 7735
rect 2823 7732 2835 7735
rect 5368 7732 5396 7772
rect 2823 7704 5396 7732
rect 2823 7701 2835 7704
rect 2777 7695 2835 7701
rect 5442 7692 5448 7744
rect 5500 7732 5506 7744
rect 5920 7732 5948 7772
rect 7098 7760 7104 7812
rect 7156 7800 7162 7812
rect 7285 7803 7343 7809
rect 7285 7800 7297 7803
rect 7156 7772 7297 7800
rect 7156 7760 7162 7772
rect 7285 7769 7297 7772
rect 7331 7769 7343 7803
rect 7285 7763 7343 7769
rect 7558 7732 7564 7744
rect 5500 7704 5545 7732
rect 5920 7704 7564 7732
rect 5500 7692 5506 7704
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 7650 7692 7656 7744
rect 7708 7732 7714 7744
rect 7760 7732 7788 7831
rect 8864 7800 8892 7908
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 9398 7936 9404 7948
rect 9180 7908 9404 7936
rect 9180 7896 9186 7908
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 10045 7939 10103 7945
rect 10045 7905 10057 7939
rect 10091 7936 10103 7939
rect 11624 7936 11652 7976
rect 11698 7964 11704 8016
rect 11756 8004 11762 8016
rect 11756 7976 12664 8004
rect 11756 7964 11762 7976
rect 12066 7936 12072 7948
rect 10091 7908 11560 7936
rect 11624 7908 12072 7936
rect 10091 7905 10103 7908
rect 10045 7899 10103 7905
rect 8938 7828 8944 7880
rect 8996 7868 9002 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 8996 7840 10333 7868
rect 8996 7828 9002 7840
rect 10321 7837 10333 7840
rect 10367 7868 10379 7871
rect 10962 7868 10968 7880
rect 10367 7840 10968 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11422 7868 11428 7880
rect 11383 7840 11428 7868
rect 11422 7828 11428 7840
rect 11480 7828 11486 7880
rect 11532 7868 11560 7908
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 12250 7896 12256 7948
rect 12308 7936 12314 7948
rect 12434 7936 12440 7948
rect 12308 7908 12440 7936
rect 12308 7896 12314 7908
rect 12434 7896 12440 7908
rect 12492 7896 12498 7948
rect 12636 7936 12664 7976
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 12768 7976 14504 8004
rect 12768 7964 12774 7976
rect 12636 7908 12940 7936
rect 12526 7868 12532 7880
rect 11532 7840 12296 7868
rect 12487 7840 12532 7868
rect 12158 7800 12164 7812
rect 8864 7772 12164 7800
rect 12158 7760 12164 7772
rect 12216 7760 12222 7812
rect 12268 7744 12296 7840
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7868 12771 7871
rect 12802 7868 12808 7880
rect 12759 7840 12808 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 12912 7868 12940 7908
rect 13170 7896 13176 7948
rect 13228 7936 13234 7948
rect 14476 7945 14504 7976
rect 13633 7939 13691 7945
rect 13633 7936 13645 7939
rect 13228 7908 13645 7936
rect 13228 7896 13234 7908
rect 13633 7905 13645 7908
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 14461 7939 14519 7945
rect 14461 7905 14473 7939
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 13817 7871 13875 7877
rect 13817 7868 13829 7871
rect 12912 7840 13829 7868
rect 13817 7837 13829 7840
rect 13863 7868 13875 7871
rect 14182 7868 14188 7880
rect 13863 7840 14188 7868
rect 13863 7837 13875 7840
rect 13817 7831 13875 7837
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 13446 7800 13452 7812
rect 12544 7772 13452 7800
rect 12544 7744 12572 7772
rect 13446 7760 13452 7772
rect 13504 7760 13510 7812
rect 13538 7760 13544 7812
rect 13596 7800 13602 7812
rect 14918 7800 14924 7812
rect 13596 7772 14924 7800
rect 13596 7760 13602 7772
rect 14918 7760 14924 7772
rect 14976 7760 14982 7812
rect 9030 7732 9036 7744
rect 7708 7704 9036 7732
rect 7708 7692 7714 7704
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9674 7692 9680 7744
rect 9732 7732 9738 7744
rect 10226 7732 10232 7744
rect 9732 7704 10232 7732
rect 9732 7692 9738 7704
rect 10226 7692 10232 7704
rect 10284 7692 10290 7744
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 11698 7732 11704 7744
rect 10652 7704 11704 7732
rect 10652 7692 10658 7704
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 12250 7692 12256 7744
rect 12308 7692 12314 7744
rect 12526 7692 12532 7744
rect 12584 7692 12590 7744
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 13265 7735 13323 7741
rect 13265 7732 13277 7735
rect 12860 7704 13277 7732
rect 12860 7692 12866 7704
rect 13265 7701 13277 7704
rect 13311 7701 13323 7735
rect 13265 7695 13323 7701
rect 13630 7692 13636 7744
rect 13688 7732 13694 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 13688 7704 14657 7732
rect 13688 7692 13694 7704
rect 14645 7701 14657 7704
rect 14691 7701 14703 7735
rect 14645 7695 14703 7701
rect 1104 7642 15824 7664
rect 1104 7590 3447 7642
rect 3499 7590 3511 7642
rect 3563 7590 3575 7642
rect 3627 7590 3639 7642
rect 3691 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 13308 7642
rect 13360 7590 13372 7642
rect 13424 7590 13436 7642
rect 13488 7590 13500 7642
rect 13552 7590 15824 7642
rect 1104 7568 15824 7590
rect 1670 7488 1676 7540
rect 1728 7528 1734 7540
rect 1857 7531 1915 7537
rect 1857 7528 1869 7531
rect 1728 7500 1869 7528
rect 1728 7488 1734 7500
rect 1857 7497 1869 7500
rect 1903 7497 1915 7531
rect 4338 7528 4344 7540
rect 1857 7491 1915 7497
rect 3068 7500 4344 7528
rect 1486 7352 1492 7404
rect 1544 7352 1550 7404
rect 2314 7392 2320 7404
rect 2275 7364 2320 7392
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 3068 7392 3096 7500
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 6270 7528 6276 7540
rect 6231 7500 6276 7528
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 7466 7528 7472 7540
rect 6380 7500 7472 7528
rect 4433 7463 4491 7469
rect 4433 7429 4445 7463
rect 4479 7460 4491 7463
rect 4706 7460 4712 7472
rect 4479 7432 4712 7460
rect 4479 7429 4491 7432
rect 4433 7423 4491 7429
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 6380 7460 6408 7500
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 7616 7500 10824 7528
rect 7616 7488 7622 7500
rect 5920 7432 6408 7460
rect 2547 7364 3096 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 1504 7200 1532 7352
rect 2222 7324 2228 7336
rect 2183 7296 2228 7324
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 3050 7324 3056 7336
rect 3011 7296 3056 7324
rect 3050 7284 3056 7296
rect 3108 7324 3114 7336
rect 4062 7324 4068 7336
rect 3108 7296 4068 7324
rect 3108 7284 3114 7296
rect 4062 7284 4068 7296
rect 4120 7324 4126 7336
rect 4890 7324 4896 7336
rect 4120 7296 4896 7324
rect 4120 7284 4126 7296
rect 4890 7284 4896 7296
rect 4948 7284 4954 7336
rect 5920 7324 5948 7432
rect 8110 7420 8116 7472
rect 8168 7460 8174 7472
rect 8205 7463 8263 7469
rect 8205 7460 8217 7463
rect 8168 7432 8217 7460
rect 8168 7420 8174 7432
rect 8205 7429 8217 7432
rect 8251 7429 8263 7463
rect 8205 7423 8263 7429
rect 9858 7420 9864 7472
rect 9916 7460 9922 7472
rect 9916 7432 10732 7460
rect 9916 7420 9922 7432
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6328 7364 6960 7392
rect 6328 7352 6334 7364
rect 5092 7296 5948 7324
rect 3320 7259 3378 7265
rect 3320 7225 3332 7259
rect 3366 7256 3378 7259
rect 5092 7256 5120 7296
rect 5994 7284 6000 7336
rect 6052 7324 6058 7336
rect 6822 7324 6828 7336
rect 6052 7296 6828 7324
rect 6052 7284 6058 7296
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 6932 7324 6960 7364
rect 8478 7352 8484 7404
rect 8536 7392 8542 7404
rect 8536 7364 8800 7392
rect 8536 7352 8542 7364
rect 7081 7327 7139 7333
rect 7081 7324 7093 7327
rect 6932 7296 7093 7324
rect 7081 7293 7093 7296
rect 7127 7293 7139 7327
rect 7081 7287 7139 7293
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7293 8723 7327
rect 8772 7324 8800 7364
rect 10134 7352 10140 7404
rect 10192 7392 10198 7404
rect 10410 7392 10416 7404
rect 10192 7364 10416 7392
rect 10192 7352 10198 7364
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 8921 7327 8979 7333
rect 8921 7324 8933 7327
rect 8772 7296 8933 7324
rect 8665 7287 8723 7293
rect 8921 7293 8933 7296
rect 8967 7324 8979 7327
rect 9490 7324 9496 7336
rect 8967 7296 9496 7324
rect 8967 7293 8979 7296
rect 8921 7287 8979 7293
rect 3366 7228 5120 7256
rect 5160 7259 5218 7265
rect 3366 7225 3378 7228
rect 3320 7219 3378 7225
rect 5160 7225 5172 7259
rect 5206 7256 5218 7259
rect 8570 7256 8576 7268
rect 5206 7228 7144 7256
rect 5206 7225 5218 7228
rect 5160 7219 5218 7225
rect 1486 7148 1492 7200
rect 1544 7148 1550 7200
rect 3878 7148 3884 7200
rect 3936 7188 3942 7200
rect 6270 7188 6276 7200
rect 3936 7160 6276 7188
rect 3936 7148 3942 7160
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 7116 7188 7144 7228
rect 8128 7228 8576 7256
rect 8128 7188 8156 7228
rect 8570 7216 8576 7228
rect 8628 7216 8634 7268
rect 8680 7256 8708 7287
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 10226 7284 10232 7336
rect 10284 7324 10290 7336
rect 10284 7296 10640 7324
rect 10284 7284 10290 7296
rect 9030 7256 9036 7268
rect 8680 7228 9036 7256
rect 9030 7216 9036 7228
rect 9088 7216 9094 7268
rect 9122 7216 9128 7268
rect 9180 7256 9186 7268
rect 9180 7228 10548 7256
rect 9180 7216 9186 7228
rect 7116 7160 8156 7188
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 9858 7188 9864 7200
rect 8260 7160 9864 7188
rect 8260 7148 8266 7160
rect 9858 7148 9864 7160
rect 9916 7188 9922 7200
rect 10520 7197 10548 7228
rect 10045 7191 10103 7197
rect 10045 7188 10057 7191
rect 9916 7160 10057 7188
rect 9916 7148 9922 7160
rect 10045 7157 10057 7160
rect 10091 7157 10103 7191
rect 10045 7151 10103 7157
rect 10505 7191 10563 7197
rect 10505 7157 10517 7191
rect 10551 7157 10563 7191
rect 10612 7188 10640 7296
rect 10704 7256 10732 7432
rect 10796 7324 10824 7500
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 11330 7528 11336 7540
rect 11112 7500 11336 7528
rect 11112 7488 11118 7500
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 11698 7488 11704 7540
rect 11756 7528 11762 7540
rect 12986 7528 12992 7540
rect 11756 7500 12992 7528
rect 11756 7488 11762 7500
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 10962 7420 10968 7472
rect 11020 7460 11026 7472
rect 11020 7432 11100 7460
rect 11020 7420 11026 7432
rect 11072 7401 11100 7432
rect 11146 7420 11152 7472
rect 11204 7460 11210 7472
rect 12437 7463 12495 7469
rect 12437 7460 12449 7463
rect 11204 7432 12449 7460
rect 11204 7420 11210 7432
rect 12437 7429 12449 7432
rect 12483 7429 12495 7463
rect 12437 7423 12495 7429
rect 12710 7420 12716 7472
rect 12768 7460 12774 7472
rect 13998 7460 14004 7472
rect 12768 7432 14004 7460
rect 12768 7420 12774 7432
rect 13998 7420 14004 7432
rect 14056 7420 14062 7472
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7361 11115 7395
rect 11698 7392 11704 7404
rect 11057 7355 11115 7361
rect 11164 7364 11704 7392
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 10796 7296 10977 7324
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 11164 7324 11192 7364
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12526 7392 12532 7404
rect 12124 7364 12532 7392
rect 12124 7352 12130 7364
rect 12526 7352 12532 7364
rect 12584 7352 12590 7404
rect 12894 7392 12900 7404
rect 12855 7364 12900 7392
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 14185 7395 14243 7401
rect 13044 7364 13089 7392
rect 13044 7352 13050 7364
rect 14185 7361 14197 7395
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 14200 7324 14228 7355
rect 10965 7287 11023 7293
rect 11072 7296 11192 7324
rect 11256 7296 14228 7324
rect 14829 7327 14887 7333
rect 11072 7256 11100 7296
rect 11256 7256 11284 7296
rect 14829 7293 14841 7327
rect 14875 7324 14887 7327
rect 14918 7324 14924 7336
rect 14875 7296 14924 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 14001 7259 14059 7265
rect 14001 7256 14013 7259
rect 10704 7228 11100 7256
rect 11164 7228 11284 7256
rect 13096 7228 14013 7256
rect 11164 7200 11192 7228
rect 10873 7191 10931 7197
rect 10873 7188 10885 7191
rect 10612 7160 10885 7188
rect 10505 7151 10563 7157
rect 10873 7157 10885 7160
rect 10919 7157 10931 7191
rect 10873 7151 10931 7157
rect 11146 7148 11152 7200
rect 11204 7148 11210 7200
rect 11701 7191 11759 7197
rect 11701 7157 11713 7191
rect 11747 7188 11759 7191
rect 12342 7188 12348 7200
rect 11747 7160 12348 7188
rect 11747 7157 11759 7160
rect 11701 7151 11759 7157
rect 12342 7148 12348 7160
rect 12400 7148 12406 7200
rect 12710 7148 12716 7200
rect 12768 7188 12774 7200
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 12768 7160 12817 7188
rect 12768 7148 12774 7160
rect 12805 7157 12817 7160
rect 12851 7157 12863 7191
rect 12805 7151 12863 7157
rect 12894 7148 12900 7200
rect 12952 7188 12958 7200
rect 13096 7188 13124 7228
rect 14001 7225 14013 7228
rect 14047 7225 14059 7259
rect 14001 7219 14059 7225
rect 13630 7188 13636 7200
rect 12952 7160 13124 7188
rect 13591 7160 13636 7188
rect 12952 7148 12958 7160
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 14093 7191 14151 7197
rect 14093 7157 14105 7191
rect 14139 7188 14151 7191
rect 14826 7188 14832 7200
rect 14139 7160 14832 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 14826 7148 14832 7160
rect 14884 7148 14890 7200
rect 14918 7148 14924 7200
rect 14976 7188 14982 7200
rect 15013 7191 15071 7197
rect 15013 7188 15025 7191
rect 14976 7160 15025 7188
rect 14976 7148 14982 7160
rect 15013 7157 15025 7160
rect 15059 7157 15071 7191
rect 15013 7151 15071 7157
rect 1104 7098 15824 7120
rect 1104 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 6104 7098
rect 6156 7046 10843 7098
rect 10895 7046 10907 7098
rect 10959 7046 10971 7098
rect 11023 7046 11035 7098
rect 11087 7046 15824 7098
rect 1104 7024 15824 7046
rect 3513 6987 3571 6993
rect 3513 6953 3525 6987
rect 3559 6984 3571 6987
rect 7006 6984 7012 6996
rect 3559 6956 7012 6984
rect 3559 6953 3571 6956
rect 3513 6947 3571 6953
rect 7006 6944 7012 6956
rect 7064 6944 7070 6996
rect 7101 6987 7159 6993
rect 7101 6953 7113 6987
rect 7147 6984 7159 6987
rect 8386 6984 8392 6996
rect 7147 6956 8392 6984
rect 7147 6953 7159 6956
rect 7101 6947 7159 6953
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 8938 6984 8944 6996
rect 8628 6956 8944 6984
rect 8628 6944 8634 6956
rect 8938 6944 8944 6956
rect 8996 6944 9002 6996
rect 9122 6944 9128 6996
rect 9180 6984 9186 6996
rect 10042 6984 10048 6996
rect 9180 6956 10048 6984
rect 9180 6944 9186 6956
rect 10042 6944 10048 6956
rect 10100 6984 10106 6996
rect 10100 6956 10272 6984
rect 10100 6944 10106 6956
rect 2314 6876 2320 6928
rect 2372 6876 2378 6928
rect 4338 6876 4344 6928
rect 4396 6916 4402 6928
rect 9766 6916 9772 6928
rect 4396 6888 9772 6916
rect 4396 6876 4402 6888
rect 9766 6876 9772 6888
rect 9824 6876 9830 6928
rect 10134 6916 10140 6928
rect 10095 6888 10140 6916
rect 10134 6876 10140 6888
rect 10192 6876 10198 6928
rect 10244 6916 10272 6956
rect 10410 6944 10416 6996
rect 10468 6984 10474 6996
rect 10873 6987 10931 6993
rect 10873 6984 10885 6987
rect 10468 6956 10885 6984
rect 10468 6944 10474 6956
rect 10873 6953 10885 6956
rect 10919 6953 10931 6987
rect 10873 6947 10931 6953
rect 12069 6987 12127 6993
rect 12069 6953 12081 6987
rect 12115 6984 12127 6987
rect 12250 6984 12256 6996
rect 12115 6956 12256 6984
rect 12115 6953 12127 6956
rect 12069 6947 12127 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 12437 6987 12495 6993
rect 12437 6984 12449 6987
rect 12400 6956 12449 6984
rect 12400 6944 12406 6956
rect 12437 6953 12449 6956
rect 12483 6953 12495 6987
rect 12437 6947 12495 6953
rect 12529 6987 12587 6993
rect 12529 6953 12541 6987
rect 12575 6984 12587 6987
rect 12802 6984 12808 6996
rect 12575 6956 12808 6984
rect 12575 6953 12587 6956
rect 12529 6947 12587 6953
rect 12802 6944 12808 6956
rect 12860 6944 12866 6996
rect 11241 6919 11299 6925
rect 11241 6916 11253 6919
rect 10244 6888 11253 6916
rect 11241 6885 11253 6888
rect 11287 6885 11299 6919
rect 11241 6879 11299 6885
rect 11333 6919 11391 6925
rect 11333 6885 11345 6919
rect 11379 6916 11391 6919
rect 11606 6916 11612 6928
rect 11379 6888 11612 6916
rect 11379 6885 11391 6888
rect 11333 6879 11391 6885
rect 11606 6876 11612 6888
rect 11664 6876 11670 6928
rect 13633 6919 13691 6925
rect 13633 6885 13645 6919
rect 13679 6916 13691 6919
rect 13722 6916 13728 6928
rect 13679 6888 13728 6916
rect 13679 6885 13691 6888
rect 13633 6879 13691 6885
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2332 6848 2360 6876
rect 1443 6820 2360 6848
rect 2400 6851 2458 6857
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2400 6817 2412 6851
rect 2446 6848 2458 6851
rect 2446 6820 3924 6848
rect 2446 6817 2458 6820
rect 2400 6811 2458 6817
rect 1486 6740 1492 6792
rect 1544 6780 1550 6792
rect 1854 6780 1860 6792
rect 1544 6752 1860 6780
rect 1544 6740 1550 6752
rect 1854 6740 1860 6752
rect 1912 6740 1918 6792
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 3896 6780 3924 6820
rect 3970 6808 3976 6860
rect 4028 6848 4034 6860
rect 4249 6851 4307 6857
rect 4249 6848 4261 6851
rect 4028 6820 4261 6848
rect 4028 6808 4034 6820
rect 4249 6817 4261 6820
rect 4295 6817 4307 6851
rect 5074 6848 5080 6860
rect 5035 6820 5080 6848
rect 4249 6811 4307 6817
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 5988 6851 6046 6857
rect 5988 6817 6000 6851
rect 6034 6848 6046 6851
rect 7650 6848 7656 6860
rect 6034 6820 7656 6848
rect 6034 6817 6046 6820
rect 5988 6811 6046 6817
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 7834 6857 7840 6860
rect 7828 6848 7840 6857
rect 7795 6820 7840 6848
rect 7828 6811 7840 6820
rect 7834 6808 7840 6811
rect 7892 6808 7898 6860
rect 8386 6808 8392 6860
rect 8444 6848 8450 6860
rect 8938 6848 8944 6860
rect 8444 6820 8944 6848
rect 8444 6808 8450 6820
rect 8938 6808 8944 6820
rect 8996 6848 9002 6860
rect 8996 6820 9987 6848
rect 8996 6808 9002 6820
rect 4706 6780 4712 6792
rect 3896 6752 4712 6780
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 4948 6752 5733 6780
rect 4948 6740 4954 6752
rect 5721 6749 5733 6752
rect 5767 6749 5779 6783
rect 7558 6780 7564 6792
rect 7519 6752 7564 6780
rect 5721 6743 5779 6749
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9674 6780 9680 6792
rect 9456 6752 9680 6780
rect 9456 6740 9462 6752
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 9959 6712 9987 6820
rect 10410 6808 10416 6860
rect 10468 6848 10474 6860
rect 10962 6848 10968 6860
rect 10468 6820 10968 6848
rect 10468 6808 10474 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11698 6808 11704 6860
rect 11756 6848 11762 6860
rect 14458 6848 14464 6860
rect 11756 6820 13860 6848
rect 14419 6820 14464 6848
rect 11756 6808 11762 6820
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 10192 6752 10241 6780
rect 10192 6740 10198 6752
rect 10229 6749 10241 6752
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 11422 6780 11428 6792
rect 10560 6752 11428 6780
rect 10560 6740 10566 6752
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11606 6740 11612 6792
rect 11664 6780 11670 6792
rect 12621 6783 12679 6789
rect 12621 6780 12633 6783
rect 11664 6752 12633 6780
rect 11664 6740 11670 6752
rect 12621 6749 12633 6752
rect 12667 6749 12679 6783
rect 12621 6743 12679 6749
rect 12802 6740 12808 6792
rect 12860 6780 12866 6792
rect 13832 6789 13860 6820
rect 14458 6808 14464 6820
rect 14516 6848 14522 6860
rect 14642 6848 14648 6860
rect 14516 6820 14648 6848
rect 14516 6808 14522 6820
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 13725 6783 13783 6789
rect 13725 6780 13737 6783
rect 12860 6752 13737 6780
rect 12860 6740 12866 6752
rect 13725 6749 13737 6752
rect 13771 6749 13783 6783
rect 13725 6743 13783 6749
rect 13817 6783 13875 6789
rect 13817 6749 13829 6783
rect 13863 6749 13875 6783
rect 13817 6743 13875 6749
rect 11054 6712 11060 6724
rect 8720 6684 9904 6712
rect 9959 6684 11060 6712
rect 8720 6672 8726 6684
rect 1486 6604 1492 6656
rect 1544 6644 1550 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1544 6616 1593 6644
rect 1544 6604 1550 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 5258 6644 5264 6656
rect 4764 6616 5264 6644
rect 4764 6604 4770 6616
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 5442 6604 5448 6656
rect 5500 6644 5506 6656
rect 9214 6644 9220 6656
rect 5500 6616 9220 6644
rect 5500 6604 5506 6616
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 9876 6644 9904 6684
rect 11054 6672 11060 6684
rect 11112 6672 11118 6724
rect 11146 6672 11152 6724
rect 11204 6712 11210 6724
rect 14645 6715 14703 6721
rect 14645 6712 14657 6715
rect 11204 6684 14657 6712
rect 11204 6672 11210 6684
rect 14645 6681 14657 6684
rect 14691 6681 14703 6715
rect 14645 6675 14703 6681
rect 13265 6647 13323 6653
rect 13265 6644 13277 6647
rect 9732 6616 9777 6644
rect 9876 6616 13277 6644
rect 9732 6604 9738 6616
rect 13265 6613 13277 6616
rect 13311 6613 13323 6647
rect 13265 6607 13323 6613
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 1857 6443 1915 6449
rect 1857 6409 1869 6443
rect 1903 6440 1915 6443
rect 3234 6440 3240 6452
rect 1903 6412 3240 6440
rect 1903 6409 1915 6412
rect 1857 6403 1915 6409
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4433 6443 4491 6449
rect 4433 6440 4445 6443
rect 4212 6412 4445 6440
rect 4212 6400 4218 6412
rect 4433 6409 4445 6412
rect 4479 6409 4491 6443
rect 8202 6440 8208 6452
rect 4433 6403 4491 6409
rect 4816 6412 8208 6440
rect 2130 6332 2136 6384
rect 2188 6372 2194 6384
rect 2188 6344 3004 6372
rect 2188 6332 2194 6344
rect 2409 6307 2467 6313
rect 2409 6304 2421 6307
rect 2148 6276 2421 6304
rect 2148 6168 2176 6276
rect 2409 6273 2421 6276
rect 2455 6273 2467 6307
rect 2409 6267 2467 6273
rect 2222 6196 2228 6248
rect 2280 6236 2286 6248
rect 2976 6236 3004 6344
rect 3050 6236 3056 6248
rect 2280 6208 2325 6236
rect 2963 6208 3056 6236
rect 2280 6196 2286 6208
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 3320 6239 3378 6245
rect 3320 6205 3332 6239
rect 3366 6236 3378 6239
rect 4816 6236 4844 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 9088 6412 9628 6440
rect 9088 6400 9094 6412
rect 6270 6372 6276 6384
rect 6231 6344 6276 6372
rect 6270 6332 6276 6344
rect 6328 6332 6334 6384
rect 9600 6372 9628 6412
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 9824 6412 10057 6440
rect 9824 6400 9830 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10045 6403 10103 6409
rect 10318 6400 10324 6452
rect 10376 6440 10382 6452
rect 12434 6440 12440 6452
rect 10376 6412 11100 6440
rect 12395 6412 12440 6440
rect 10376 6400 10382 6412
rect 10505 6375 10563 6381
rect 10505 6372 10517 6375
rect 9600 6344 10517 6372
rect 10505 6341 10517 6344
rect 10551 6341 10563 6375
rect 11072 6372 11100 6412
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 11072 6344 12664 6372
rect 10505 6335 10563 6341
rect 4890 6264 4896 6316
rect 4948 6304 4954 6316
rect 4948 6276 4993 6304
rect 4948 6264 4954 6276
rect 7834 6264 7840 6316
rect 7892 6304 7898 6316
rect 7892 6276 8800 6304
rect 7892 6264 7898 6276
rect 6822 6236 6828 6248
rect 3366 6208 4844 6236
rect 6735 6208 6828 6236
rect 3366 6205 3378 6208
rect 3320 6199 3378 6205
rect 6822 6196 6828 6208
rect 6880 6236 6886 6248
rect 7558 6236 7564 6248
rect 6880 6208 7564 6236
rect 6880 6196 6886 6208
rect 7558 6196 7564 6208
rect 7616 6236 7622 6248
rect 8665 6239 8723 6245
rect 8665 6236 8677 6239
rect 7616 6208 8677 6236
rect 7616 6196 7622 6208
rect 8665 6205 8677 6208
rect 8711 6205 8723 6239
rect 8772 6236 8800 6276
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 11057 6307 11115 6313
rect 11057 6304 11069 6307
rect 10284 6276 11069 6304
rect 10284 6264 10290 6276
rect 11057 6273 11069 6276
rect 11103 6273 11115 6307
rect 11057 6267 11115 6273
rect 11701 6307 11759 6313
rect 11701 6273 11713 6307
rect 11747 6304 11759 6307
rect 12526 6304 12532 6316
rect 11747 6276 12532 6304
rect 11747 6273 11759 6276
rect 11701 6267 11759 6273
rect 12526 6264 12532 6276
rect 12584 6264 12590 6316
rect 12636 6304 12664 6344
rect 12710 6332 12716 6384
rect 12768 6372 12774 6384
rect 12768 6344 13124 6372
rect 12768 6332 12774 6344
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12636 6276 13001 6304
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 13096 6248 13124 6344
rect 14274 6304 14280 6316
rect 14235 6276 14280 6304
rect 14274 6264 14280 6276
rect 14332 6264 14338 6316
rect 8921 6239 8979 6245
rect 8921 6236 8933 6239
rect 8772 6208 8933 6236
rect 8665 6199 8723 6205
rect 8921 6205 8933 6208
rect 8967 6236 8979 6239
rect 10318 6236 10324 6248
rect 8967 6208 10324 6236
rect 8967 6205 8979 6208
rect 8921 6199 8979 6205
rect 10318 6196 10324 6208
rect 10376 6196 10382 6248
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 10652 6208 10885 6236
rect 10652 6196 10658 6208
rect 10873 6205 10885 6208
rect 10919 6205 10931 6239
rect 10873 6199 10931 6205
rect 10962 6196 10968 6248
rect 11020 6236 11026 6248
rect 11020 6208 11065 6236
rect 11020 6196 11026 6208
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 12897 6239 12955 6245
rect 12897 6236 12909 6239
rect 12492 6208 12909 6236
rect 12492 6196 12498 6208
rect 12897 6205 12909 6208
rect 12943 6205 12955 6239
rect 12897 6199 12955 6205
rect 13078 6196 13084 6248
rect 13136 6196 13142 6248
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6236 14887 6239
rect 15470 6236 15476 6248
rect 14875 6208 15476 6236
rect 14875 6205 14887 6208
rect 14829 6199 14887 6205
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 5138 6171 5196 6177
rect 5138 6168 5150 6171
rect 2148 6140 5150 6168
rect 5138 6137 5150 6140
rect 5184 6168 5196 6171
rect 5442 6168 5448 6180
rect 5184 6140 5448 6168
rect 5184 6137 5196 6140
rect 5138 6131 5196 6137
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 5534 6128 5540 6180
rect 5592 6168 5598 6180
rect 6454 6168 6460 6180
rect 5592 6140 6460 6168
rect 5592 6128 5598 6140
rect 6454 6128 6460 6140
rect 6512 6128 6518 6180
rect 7092 6171 7150 6177
rect 7092 6137 7104 6171
rect 7138 6168 7150 6171
rect 8110 6168 8116 6180
rect 7138 6140 8116 6168
rect 7138 6137 7150 6140
rect 7092 6131 7150 6137
rect 8110 6128 8116 6140
rect 8168 6128 8174 6180
rect 9490 6128 9496 6180
rect 9548 6168 9554 6180
rect 13354 6168 13360 6180
rect 9548 6140 10824 6168
rect 9548 6128 9554 6140
rect 1302 6060 1308 6112
rect 1360 6100 1366 6112
rect 2317 6103 2375 6109
rect 2317 6100 2329 6103
rect 1360 6072 2329 6100
rect 1360 6060 1366 6072
rect 2317 6069 2329 6072
rect 2363 6100 2375 6103
rect 3878 6100 3884 6112
rect 2363 6072 3884 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 3878 6060 3884 6072
rect 3936 6060 3942 6112
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 7558 6100 7564 6112
rect 4212 6072 7564 6100
rect 4212 6060 4218 6072
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 7650 6060 7656 6112
rect 7708 6100 7714 6112
rect 8202 6100 8208 6112
rect 7708 6072 8208 6100
rect 7708 6060 7714 6072
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 10686 6100 10692 6112
rect 8628 6072 10692 6100
rect 8628 6060 8634 6072
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 10796 6100 10824 6140
rect 12636 6140 13360 6168
rect 12636 6100 12664 6140
rect 13354 6128 13360 6140
rect 13412 6128 13418 6180
rect 14093 6171 14151 6177
rect 14093 6137 14105 6171
rect 14139 6168 14151 6171
rect 15102 6168 15108 6180
rect 14139 6140 15108 6168
rect 14139 6137 14151 6140
rect 14093 6131 14151 6137
rect 15102 6128 15108 6140
rect 15160 6128 15166 6180
rect 10796 6072 12664 6100
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 12768 6072 12817 6100
rect 12768 6060 12774 6072
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 13630 6100 13636 6112
rect 13591 6072 13636 6100
rect 12805 6063 12863 6069
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14001 6103 14059 6109
rect 14001 6100 14013 6103
rect 13872 6072 14013 6100
rect 13872 6060 13878 6072
rect 14001 6069 14013 6072
rect 14047 6069 14059 6103
rect 14001 6063 14059 6069
rect 14182 6060 14188 6112
rect 14240 6100 14246 6112
rect 15013 6103 15071 6109
rect 15013 6100 15025 6103
rect 14240 6072 15025 6100
rect 14240 6060 14246 6072
rect 15013 6069 15025 6072
rect 15059 6069 15071 6103
rect 15013 6063 15071 6069
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 4617 5899 4675 5905
rect 4617 5865 4629 5899
rect 4663 5896 4675 5899
rect 4663 5868 9076 5896
rect 4663 5865 4675 5868
rect 4617 5859 4675 5865
rect 2222 5828 2228 5840
rect 1412 5800 2228 5828
rect 1412 5769 1440 5800
rect 2222 5788 2228 5800
rect 2280 5788 2286 5840
rect 4709 5831 4767 5837
rect 4709 5797 4721 5831
rect 4755 5828 4767 5831
rect 5534 5828 5540 5840
rect 4755 5800 5540 5828
rect 4755 5797 4767 5800
rect 4709 5791 4767 5797
rect 5534 5788 5540 5800
rect 5592 5788 5598 5840
rect 5626 5788 5632 5840
rect 5684 5837 5690 5840
rect 5684 5831 5748 5837
rect 5684 5797 5702 5831
rect 5736 5797 5748 5831
rect 5684 5791 5748 5797
rect 5684 5788 5690 5791
rect 7282 5788 7288 5840
rect 7340 5828 7346 5840
rect 8570 5828 8576 5840
rect 7340 5800 8576 5828
rect 7340 5788 7346 5800
rect 8570 5788 8576 5800
rect 8628 5788 8634 5840
rect 9048 5828 9076 5868
rect 10042 5856 10048 5908
rect 10100 5896 10106 5908
rect 11330 5896 11336 5908
rect 10100 5868 11336 5896
rect 10100 5856 10106 5868
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 11882 5896 11888 5908
rect 11795 5868 11888 5896
rect 11882 5856 11888 5868
rect 11940 5896 11946 5908
rect 12526 5896 12532 5908
rect 11940 5868 12532 5896
rect 11940 5856 11946 5868
rect 12526 5856 12532 5868
rect 12584 5856 12590 5908
rect 12710 5896 12716 5908
rect 12671 5868 12716 5896
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 12894 5856 12900 5908
rect 12952 5896 12958 5908
rect 14369 5899 14427 5905
rect 14369 5896 14381 5899
rect 12952 5868 14381 5896
rect 12952 5856 12958 5868
rect 14369 5865 14381 5868
rect 14415 5865 14427 5899
rect 14369 5859 14427 5865
rect 9766 5828 9772 5840
rect 9048 5800 9772 5828
rect 9766 5788 9772 5800
rect 9824 5788 9830 5840
rect 9876 5800 10732 5828
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5729 1455 5763
rect 2130 5760 2136 5772
rect 2091 5732 2136 5760
rect 1397 5723 1455 5729
rect 2130 5720 2136 5732
rect 2188 5720 2194 5772
rect 2400 5763 2458 5769
rect 2400 5729 2412 5763
rect 2446 5760 2458 5763
rect 4614 5760 4620 5772
rect 2446 5732 4620 5760
rect 2446 5729 2458 5732
rect 2400 5723 2458 5729
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 6730 5760 6736 5772
rect 5460 5732 6736 5760
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5692 4951 5695
rect 5166 5692 5172 5704
rect 4939 5664 5172 5692
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 5460 5701 5488 5732
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 7541 5763 7599 5769
rect 7541 5760 7553 5763
rect 7248 5732 7553 5760
rect 7248 5720 7254 5732
rect 7541 5729 7553 5732
rect 7587 5729 7599 5763
rect 7541 5723 7599 5729
rect 8846 5720 8852 5772
rect 8904 5760 8910 5772
rect 9309 5763 9367 5769
rect 9309 5760 9321 5763
rect 8904 5732 9321 5760
rect 8904 5720 8910 5732
rect 9309 5729 9321 5732
rect 9355 5729 9367 5763
rect 9876 5760 9904 5800
rect 9309 5723 9367 5729
rect 9416 5732 9904 5760
rect 9944 5763 10002 5769
rect 5445 5695 5503 5701
rect 5445 5661 5457 5695
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 6822 5652 6828 5704
rect 6880 5692 6886 5704
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 6880 5664 7297 5692
rect 6880 5652 6886 5664
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 3878 5584 3884 5636
rect 3936 5624 3942 5636
rect 5074 5624 5080 5636
rect 3936 5596 5080 5624
rect 3936 5584 3942 5596
rect 5074 5584 5080 5596
rect 5132 5584 5138 5636
rect 8294 5584 8300 5636
rect 8352 5624 8358 5636
rect 8665 5627 8723 5633
rect 8665 5624 8677 5627
rect 8352 5596 8677 5624
rect 8352 5584 8358 5596
rect 8665 5593 8677 5596
rect 8711 5593 8723 5627
rect 8665 5587 8723 5593
rect 8846 5584 8852 5636
rect 8904 5624 8910 5636
rect 9125 5627 9183 5633
rect 9125 5624 9137 5627
rect 8904 5596 9137 5624
rect 8904 5584 8910 5596
rect 9125 5593 9137 5596
rect 9171 5624 9183 5627
rect 9306 5624 9312 5636
rect 9171 5596 9312 5624
rect 9171 5593 9183 5596
rect 9125 5587 9183 5593
rect 9306 5584 9312 5596
rect 9364 5584 9370 5636
rect 1394 5516 1400 5568
rect 1452 5556 1458 5568
rect 1581 5559 1639 5565
rect 1581 5556 1593 5559
rect 1452 5528 1593 5556
rect 1452 5516 1458 5528
rect 1581 5525 1593 5528
rect 1627 5525 1639 5559
rect 1581 5519 1639 5525
rect 1854 5516 1860 5568
rect 1912 5556 1918 5568
rect 2406 5556 2412 5568
rect 1912 5528 2412 5556
rect 1912 5516 1918 5528
rect 2406 5516 2412 5528
rect 2464 5556 2470 5568
rect 3513 5559 3571 5565
rect 3513 5556 3525 5559
rect 2464 5528 3525 5556
rect 2464 5516 2470 5528
rect 3513 5525 3525 5528
rect 3559 5525 3571 5559
rect 3513 5519 3571 5525
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 4249 5559 4307 5565
rect 4249 5556 4261 5559
rect 4120 5528 4261 5556
rect 4120 5516 4126 5528
rect 4249 5525 4261 5528
rect 4295 5525 4307 5559
rect 4249 5519 4307 5525
rect 5442 5516 5448 5568
rect 5500 5556 5506 5568
rect 6825 5559 6883 5565
rect 6825 5556 6837 5559
rect 5500 5528 6837 5556
rect 5500 5516 5506 5528
rect 6825 5525 6837 5528
rect 6871 5525 6883 5559
rect 6825 5519 6883 5525
rect 7558 5516 7564 5568
rect 7616 5556 7622 5568
rect 9416 5556 9444 5732
rect 9944 5729 9956 5763
rect 9990 5760 10002 5763
rect 10502 5760 10508 5772
rect 9990 5732 10508 5760
rect 9990 5729 10002 5732
rect 9944 5723 10002 5729
rect 10502 5720 10508 5732
rect 10560 5720 10566 5772
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 10704 5692 10732 5800
rect 11054 5788 11060 5840
rect 11112 5828 11118 5840
rect 12158 5828 12164 5840
rect 11112 5800 12164 5828
rect 11112 5788 11118 5800
rect 12158 5788 12164 5800
rect 12216 5788 12222 5840
rect 10778 5720 10784 5772
rect 10836 5760 10842 5772
rect 11606 5760 11612 5772
rect 10836 5732 11612 5760
rect 10836 5720 10842 5732
rect 11606 5720 11612 5732
rect 11664 5760 11670 5772
rect 11977 5763 12035 5769
rect 11977 5760 11989 5763
rect 11664 5732 11989 5760
rect 11664 5720 11670 5732
rect 11977 5729 11989 5732
rect 12023 5729 12035 5763
rect 11977 5723 12035 5729
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 13081 5763 13139 5769
rect 13081 5760 13093 5763
rect 12492 5732 13093 5760
rect 12492 5720 12498 5732
rect 13081 5729 13093 5732
rect 13127 5729 13139 5763
rect 13081 5723 13139 5729
rect 13173 5763 13231 5769
rect 13173 5729 13185 5763
rect 13219 5760 13231 5763
rect 13906 5760 13912 5772
rect 13219 5732 13912 5760
rect 13219 5729 13231 5732
rect 13173 5723 13231 5729
rect 13906 5720 13912 5732
rect 13964 5720 13970 5772
rect 14277 5763 14335 5769
rect 14277 5729 14289 5763
rect 14323 5760 14335 5763
rect 15102 5760 15108 5772
rect 14323 5732 15108 5760
rect 14323 5729 14335 5732
rect 14277 5723 14335 5729
rect 12158 5692 12164 5704
rect 10704 5664 11192 5692
rect 12119 5664 12164 5692
rect 9677 5655 9735 5661
rect 7616 5528 9444 5556
rect 9692 5556 9720 5655
rect 11054 5624 11060 5636
rect 11015 5596 11060 5624
rect 11054 5584 11060 5596
rect 11112 5584 11118 5636
rect 11164 5624 11192 5664
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 12986 5652 12992 5704
rect 13044 5692 13050 5704
rect 13265 5695 13323 5701
rect 13265 5692 13277 5695
rect 13044 5664 13277 5692
rect 13044 5652 13050 5664
rect 13265 5661 13277 5664
rect 13311 5661 13323 5695
rect 13265 5655 13323 5661
rect 13354 5652 13360 5704
rect 13412 5692 13418 5704
rect 14292 5692 14320 5723
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 14458 5692 14464 5704
rect 13412 5664 14320 5692
rect 14419 5664 14464 5692
rect 13412 5652 13418 5664
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 14182 5624 14188 5636
rect 11164 5596 14188 5624
rect 14182 5584 14188 5596
rect 14240 5584 14246 5636
rect 10410 5556 10416 5568
rect 9692 5528 10416 5556
rect 7616 5516 7622 5528
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 11517 5559 11575 5565
rect 11517 5556 11529 5559
rect 11204 5528 11529 5556
rect 11204 5516 11210 5528
rect 11517 5525 11529 5528
rect 11563 5525 11575 5559
rect 13906 5556 13912 5568
rect 13867 5528 13912 5556
rect 11517 5519 11575 5525
rect 13906 5516 13912 5528
rect 13964 5516 13970 5568
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 1857 5355 1915 5361
rect 1857 5321 1869 5355
rect 1903 5352 1915 5355
rect 3234 5352 3240 5364
rect 1903 5324 3240 5352
rect 1903 5321 1915 5324
rect 1857 5315 1915 5321
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 4338 5312 4344 5364
rect 4396 5352 4402 5364
rect 4396 5324 7788 5352
rect 4396 5312 4402 5324
rect 3050 5284 3056 5296
rect 2240 5256 3056 5284
rect 2240 5157 2268 5256
rect 3050 5244 3056 5256
rect 3108 5244 3114 5296
rect 4433 5287 4491 5293
rect 4433 5253 4445 5287
rect 4479 5284 4491 5287
rect 4614 5284 4620 5296
rect 4479 5256 4620 5284
rect 4479 5253 4491 5256
rect 4433 5247 4491 5253
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 6638 5244 6644 5296
rect 6696 5284 6702 5296
rect 6822 5284 6828 5296
rect 6696 5256 6828 5284
rect 6696 5244 6702 5256
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 7760 5284 7788 5324
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 8168 5324 8217 5352
rect 8168 5312 8174 5324
rect 8205 5321 8217 5324
rect 8251 5352 8263 5355
rect 10226 5352 10232 5364
rect 8251 5324 10232 5352
rect 8251 5321 8263 5324
rect 8205 5315 8263 5321
rect 10226 5312 10232 5324
rect 10284 5352 10290 5364
rect 11054 5352 11060 5364
rect 10284 5324 11060 5352
rect 10284 5312 10290 5324
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11514 5312 11520 5364
rect 11572 5352 11578 5364
rect 11882 5352 11888 5364
rect 11572 5324 11888 5352
rect 11572 5312 11578 5324
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 12342 5312 12348 5364
rect 12400 5352 12406 5364
rect 12437 5355 12495 5361
rect 12437 5352 12449 5355
rect 12400 5324 12449 5352
rect 12400 5312 12406 5324
rect 12437 5321 12449 5324
rect 12483 5321 12495 5355
rect 13630 5352 13636 5364
rect 13591 5324 13636 5352
rect 12437 5315 12495 5321
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 8662 5284 8668 5296
rect 7760 5256 8668 5284
rect 8662 5244 8668 5256
rect 8720 5244 8726 5296
rect 10045 5287 10103 5293
rect 10045 5253 10057 5287
rect 10091 5284 10103 5287
rect 11422 5284 11428 5296
rect 10091 5256 11428 5284
rect 10091 5253 10103 5256
rect 10045 5247 10103 5253
rect 11422 5244 11428 5256
rect 11480 5244 11486 5296
rect 12618 5244 12624 5296
rect 12676 5284 12682 5296
rect 15013 5287 15071 5293
rect 15013 5284 15025 5287
rect 12676 5256 15025 5284
rect 12676 5244 12682 5256
rect 15013 5253 15025 5256
rect 15059 5253 15071 5287
rect 15013 5247 15071 5253
rect 2498 5216 2504 5228
rect 2411 5188 2504 5216
rect 2498 5176 2504 5188
rect 2556 5216 2562 5228
rect 2556 5188 3004 5216
rect 2556 5176 2562 5188
rect 2225 5151 2283 5157
rect 2225 5117 2237 5151
rect 2271 5117 2283 5151
rect 2225 5111 2283 5117
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2976 5012 3004 5188
rect 9950 5176 9956 5228
rect 10008 5176 10014 5228
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 11054 5216 11060 5228
rect 10560 5188 10732 5216
rect 11015 5188 11060 5216
rect 10560 5176 10566 5188
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 4890 5148 4896 5160
rect 3099 5120 4896 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 5160 5151 5218 5157
rect 5160 5117 5172 5151
rect 5206 5148 5218 5151
rect 5442 5148 5448 5160
rect 5206 5120 5448 5148
rect 5206 5117 5218 5120
rect 5160 5111 5218 5117
rect 3320 5083 3378 5089
rect 3320 5049 3332 5083
rect 3366 5080 3378 5083
rect 3418 5080 3424 5092
rect 3366 5052 3424 5080
rect 3366 5049 3378 5052
rect 3320 5043 3378 5049
rect 3418 5040 3424 5052
rect 3476 5040 3482 5092
rect 5175 5080 5203 5111
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6788 5120 6837 5148
rect 6788 5108 6794 5120
rect 6825 5117 6837 5120
rect 6871 5148 6883 5151
rect 6914 5148 6920 5160
rect 6871 5120 6920 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7098 5157 7104 5160
rect 7092 5111 7104 5157
rect 7156 5148 7162 5160
rect 7156 5120 7192 5148
rect 7098 5108 7104 5111
rect 7156 5108 7162 5120
rect 7650 5108 7656 5160
rect 7708 5148 7714 5160
rect 8938 5157 8944 5160
rect 8665 5151 8723 5157
rect 8665 5148 8677 5151
rect 7708 5120 8677 5148
rect 7708 5108 7714 5120
rect 8665 5117 8677 5120
rect 8711 5117 8723 5151
rect 8932 5148 8944 5157
rect 8899 5120 8944 5148
rect 8665 5111 8723 5117
rect 8932 5111 8944 5120
rect 8938 5108 8944 5111
rect 8996 5108 9002 5160
rect 9968 5148 9996 5176
rect 10594 5148 10600 5160
rect 9968 5120 10600 5148
rect 10594 5108 10600 5120
rect 10652 5108 10658 5160
rect 10704 5148 10732 5188
rect 11054 5176 11060 5188
rect 11112 5216 11118 5228
rect 12158 5216 12164 5228
rect 11112 5188 12164 5216
rect 11112 5176 11118 5188
rect 11624 5160 11652 5188
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 12986 5216 12992 5228
rect 12947 5188 12992 5216
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 13446 5216 13452 5228
rect 13407 5188 13452 5216
rect 13446 5176 13452 5188
rect 13504 5216 13510 5228
rect 14182 5216 14188 5228
rect 13504 5188 14044 5216
rect 14143 5188 14188 5216
rect 13504 5176 13510 5188
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10704 5120 10885 5148
rect 10873 5117 10885 5120
rect 10919 5148 10931 5151
rect 11238 5148 11244 5160
rect 10919 5120 11244 5148
rect 10919 5117 10931 5120
rect 10873 5111 10931 5117
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 11606 5108 11612 5160
rect 11664 5108 11670 5160
rect 11701 5151 11759 5157
rect 11701 5117 11713 5151
rect 11747 5148 11759 5151
rect 13814 5148 13820 5160
rect 11747 5120 13820 5148
rect 11747 5117 11759 5120
rect 11701 5111 11759 5117
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14016 5157 14044 5188
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5117 14059 5151
rect 14001 5111 14059 5117
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5148 14887 5151
rect 14918 5148 14924 5160
rect 14875 5120 14924 5148
rect 14875 5117 14887 5120
rect 14829 5111 14887 5117
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 3528 5052 5203 5080
rect 3528 5012 3556 5052
rect 5626 5040 5632 5092
rect 5684 5080 5690 5092
rect 5684 5052 6960 5080
rect 5684 5040 5690 5052
rect 6932 5024 6960 5052
rect 8110 5040 8116 5092
rect 8168 5080 8174 5092
rect 9122 5080 9128 5092
rect 8168 5052 9128 5080
rect 8168 5040 8174 5052
rect 9122 5040 9128 5052
rect 9180 5040 9186 5092
rect 9490 5040 9496 5092
rect 9548 5080 9554 5092
rect 10962 5080 10968 5092
rect 9548 5052 10640 5080
rect 10923 5052 10968 5080
rect 9548 5040 9554 5052
rect 6270 5012 6276 5024
rect 2372 4984 2417 5012
rect 2976 4984 3556 5012
rect 6231 4984 6276 5012
rect 2372 4972 2378 4984
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6914 4972 6920 5024
rect 6972 4972 6978 5024
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 9214 5012 9220 5024
rect 8628 4984 9220 5012
rect 8628 4972 8634 4984
rect 9214 4972 9220 4984
rect 9272 4972 9278 5024
rect 9306 4972 9312 5024
rect 9364 5012 9370 5024
rect 10042 5012 10048 5024
rect 9364 4984 10048 5012
rect 9364 4972 9370 4984
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 10134 4972 10140 5024
rect 10192 5012 10198 5024
rect 10505 5015 10563 5021
rect 10505 5012 10517 5015
rect 10192 4984 10517 5012
rect 10192 4972 10198 4984
rect 10505 4981 10517 4984
rect 10551 4981 10563 5015
rect 10612 5012 10640 5052
rect 10962 5040 10968 5052
rect 11020 5040 11026 5092
rect 11790 5040 11796 5092
rect 11848 5080 11854 5092
rect 12805 5083 12863 5089
rect 12805 5080 12817 5083
rect 11848 5052 12817 5080
rect 11848 5040 11854 5052
rect 12805 5049 12817 5052
rect 12851 5080 12863 5083
rect 13262 5080 13268 5092
rect 12851 5052 13268 5080
rect 12851 5049 12863 5052
rect 12805 5043 12863 5049
rect 13262 5040 13268 5052
rect 13320 5040 13326 5092
rect 13630 5040 13636 5092
rect 13688 5080 13694 5092
rect 14093 5083 14151 5089
rect 14093 5080 14105 5083
rect 13688 5052 14105 5080
rect 13688 5040 13694 5052
rect 14093 5049 14105 5052
rect 14139 5049 14151 5083
rect 14093 5043 14151 5049
rect 12434 5012 12440 5024
rect 10612 4984 12440 5012
rect 10505 4975 10563 4981
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 12897 5015 12955 5021
rect 12897 4981 12909 5015
rect 12943 5012 12955 5015
rect 13814 5012 13820 5024
rect 12943 4984 13820 5012
rect 12943 4981 12955 4984
rect 12897 4975 12955 4981
rect 13814 4972 13820 4984
rect 13872 5012 13878 5024
rect 14642 5012 14648 5024
rect 13872 4984 14648 5012
rect 13872 4972 13878 4984
rect 14642 4972 14648 4984
rect 14700 4972 14706 5024
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 3050 4768 3056 4820
rect 3108 4808 3114 4820
rect 10042 4808 10048 4820
rect 3108 4780 9720 4808
rect 10003 4780 10048 4808
rect 3108 4768 3114 4780
rect 2406 4749 2412 4752
rect 2400 4740 2412 4749
rect 2367 4712 2412 4740
rect 2400 4703 2412 4712
rect 2406 4700 2412 4703
rect 2464 4700 2470 4752
rect 2682 4700 2688 4752
rect 2740 4740 2746 4752
rect 4338 4740 4344 4752
rect 2740 4712 4344 4740
rect 2740 4700 2746 4712
rect 4338 4700 4344 4712
rect 4396 4700 4402 4752
rect 4525 4743 4583 4749
rect 4525 4709 4537 4743
rect 4571 4740 4583 4743
rect 6822 4740 6828 4752
rect 4571 4712 6828 4740
rect 4571 4709 4583 4712
rect 4525 4703 4583 4709
rect 6822 4700 6828 4712
rect 6880 4700 6886 4752
rect 7006 4700 7012 4752
rect 7064 4740 7070 4752
rect 7650 4740 7656 4752
rect 7064 4712 7656 4740
rect 7064 4700 7070 4712
rect 7650 4700 7656 4712
rect 7708 4700 7714 4752
rect 7742 4700 7748 4752
rect 7800 4740 7806 4752
rect 8846 4740 8852 4752
rect 7800 4712 8852 4740
rect 7800 4700 7806 4712
rect 8846 4700 8852 4712
rect 8904 4700 8910 4752
rect 8941 4743 8999 4749
rect 8941 4709 8953 4743
rect 8987 4740 8999 4743
rect 9398 4740 9404 4752
rect 8987 4712 9404 4740
rect 8987 4709 8999 4712
rect 8941 4703 8999 4709
rect 9398 4700 9404 4712
rect 9456 4700 9462 4752
rect 9582 4740 9588 4752
rect 9508 4712 9588 4740
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1854 4672 1860 4684
rect 1443 4644 1860 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1854 4632 1860 4644
rect 1912 4632 1918 4684
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4672 2191 4675
rect 2866 4672 2872 4684
rect 2179 4644 2872 4672
rect 2179 4641 2191 4644
rect 2133 4635 2191 4641
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 2958 4632 2964 4684
rect 3016 4672 3022 4684
rect 3786 4672 3792 4684
rect 3016 4644 3792 4672
rect 3016 4632 3022 4644
rect 3786 4632 3792 4644
rect 3844 4632 3850 4684
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 5350 4672 5356 4684
rect 4479 4644 5356 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 5534 4681 5540 4684
rect 5528 4672 5540 4681
rect 5495 4644 5540 4672
rect 5528 4635 5540 4644
rect 5534 4632 5540 4635
rect 5592 4632 5598 4684
rect 7374 4681 7380 4684
rect 7368 4672 7380 4681
rect 7335 4644 7380 4672
rect 7368 4635 7380 4644
rect 7374 4632 7380 4635
rect 7432 4632 7438 4684
rect 8202 4632 8208 4684
rect 8260 4672 8266 4684
rect 9508 4672 9536 4712
rect 9582 4700 9588 4712
rect 9640 4700 9646 4752
rect 9692 4740 9720 4780
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 10137 4811 10195 4817
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 11238 4808 11244 4820
rect 10183 4780 11244 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 11072 4752 11100 4780
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 11330 4768 11336 4820
rect 11388 4808 11394 4820
rect 12529 4811 12587 4817
rect 12529 4808 12541 4811
rect 11388 4780 12541 4808
rect 11388 4768 11394 4780
rect 12529 4777 12541 4780
rect 12575 4808 12587 4811
rect 12575 4780 13124 4808
rect 12575 4777 12587 4780
rect 12529 4771 12587 4777
rect 9950 4740 9956 4752
rect 9692 4712 9956 4740
rect 9950 4700 9956 4712
rect 10008 4700 10014 4752
rect 11054 4700 11060 4752
rect 11112 4700 11118 4752
rect 11882 4700 11888 4752
rect 11940 4740 11946 4752
rect 12434 4740 12440 4752
rect 11940 4712 12440 4740
rect 11940 4700 11946 4712
rect 12434 4700 12440 4712
rect 12492 4700 12498 4752
rect 12710 4700 12716 4752
rect 12768 4740 12774 4752
rect 13096 4740 13124 4780
rect 13170 4768 13176 4820
rect 13228 4808 13234 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 13228 4780 13277 4808
rect 13228 4768 13234 4780
rect 13265 4777 13277 4780
rect 13311 4777 13323 4811
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 13265 4771 13323 4777
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 12768 4712 12848 4740
rect 13096 4712 14504 4740
rect 12768 4700 12774 4712
rect 10962 4672 10968 4684
rect 8260 4644 9536 4672
rect 9784 4644 10968 4672
rect 8260 4632 8266 4644
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 3513 4539 3571 4545
rect 3513 4505 3525 4539
rect 3559 4536 3571 4539
rect 4614 4536 4620 4548
rect 3559 4508 4620 4536
rect 3559 4505 3571 4508
rect 3513 4499 3571 4505
rect 4614 4496 4620 4508
rect 4672 4496 4678 4548
rect 1581 4471 1639 4477
rect 1581 4437 1593 4471
rect 1627 4468 1639 4471
rect 2406 4468 2412 4480
rect 1627 4440 2412 4468
rect 1627 4437 1639 4440
rect 1581 4431 1639 4437
rect 2406 4428 2412 4440
rect 2464 4428 2470 4480
rect 4065 4471 4123 4477
rect 4065 4437 4077 4471
rect 4111 4468 4123 4471
rect 4338 4468 4344 4480
rect 4111 4440 4344 4468
rect 4111 4437 4123 4440
rect 4065 4431 4123 4437
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 4724 4468 4752 4567
rect 5074 4564 5080 4616
rect 5132 4604 5138 4616
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 5132 4576 5273 4604
rect 5132 4564 5138 4576
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 7101 4607 7159 4613
rect 7101 4604 7113 4607
rect 6788 4576 7113 4604
rect 6788 4564 6794 4576
rect 7101 4573 7113 4576
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 8846 4564 8852 4616
rect 8904 4604 8910 4616
rect 9784 4604 9812 4644
rect 10962 4632 10968 4644
rect 11020 4632 11026 4684
rect 11238 4672 11244 4684
rect 11199 4644 11244 4672
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 11514 4632 11520 4684
rect 11572 4672 11578 4684
rect 11790 4672 11796 4684
rect 11572 4644 11796 4672
rect 11572 4632 11578 4644
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 8904 4576 9812 4604
rect 8904 4564 8910 4576
rect 9858 4564 9864 4616
rect 9916 4604 9922 4616
rect 10042 4604 10048 4616
rect 9916 4576 10048 4604
rect 9916 4564 9922 4576
rect 10042 4564 10048 4576
rect 10100 4604 10106 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 10100 4576 10241 4604
rect 10100 4564 10106 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 10778 4564 10784 4616
rect 10836 4604 10842 4616
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 10836 4576 11345 4604
rect 10836 4564 10842 4576
rect 11333 4573 11345 4576
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4604 11483 4607
rect 11606 4604 11612 4616
rect 11471 4576 11612 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 11698 4564 11704 4616
rect 11756 4604 11762 4616
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 11756 4576 12633 4604
rect 11756 4564 11762 4576
rect 12621 4573 12633 4576
rect 12667 4573 12679 4607
rect 12820 4604 12848 4712
rect 14476 4681 14504 4712
rect 13725 4675 13783 4681
rect 13725 4672 13737 4675
rect 13648 4644 13737 4672
rect 13648 4604 13676 4644
rect 13725 4641 13737 4644
rect 13771 4641 13783 4675
rect 13725 4635 13783 4641
rect 14461 4675 14519 4681
rect 14461 4641 14473 4675
rect 14507 4641 14519 4675
rect 14461 4635 14519 4641
rect 12820 4576 13676 4604
rect 13817 4607 13875 4613
rect 12621 4567 12679 4573
rect 13817 4573 13829 4607
rect 13863 4604 13875 4607
rect 14182 4604 14188 4616
rect 13863 4576 14188 4604
rect 13863 4573 13875 4576
rect 13817 4567 13875 4573
rect 8294 4496 8300 4548
rect 8352 4496 8358 4548
rect 8478 4536 8484 4548
rect 8439 4508 8484 4536
rect 8478 4496 8484 4508
rect 8536 4496 8542 4548
rect 8662 4496 8668 4548
rect 8720 4536 8726 4548
rect 12069 4539 12127 4545
rect 12069 4536 12081 4539
rect 8720 4508 12081 4536
rect 8720 4496 8726 4508
rect 12069 4505 12081 4508
rect 12115 4505 12127 4539
rect 12069 4499 12127 4505
rect 12986 4496 12992 4548
rect 13044 4536 13050 4548
rect 13832 4536 13860 4567
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14642 4536 14648 4548
rect 13044 4508 13860 4536
rect 14603 4508 14648 4536
rect 13044 4496 13050 4508
rect 14642 4496 14648 4508
rect 14700 4496 14706 4548
rect 5074 4468 5080 4480
rect 4724 4440 5080 4468
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 6641 4471 6699 4477
rect 6641 4437 6653 4471
rect 6687 4468 6699 4471
rect 7374 4468 7380 4480
rect 6687 4440 7380 4468
rect 6687 4437 6699 4440
rect 6641 4431 6699 4437
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 8312 4468 8340 4496
rect 9674 4468 9680 4480
rect 7524 4440 8340 4468
rect 9635 4440 9680 4468
rect 7524 4428 7530 4440
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 10318 4428 10324 4480
rect 10376 4468 10382 4480
rect 10873 4471 10931 4477
rect 10873 4468 10885 4471
rect 10376 4440 10885 4468
rect 10376 4428 10382 4440
rect 10873 4437 10885 4440
rect 10919 4437 10931 4471
rect 10873 4431 10931 4437
rect 10962 4428 10968 4480
rect 11020 4468 11026 4480
rect 11882 4468 11888 4480
rect 11020 4440 11888 4468
rect 11020 4428 11026 4440
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 2866 4224 2872 4276
rect 2924 4264 2930 4276
rect 4890 4264 4896 4276
rect 2924 4236 4896 4264
rect 2924 4224 2930 4236
rect 2498 4128 2504 4140
rect 2459 4100 2504 4128
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 3068 4137 3096 4236
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 5074 4224 5080 4276
rect 5132 4264 5138 4276
rect 7006 4264 7012 4276
rect 5132 4236 7012 4264
rect 5132 4224 5138 4236
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 7156 4236 7788 4264
rect 7156 4224 7162 4236
rect 4246 4156 4252 4208
rect 4304 4196 4310 4208
rect 4433 4199 4491 4205
rect 4433 4196 4445 4199
rect 4304 4168 4445 4196
rect 4304 4156 4310 4168
rect 4433 4165 4445 4168
rect 4479 4196 4491 4199
rect 4614 4196 4620 4208
rect 4479 4168 4620 4196
rect 4479 4165 4491 4168
rect 4433 4159 4491 4165
rect 4614 4156 4620 4168
rect 4672 4156 4678 4208
rect 7760 4196 7788 4236
rect 7834 4224 7840 4276
rect 7892 4264 7898 4276
rect 9214 4264 9220 4276
rect 7892 4236 9220 4264
rect 7892 4224 7898 4236
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 9306 4224 9312 4276
rect 9364 4264 9370 4276
rect 10226 4264 10232 4276
rect 9364 4236 10232 4264
rect 9364 4224 9370 4236
rect 10226 4224 10232 4236
rect 10284 4224 10290 4276
rect 11057 4267 11115 4273
rect 11057 4233 11069 4267
rect 11103 4264 11115 4267
rect 11238 4264 11244 4276
rect 11103 4236 11244 4264
rect 11103 4233 11115 4236
rect 11057 4227 11115 4233
rect 11238 4224 11244 4236
rect 11296 4224 11302 4276
rect 11422 4224 11428 4276
rect 11480 4264 11486 4276
rect 11480 4236 12112 4264
rect 11480 4224 11486 4236
rect 7760 4168 7860 4196
rect 3053 4131 3111 4137
rect 3053 4097 3065 4131
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 7832 4128 7860 4168
rect 8110 4156 8116 4208
rect 8168 4196 8174 4208
rect 8570 4196 8576 4208
rect 8168 4168 8576 4196
rect 8168 4156 8174 4168
rect 8570 4156 8576 4168
rect 8628 4156 8634 4208
rect 8665 4199 8723 4205
rect 8665 4165 8677 4199
rect 8711 4196 8723 4199
rect 8711 4168 9720 4196
rect 8711 4165 8723 4168
rect 8665 4159 8723 4165
rect 9306 4128 9312 4140
rect 4212 4100 5028 4128
rect 4212 4088 4218 4100
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4060 2283 4063
rect 4890 4060 4896 4072
rect 2271 4032 4752 4060
rect 4851 4032 4896 4060
rect 2271 4029 2283 4032
rect 2225 4023 2283 4029
rect 3320 3995 3378 4001
rect 3320 3961 3332 3995
rect 3366 3992 3378 3995
rect 4246 3992 4252 4004
rect 3366 3964 4252 3992
rect 3366 3961 3378 3964
rect 3320 3955 3378 3961
rect 4246 3952 4252 3964
rect 4304 3952 4310 4004
rect 1857 3927 1915 3933
rect 1857 3893 1869 3927
rect 1903 3924 1915 3927
rect 2130 3924 2136 3936
rect 1903 3896 2136 3924
rect 1903 3893 1915 3896
rect 1857 3887 1915 3893
rect 2130 3884 2136 3896
rect 2188 3884 2194 3936
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 4154 3924 4160 3936
rect 2363 3896 4160 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 4724 3924 4752 4032
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 5000 4060 5028 4100
rect 6003 4100 6960 4128
rect 7832 4100 9312 4128
rect 6003 4060 6031 4100
rect 5000 4032 6031 4060
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6788 4032 6837 4060
rect 6788 4020 6794 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6932 4060 6960 4100
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 8662 4060 8668 4072
rect 6932 4032 8668 4060
rect 6825 4023 6883 4029
rect 5166 4001 5172 4004
rect 5160 3992 5172 4001
rect 5079 3964 5172 3992
rect 5160 3955 5172 3964
rect 5224 3992 5230 4004
rect 6840 3992 6868 4023
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 9692 4060 9720 4168
rect 9766 4156 9772 4208
rect 9824 4196 9830 4208
rect 9861 4199 9919 4205
rect 9861 4196 9873 4199
rect 9824 4168 9873 4196
rect 9824 4156 9830 4168
rect 9861 4165 9873 4168
rect 9907 4165 9919 4199
rect 10244 4196 10272 4224
rect 12084 4196 12112 4236
rect 12158 4224 12164 4276
rect 12216 4264 12222 4276
rect 13630 4264 13636 4276
rect 12216 4236 13636 4264
rect 12216 4224 12222 4236
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 14458 4196 14464 4208
rect 10244 4168 11652 4196
rect 12084 4168 14464 4196
rect 9861 4159 9919 4165
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10413 4131 10471 4137
rect 10413 4128 10425 4131
rect 10100 4100 10425 4128
rect 10100 4088 10106 4100
rect 10413 4097 10425 4100
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 11330 4088 11336 4140
rect 11388 4128 11394 4140
rect 11624 4137 11652 4168
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 11388 4100 11529 4128
rect 11388 4088 11394 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 11609 4131 11667 4137
rect 11609 4097 11621 4131
rect 11655 4097 11667 4131
rect 11609 4091 11667 4097
rect 11882 4088 11888 4140
rect 11940 4128 11946 4140
rect 12986 4128 12992 4140
rect 11940 4100 12992 4128
rect 11940 4088 11946 4100
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 13078 4088 13084 4140
rect 13136 4128 13142 4140
rect 14200 4137 14228 4168
rect 14458 4156 14464 4168
rect 14516 4156 14522 4208
rect 14093 4131 14151 4137
rect 14093 4128 14105 4131
rect 13136 4100 14105 4128
rect 13136 4088 13142 4100
rect 14093 4097 14105 4100
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 14185 4131 14243 4137
rect 14185 4097 14197 4131
rect 14231 4097 14243 4131
rect 14185 4091 14243 4097
rect 10226 4060 10232 4072
rect 9692 4032 9996 4060
rect 10187 4032 10232 4060
rect 6914 3992 6920 4004
rect 5224 3964 6408 3992
rect 6840 3964 6920 3992
rect 5166 3952 5172 3955
rect 5224 3952 5230 3964
rect 5442 3924 5448 3936
rect 4724 3896 5448 3924
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 5534 3884 5540 3936
rect 5592 3924 5598 3936
rect 6273 3927 6331 3933
rect 6273 3924 6285 3927
rect 5592 3896 6285 3924
rect 5592 3884 5598 3896
rect 6273 3893 6285 3896
rect 6319 3893 6331 3927
rect 6380 3924 6408 3964
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 7006 3952 7012 4004
rect 7064 4001 7070 4004
rect 7064 3995 7128 4001
rect 7064 3961 7082 3995
rect 7116 3992 7128 3995
rect 7466 3992 7472 4004
rect 7116 3964 7472 3992
rect 7116 3961 7128 3964
rect 7064 3955 7128 3961
rect 7064 3952 7070 3955
rect 7466 3952 7472 3964
rect 7524 3992 7530 4004
rect 8110 3992 8116 4004
rect 7524 3964 8116 3992
rect 7524 3952 7530 3964
rect 8110 3952 8116 3964
rect 8168 3952 8174 4004
rect 8478 3952 8484 4004
rect 8536 3992 8542 4004
rect 9674 3992 9680 4004
rect 8536 3964 9680 3992
rect 8536 3952 8542 3964
rect 9674 3952 9680 3964
rect 9732 3952 9738 4004
rect 9968 3992 9996 4032
rect 10226 4020 10232 4032
rect 10284 4020 10290 4072
rect 10321 4063 10379 4069
rect 10321 4029 10333 4063
rect 10367 4060 10379 4063
rect 10686 4060 10692 4072
rect 10367 4032 10692 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 12434 4060 12440 4072
rect 11624 4032 12440 4060
rect 11624 4004 11652 4032
rect 12434 4020 12440 4032
rect 12492 4060 12498 4072
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12492 4032 12817 4060
rect 12492 4020 12498 4032
rect 12805 4029 12817 4032
rect 12851 4029 12863 4063
rect 12805 4023 12863 4029
rect 12897 4063 12955 4069
rect 12897 4029 12909 4063
rect 12943 4060 12955 4063
rect 13262 4060 13268 4072
rect 12943 4032 13268 4060
rect 12943 4029 12955 4032
rect 12897 4023 12955 4029
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 14829 4063 14887 4069
rect 14829 4029 14841 4063
rect 14875 4060 14887 4063
rect 15194 4060 15200 4072
rect 14875 4032 15200 4060
rect 14875 4029 14887 4032
rect 14829 4023 14887 4029
rect 15194 4020 15200 4032
rect 15252 4020 15258 4072
rect 10778 3992 10784 4004
rect 9968 3964 10784 3992
rect 10778 3952 10784 3964
rect 10836 3952 10842 4004
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 11112 3964 11468 3992
rect 11112 3952 11118 3964
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 6380 3896 8217 3924
rect 6273 3887 6331 3893
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 9030 3924 9036 3936
rect 8991 3896 9036 3924
rect 8205 3887 8263 3893
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 9125 3927 9183 3933
rect 9125 3893 9137 3927
rect 9171 3924 9183 3927
rect 9214 3924 9220 3936
rect 9171 3896 9220 3924
rect 9171 3893 9183 3896
rect 9125 3887 9183 3893
rect 9214 3884 9220 3896
rect 9272 3924 9278 3936
rect 9490 3924 9496 3936
rect 9272 3896 9496 3924
rect 9272 3884 9278 3896
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 11238 3924 11244 3936
rect 10100 3896 11244 3924
rect 10100 3884 10106 3896
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 11440 3933 11468 3964
rect 11606 3952 11612 4004
rect 11664 3952 11670 4004
rect 14001 3995 14059 4001
rect 14001 3961 14013 3995
rect 14047 3961 14059 3995
rect 14001 3955 14059 3961
rect 11425 3927 11483 3933
rect 11425 3893 11437 3927
rect 11471 3924 11483 3927
rect 11790 3924 11796 3936
rect 11471 3896 11796 3924
rect 11471 3893 11483 3896
rect 11425 3887 11483 3893
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12492 3896 12537 3924
rect 12492 3884 12498 3896
rect 13262 3884 13268 3936
rect 13320 3924 13326 3936
rect 13633 3927 13691 3933
rect 13633 3924 13645 3927
rect 13320 3896 13645 3924
rect 13320 3884 13326 3896
rect 13633 3893 13645 3896
rect 13679 3893 13691 3927
rect 14016 3924 14044 3955
rect 14458 3924 14464 3936
rect 14016 3896 14464 3924
rect 13633 3887 13691 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 14642 3884 14648 3936
rect 14700 3924 14706 3936
rect 15013 3927 15071 3933
rect 15013 3924 15025 3927
rect 14700 3896 15025 3924
rect 14700 3884 14706 3896
rect 15013 3893 15025 3896
rect 15059 3893 15071 3927
rect 15013 3887 15071 3893
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 1946 3720 1952 3732
rect 1907 3692 1952 3720
rect 1946 3680 1952 3692
rect 2004 3680 2010 3732
rect 2130 3680 2136 3732
rect 2188 3720 2194 3732
rect 3145 3723 3203 3729
rect 3145 3720 3157 3723
rect 2188 3692 3157 3720
rect 2188 3680 2194 3692
rect 3145 3689 3157 3692
rect 3191 3689 3203 3723
rect 3145 3683 3203 3689
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 3292 3692 3337 3720
rect 3292 3680 3298 3692
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 4430 3720 4436 3732
rect 4304 3692 4436 3720
rect 4304 3680 4310 3692
rect 4430 3680 4436 3692
rect 4488 3680 4494 3732
rect 4982 3720 4988 3732
rect 4943 3692 4988 3720
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 5500 3692 8616 3720
rect 5500 3680 5506 3692
rect 2041 3655 2099 3661
rect 2041 3621 2053 3655
rect 2087 3652 2099 3655
rect 2682 3652 2688 3664
rect 2087 3624 2688 3652
rect 2087 3621 2099 3624
rect 2041 3615 2099 3621
rect 2682 3612 2688 3624
rect 2740 3612 2746 3664
rect 4893 3655 4951 3661
rect 4893 3621 4905 3655
rect 4939 3652 4951 3655
rect 8478 3652 8484 3664
rect 4939 3624 8484 3652
rect 4939 3621 4951 3624
rect 4893 3615 4951 3621
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 8588 3652 8616 3692
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 8904 3692 8953 3720
rect 8904 3680 8910 3692
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 9674 3720 9680 3732
rect 8941 3683 8999 3689
rect 9048 3692 9680 3720
rect 9048 3652 9076 3692
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10873 3723 10931 3729
rect 10873 3720 10885 3723
rect 10008 3692 10885 3720
rect 10008 3680 10014 3692
rect 10873 3689 10885 3692
rect 10919 3689 10931 3723
rect 11238 3720 11244 3732
rect 11199 3692 11244 3720
rect 10873 3683 10931 3689
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 12066 3720 12072 3732
rect 12027 3692 12072 3720
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 12437 3723 12495 3729
rect 12437 3689 12449 3723
rect 12483 3720 12495 3723
rect 13262 3720 13268 3732
rect 12483 3692 13268 3720
rect 12483 3689 12495 3692
rect 12437 3683 12495 3689
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 13630 3720 13636 3732
rect 13591 3692 13636 3720
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 13906 3720 13912 3732
rect 13740 3692 13912 3720
rect 10045 3655 10103 3661
rect 10045 3652 10057 3655
rect 8588 3624 9076 3652
rect 9416 3624 10057 3652
rect 5988 3587 6046 3593
rect 5988 3584 6000 3587
rect 3436 3556 6000 3584
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 3234 3516 3240 3528
rect 2271 3488 3240 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 3436 3525 3464 3556
rect 5988 3553 6000 3556
rect 6034 3584 6046 3587
rect 6270 3584 6276 3596
rect 6034 3556 6276 3584
rect 6034 3553 6046 3556
rect 5988 3547 6046 3553
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 6914 3584 6920 3596
rect 6788 3556 6920 3584
rect 6788 3544 6794 3556
rect 6914 3544 6920 3556
rect 6972 3584 6978 3596
rect 7558 3584 7564 3596
rect 6972 3556 7564 3584
rect 6972 3544 6978 3556
rect 7558 3544 7564 3556
rect 7616 3544 7622 3596
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 7817 3587 7875 3593
rect 7817 3584 7829 3587
rect 7708 3556 7829 3584
rect 7708 3544 7714 3556
rect 7817 3553 7829 3556
rect 7863 3553 7875 3587
rect 7817 3547 7875 3553
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 9416 3584 9444 3624
rect 10045 3621 10057 3624
rect 10091 3652 10103 3655
rect 12529 3655 12587 3661
rect 10091 3624 10272 3652
rect 10091 3621 10103 3624
rect 10045 3615 10103 3621
rect 9180 3556 9444 3584
rect 9180 3544 9186 3556
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 10244 3584 10272 3624
rect 12529 3621 12541 3655
rect 12575 3652 12587 3655
rect 13740 3652 13768 3692
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 12575 3624 13768 3652
rect 12575 3621 12587 3624
rect 12529 3615 12587 3621
rect 13814 3612 13820 3664
rect 13872 3652 13878 3664
rect 14182 3652 14188 3664
rect 13872 3624 14188 3652
rect 13872 3612 13878 3624
rect 14182 3612 14188 3624
rect 14240 3612 14246 3664
rect 9548 3556 10088 3584
rect 10244 3556 10364 3584
rect 9548 3544 9554 3556
rect 10060 3528 10088 3556
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3485 3479 3519
rect 5166 3516 5172 3528
rect 5127 3488 5172 3516
rect 3421 3479 3479 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5500 3488 5733 3516
rect 5500 3476 5506 3488
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 8864 3488 9720 3516
rect 2774 3408 2780 3460
rect 2832 3448 2838 3460
rect 2832 3420 2877 3448
rect 2832 3408 2838 3420
rect 3142 3408 3148 3460
rect 3200 3448 3206 3460
rect 5626 3448 5632 3460
rect 3200 3420 5632 3448
rect 3200 3408 3206 3420
rect 5626 3408 5632 3420
rect 5684 3408 5690 3460
rect 6822 3408 6828 3460
rect 6880 3448 6886 3460
rect 6880 3420 7604 3448
rect 6880 3408 6886 3420
rect 750 3340 756 3392
rect 808 3380 814 3392
rect 1486 3380 1492 3392
rect 808 3352 1492 3380
rect 808 3340 814 3352
rect 1486 3340 1492 3352
rect 1544 3340 1550 3392
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 4525 3383 4583 3389
rect 4525 3380 4537 3383
rect 4212 3352 4537 3380
rect 4212 3340 4218 3352
rect 4525 3349 4537 3352
rect 4571 3349 4583 3383
rect 7098 3380 7104 3392
rect 7059 3352 7104 3380
rect 4525 3343 4583 3349
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 7576 3380 7604 3420
rect 8864 3380 8892 3488
rect 9692 3457 9720 3488
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10137 3519 10195 3525
rect 10137 3516 10149 3519
rect 10100 3488 10149 3516
rect 10100 3476 10106 3488
rect 10137 3485 10149 3488
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 10229 3519 10287 3525
rect 10229 3485 10241 3519
rect 10275 3485 10287 3519
rect 10336 3516 10364 3556
rect 10410 3544 10416 3596
rect 10468 3584 10474 3596
rect 11146 3584 11152 3596
rect 10468 3556 11152 3584
rect 10468 3544 10474 3556
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 11333 3587 11391 3593
rect 11333 3584 11345 3587
rect 11296 3556 11345 3584
rect 11296 3544 11302 3556
rect 11333 3553 11345 3556
rect 11379 3553 11391 3587
rect 11333 3547 11391 3553
rect 14090 3544 14096 3596
rect 14148 3584 14154 3596
rect 14461 3587 14519 3593
rect 14461 3584 14473 3587
rect 14148 3556 14473 3584
rect 14148 3544 14154 3556
rect 14461 3553 14473 3556
rect 14507 3553 14519 3587
rect 14461 3547 14519 3553
rect 10778 3516 10784 3528
rect 10336 3488 10784 3516
rect 10229 3479 10287 3485
rect 9677 3451 9735 3457
rect 9677 3417 9689 3451
rect 9723 3417 9735 3451
rect 10244 3448 10272 3479
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 10870 3476 10876 3528
rect 10928 3516 10934 3528
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 10928 3488 11437 3516
rect 10928 3476 10934 3488
rect 11425 3485 11437 3488
rect 11471 3516 11483 3519
rect 11698 3516 11704 3528
rect 11471 3488 11704 3516
rect 11471 3485 11483 3488
rect 11425 3479 11483 3485
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 11882 3476 11888 3528
rect 11940 3516 11946 3528
rect 12621 3519 12679 3525
rect 12621 3516 12633 3519
rect 11940 3488 12633 3516
rect 11940 3476 11946 3488
rect 12621 3485 12633 3488
rect 12667 3485 12679 3519
rect 13725 3519 13783 3525
rect 12621 3479 12679 3485
rect 12728 3488 13676 3516
rect 9677 3411 9735 3417
rect 9784 3420 10272 3448
rect 7576 3352 8892 3380
rect 9214 3340 9220 3392
rect 9272 3380 9278 3392
rect 9784 3380 9812 3420
rect 10686 3408 10692 3460
rect 10744 3448 10750 3460
rect 10744 3420 11560 3448
rect 10744 3408 10750 3420
rect 9272 3352 9812 3380
rect 9272 3340 9278 3352
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 11422 3380 11428 3392
rect 10100 3352 11428 3380
rect 10100 3340 10106 3352
rect 11422 3340 11428 3352
rect 11480 3340 11486 3392
rect 11532 3380 11560 3420
rect 12250 3408 12256 3460
rect 12308 3448 12314 3460
rect 12728 3448 12756 3488
rect 13262 3448 13268 3460
rect 12308 3420 12756 3448
rect 13223 3420 13268 3448
rect 12308 3408 12314 3420
rect 13262 3408 13268 3420
rect 13320 3408 13326 3460
rect 13648 3448 13676 3488
rect 13725 3485 13737 3519
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3485 13967 3519
rect 13909 3479 13967 3485
rect 13740 3448 13768 3479
rect 13648 3420 13768 3448
rect 13814 3408 13820 3460
rect 13872 3448 13878 3460
rect 13924 3448 13952 3479
rect 13872 3420 13952 3448
rect 13872 3408 13878 3420
rect 14645 3383 14703 3389
rect 14645 3380 14657 3383
rect 11532 3352 14657 3380
rect 14645 3349 14657 3352
rect 14691 3349 14703 3383
rect 14645 3343 14703 3349
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 2314 3136 2320 3188
rect 2372 3176 2378 3188
rect 2501 3179 2559 3185
rect 2501 3176 2513 3179
rect 2372 3148 2513 3176
rect 2372 3136 2378 3148
rect 2501 3145 2513 3148
rect 2547 3145 2559 3179
rect 2501 3139 2559 3145
rect 3697 3179 3755 3185
rect 3697 3145 3709 3179
rect 3743 3176 3755 3179
rect 4246 3176 4252 3188
rect 3743 3148 4252 3176
rect 3743 3145 3755 3148
rect 3697 3139 3755 3145
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 5534 3176 5540 3188
rect 4356 3148 5540 3176
rect 3234 3068 3240 3120
rect 3292 3108 3298 3120
rect 3292 3080 4292 3108
rect 3292 3068 3298 3080
rect 1118 3000 1124 3052
rect 1176 3000 1182 3052
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 2498 3040 2504 3052
rect 1903 3012 2504 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 3142 3040 3148 3052
rect 3103 3012 3148 3040
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 4154 3040 4160 3052
rect 4115 3012 4160 3040
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 1136 2972 1164 3000
rect 1581 2975 1639 2981
rect 1581 2972 1593 2975
rect 1136 2944 1593 2972
rect 1581 2941 1593 2944
rect 1627 2941 1639 2975
rect 4062 2972 4068 2984
rect 4023 2944 4068 2972
rect 1581 2935 1639 2941
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 4264 2972 4292 3080
rect 4356 3049 4384 3148
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 6273 3179 6331 3185
rect 6273 3145 6285 3179
rect 6319 3176 6331 3179
rect 7190 3176 7196 3188
rect 6319 3148 7196 3176
rect 6319 3145 6331 3148
rect 6273 3139 6331 3145
rect 7190 3136 7196 3148
rect 7248 3176 7254 3188
rect 8110 3176 8116 3188
rect 7248 3148 8116 3176
rect 7248 3136 7254 3148
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 12253 3179 12311 3185
rect 12253 3176 12265 3179
rect 8312 3148 12265 3176
rect 4890 3068 4896 3120
rect 4948 3068 4954 3120
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 4614 3040 4620 3052
rect 4488 3012 4620 3040
rect 4488 3000 4494 3012
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 4908 2981 4936 3068
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 6546 3040 6552 3052
rect 6328 3012 6552 3040
rect 6328 3000 6334 3012
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6788 3012 6837 3040
rect 6788 3000 6794 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 4893 2975 4951 2981
rect 4264 2944 4844 2972
rect 2961 2907 3019 2913
rect 2961 2873 2973 2907
rect 3007 2904 3019 2907
rect 4816 2904 4844 2944
rect 4893 2941 4905 2975
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 5626 2932 5632 2984
rect 5684 2972 5690 2984
rect 5684 2944 6868 2972
rect 5684 2932 5690 2944
rect 5138 2907 5196 2913
rect 5138 2904 5150 2907
rect 3007 2876 4752 2904
rect 4816 2876 5150 2904
rect 3007 2873 3019 2876
rect 2961 2867 3019 2873
rect 382 2796 388 2848
rect 440 2836 446 2848
rect 1394 2836 1400 2848
rect 440 2808 1400 2836
rect 440 2796 446 2808
rect 1394 2796 1400 2808
rect 1452 2796 1458 2848
rect 2869 2839 2927 2845
rect 2869 2805 2881 2839
rect 2915 2836 2927 2839
rect 3050 2836 3056 2848
rect 2915 2808 3056 2836
rect 2915 2805 2927 2808
rect 2869 2799 2927 2805
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 4724 2836 4752 2876
rect 5138 2873 5150 2876
rect 5184 2904 5196 2907
rect 5718 2904 5724 2916
rect 5184 2876 5724 2904
rect 5184 2873 5196 2876
rect 5138 2867 5196 2873
rect 5718 2864 5724 2876
rect 5776 2864 5782 2916
rect 6362 2864 6368 2916
rect 6420 2864 6426 2916
rect 5534 2836 5540 2848
rect 4724 2808 5540 2836
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 5626 2796 5632 2848
rect 5684 2836 5690 2848
rect 6380 2836 6408 2864
rect 5684 2808 6408 2836
rect 6840 2836 6868 2944
rect 7558 2932 7564 2984
rect 7616 2972 7622 2984
rect 8312 2972 8340 3148
rect 12253 3145 12265 3148
rect 12299 3176 12311 3179
rect 13078 3176 13084 3188
rect 12299 3148 13084 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 13633 3179 13691 3185
rect 13633 3145 13645 3179
rect 13679 3176 13691 3179
rect 13722 3176 13728 3188
rect 13679 3148 13728 3176
rect 13679 3145 13691 3148
rect 13633 3139 13691 3145
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 8662 3108 8668 3120
rect 8623 3080 8668 3108
rect 8662 3068 8668 3080
rect 8720 3068 8726 3120
rect 9766 3108 9772 3120
rect 9140 3080 9444 3108
rect 9727 3080 9772 3108
rect 9140 3049 9168 3080
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3009 9183 3043
rect 9306 3040 9312 3052
rect 9267 3012 9312 3040
rect 9125 3003 9183 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 9416 3040 9444 3080
rect 9766 3068 9772 3080
rect 9824 3108 9830 3120
rect 10042 3108 10048 3120
rect 9824 3080 10048 3108
rect 9824 3068 9830 3080
rect 10042 3068 10048 3080
rect 10100 3068 10106 3120
rect 10778 3108 10784 3120
rect 10520 3080 10784 3108
rect 10410 3040 10416 3052
rect 9416 3012 10416 3040
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 10520 3049 10548 3080
rect 10778 3068 10784 3080
rect 10836 3068 10842 3120
rect 11790 3068 11796 3120
rect 11848 3108 11854 3120
rect 11848 3080 14872 3108
rect 11848 3068 11854 3080
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 11609 3043 11667 3049
rect 11609 3040 11621 3043
rect 11020 3012 11621 3040
rect 11020 3000 11026 3012
rect 11609 3009 11621 3012
rect 11655 3040 11667 3043
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 11655 3012 13001 3040
rect 11655 3009 11667 3012
rect 11609 3003 11667 3009
rect 12989 3009 13001 3012
rect 13035 3040 13047 3043
rect 13814 3040 13820 3052
rect 13035 3012 13820 3040
rect 13035 3009 13047 3012
rect 12989 3003 13047 3009
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 14090 3040 14096 3052
rect 14051 3012 14096 3040
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 7616 2944 8340 2972
rect 7616 2932 7622 2944
rect 8386 2932 8392 2984
rect 8444 2972 8450 2984
rect 9324 2972 9352 3000
rect 8444 2944 9352 2972
rect 8444 2932 8450 2944
rect 10042 2932 10048 2984
rect 10100 2972 10106 2984
rect 10229 2975 10287 2981
rect 10229 2972 10241 2975
rect 10100 2944 10241 2972
rect 10100 2932 10106 2944
rect 10229 2941 10241 2944
rect 10275 2941 10287 2975
rect 11514 2972 11520 2984
rect 10229 2935 10287 2941
rect 10888 2944 11520 2972
rect 7006 2864 7012 2916
rect 7064 2913 7070 2916
rect 7064 2907 7128 2913
rect 7064 2873 7082 2907
rect 7116 2873 7128 2907
rect 7064 2867 7128 2873
rect 7064 2864 7070 2867
rect 7190 2864 7196 2916
rect 7248 2904 7254 2916
rect 7834 2904 7840 2916
rect 7248 2876 7840 2904
rect 7248 2864 7254 2876
rect 7834 2864 7840 2876
rect 7892 2864 7898 2916
rect 8110 2864 8116 2916
rect 8168 2904 8174 2916
rect 9214 2904 9220 2916
rect 8168 2876 9220 2904
rect 8168 2864 8174 2876
rect 9214 2864 9220 2876
rect 9272 2864 9278 2916
rect 10321 2907 10379 2913
rect 10321 2873 10333 2907
rect 10367 2904 10379 2907
rect 10888 2904 10916 2944
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 11790 2932 11796 2984
rect 11848 2972 11854 2984
rect 12805 2975 12863 2981
rect 12805 2972 12817 2975
rect 11848 2944 12817 2972
rect 11848 2932 11854 2944
rect 12805 2941 12817 2944
rect 12851 2972 12863 2975
rect 12851 2944 13124 2972
rect 12851 2941 12863 2944
rect 12805 2935 12863 2941
rect 10367 2876 10916 2904
rect 10367 2873 10379 2876
rect 10321 2867 10379 2873
rect 10962 2864 10968 2916
rect 11020 2864 11026 2916
rect 12986 2904 12992 2916
rect 11072 2876 12992 2904
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 6840 2808 8217 2836
rect 5684 2796 5690 2808
rect 8205 2805 8217 2808
rect 8251 2836 8263 2839
rect 8846 2836 8852 2848
rect 8251 2808 8852 2836
rect 8251 2805 8263 2808
rect 8205 2799 8263 2805
rect 8846 2796 8852 2808
rect 8904 2796 8910 2848
rect 8938 2796 8944 2848
rect 8996 2836 9002 2848
rect 9033 2839 9091 2845
rect 9033 2836 9045 2839
rect 8996 2808 9045 2836
rect 8996 2796 9002 2808
rect 9033 2805 9045 2808
rect 9079 2805 9091 2839
rect 9858 2836 9864 2848
rect 9819 2808 9864 2836
rect 9033 2799 9091 2805
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 10042 2796 10048 2848
rect 10100 2836 10106 2848
rect 10980 2836 11008 2864
rect 11072 2845 11100 2876
rect 12986 2864 12992 2876
rect 13044 2864 13050 2916
rect 13096 2904 13124 2944
rect 13906 2932 13912 2984
rect 13964 2972 13970 2984
rect 14292 2972 14320 3000
rect 14844 2981 14872 3080
rect 13964 2944 14320 2972
rect 14829 2975 14887 2981
rect 13964 2932 13970 2944
rect 14829 2941 14841 2975
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 15102 2904 15108 2916
rect 13096 2876 15108 2904
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 10100 2808 11008 2836
rect 11057 2839 11115 2845
rect 10100 2796 10106 2808
rect 11057 2805 11069 2839
rect 11103 2805 11115 2839
rect 11422 2836 11428 2848
rect 11383 2808 11428 2836
rect 11057 2799 11115 2805
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2836 11575 2839
rect 12253 2839 12311 2845
rect 12253 2836 12265 2839
rect 11563 2808 12265 2836
rect 11563 2805 11575 2808
rect 11517 2799 11575 2805
rect 12253 2805 12265 2808
rect 12299 2805 12311 2839
rect 12253 2799 12311 2805
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12894 2836 12900 2848
rect 12492 2808 12537 2836
rect 12855 2808 12900 2836
rect 12492 2796 12498 2808
rect 12894 2796 12900 2808
rect 12952 2796 12958 2848
rect 13630 2796 13636 2848
rect 13688 2836 13694 2848
rect 14001 2839 14059 2845
rect 14001 2836 14013 2839
rect 13688 2808 14013 2836
rect 13688 2796 13694 2808
rect 14001 2805 14013 2808
rect 14047 2805 14059 2839
rect 14001 2799 14059 2805
rect 14090 2796 14096 2848
rect 14148 2836 14154 2848
rect 15013 2839 15071 2845
rect 15013 2836 15025 2839
rect 14148 2808 15025 2836
rect 14148 2796 14154 2808
rect 15013 2805 15025 2808
rect 15059 2805 15071 2839
rect 15013 2799 15071 2805
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 5718 2592 5724 2644
rect 5776 2632 5782 2644
rect 6365 2635 6423 2641
rect 6365 2632 6377 2635
rect 5776 2604 6377 2632
rect 5776 2592 5782 2604
rect 6365 2601 6377 2604
rect 6411 2601 6423 2635
rect 6365 2595 6423 2601
rect 6454 2592 6460 2644
rect 6512 2632 6518 2644
rect 6917 2635 6975 2641
rect 6917 2632 6929 2635
rect 6512 2604 6929 2632
rect 6512 2592 6518 2604
rect 6917 2601 6929 2604
rect 6963 2601 6975 2635
rect 6917 2595 6975 2601
rect 7377 2635 7435 2641
rect 7377 2601 7389 2635
rect 7423 2632 7435 2635
rect 8018 2632 8024 2644
rect 7423 2604 8024 2632
rect 7423 2601 7435 2604
rect 7377 2595 7435 2601
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 8113 2635 8171 2641
rect 8113 2601 8125 2635
rect 8159 2601 8171 2635
rect 8113 2595 8171 2601
rect 4430 2524 4436 2576
rect 4488 2564 4494 2576
rect 5230 2567 5288 2573
rect 5230 2564 5242 2567
rect 4488 2536 5242 2564
rect 4488 2524 4494 2536
rect 5230 2533 5242 2536
rect 5276 2533 5288 2567
rect 5230 2527 5288 2533
rect 5442 2524 5448 2576
rect 5500 2524 5506 2576
rect 5534 2524 5540 2576
rect 5592 2564 5598 2576
rect 8128 2564 8156 2595
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 10134 2632 10140 2644
rect 9732 2604 9812 2632
rect 10095 2604 10140 2632
rect 9732 2592 9738 2604
rect 9784 2564 9812 2604
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10318 2632 10324 2644
rect 10275 2604 10324 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 11422 2632 11428 2644
rect 11383 2604 11428 2632
rect 11422 2592 11428 2604
rect 11480 2632 11486 2644
rect 12250 2632 12256 2644
rect 11480 2604 12256 2632
rect 11480 2592 11486 2604
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 13081 2635 13139 2641
rect 13081 2632 13093 2635
rect 12492 2604 13093 2632
rect 12492 2592 12498 2604
rect 13081 2601 13093 2604
rect 13127 2601 13139 2635
rect 13081 2595 13139 2601
rect 14182 2592 14188 2644
rect 14240 2632 14246 2644
rect 14277 2635 14335 2641
rect 14277 2632 14289 2635
rect 14240 2604 14289 2632
rect 14240 2592 14246 2604
rect 14277 2601 14289 2604
rect 14323 2601 14335 2635
rect 14277 2595 14335 2601
rect 10686 2564 10692 2576
rect 5592 2536 8156 2564
rect 8404 2536 9720 2564
rect 9784 2536 10692 2564
rect 5592 2524 5598 2536
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 2400 2499 2458 2505
rect 2400 2465 2412 2499
rect 2446 2496 2458 2499
rect 2866 2496 2872 2508
rect 2446 2468 2872 2496
rect 2446 2465 2458 2468
rect 2400 2459 2458 2465
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 3970 2456 3976 2508
rect 4028 2496 4034 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 4028 2468 4077 2496
rect 4028 2456 4034 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4614 2456 4620 2508
rect 4672 2496 4678 2508
rect 5460 2496 5488 2524
rect 4672 2468 5488 2496
rect 7285 2499 7343 2505
rect 4672 2456 4678 2468
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2397 2191 2431
rect 4338 2428 4344 2440
rect 4299 2400 4344 2428
rect 2133 2391 2191 2397
rect 106 2252 112 2304
rect 164 2292 170 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 164 2264 1593 2292
rect 164 2252 170 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 2148 2292 2176 2391
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 4632 2360 4660 2456
rect 5000 2440 5028 2468
rect 7285 2465 7297 2499
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 4982 2428 4988 2440
rect 4943 2400 4988 2428
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 3344 2332 4660 2360
rect 3344 2292 3372 2332
rect 2148 2264 3372 2292
rect 3513 2295 3571 2301
rect 1581 2255 1639 2261
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 7006 2292 7012 2304
rect 3559 2264 7012 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 7300 2292 7328 2459
rect 7650 2456 7656 2508
rect 7708 2496 7714 2508
rect 8404 2496 8432 2536
rect 7708 2468 8432 2496
rect 8481 2499 8539 2505
rect 7708 2456 7714 2468
rect 8481 2465 8493 2499
rect 8527 2496 8539 2499
rect 9030 2496 9036 2508
rect 8527 2468 9036 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 9030 2456 9036 2468
rect 9088 2456 9094 2508
rect 9490 2496 9496 2508
rect 9451 2468 9496 2496
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 9692 2496 9720 2536
rect 10686 2524 10692 2536
rect 10744 2524 10750 2576
rect 11333 2567 11391 2573
rect 11333 2533 11345 2567
rect 11379 2564 11391 2567
rect 12158 2564 12164 2576
rect 11379 2536 12164 2564
rect 11379 2533 11391 2536
rect 11333 2527 11391 2533
rect 12158 2524 12164 2536
rect 12216 2524 12222 2576
rect 12710 2564 12716 2576
rect 12268 2536 12716 2564
rect 9692 2468 11560 2496
rect 7466 2428 7472 2440
rect 7427 2400 7472 2428
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 8570 2428 8576 2440
rect 8168 2400 8576 2428
rect 8168 2388 8174 2400
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 7374 2320 7380 2372
rect 7432 2360 7438 2372
rect 8680 2360 8708 2391
rect 9306 2388 9312 2440
rect 9364 2428 9370 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 9364 2400 10333 2428
rect 9364 2388 9370 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 11330 2388 11336 2440
rect 11388 2428 11394 2440
rect 11532 2437 11560 2468
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 11388 2400 11529 2428
rect 11388 2388 11394 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 10410 2360 10416 2372
rect 7432 2332 8708 2360
rect 9232 2332 10416 2360
rect 7432 2320 7438 2332
rect 9232 2292 9260 2332
rect 10410 2320 10416 2332
rect 10468 2320 10474 2372
rect 10965 2363 11023 2369
rect 10965 2329 10977 2363
rect 11011 2360 11023 2363
rect 12268 2360 12296 2536
rect 12710 2524 12716 2536
rect 12768 2524 12774 2576
rect 12986 2564 12992 2576
rect 12947 2536 12992 2564
rect 12986 2524 12992 2536
rect 13044 2524 13050 2576
rect 12345 2499 12403 2505
rect 12345 2465 12357 2499
rect 12391 2465 12403 2499
rect 12345 2459 12403 2465
rect 11011 2332 12296 2360
rect 11011 2329 11023 2332
rect 10965 2323 11023 2329
rect 7300 2264 9260 2292
rect 9306 2252 9312 2304
rect 9364 2292 9370 2304
rect 9766 2292 9772 2304
rect 9364 2264 9409 2292
rect 9727 2264 9772 2292
rect 9364 2252 9370 2264
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 10428 2292 10456 2320
rect 11330 2292 11336 2304
rect 10428 2264 11336 2292
rect 11330 2252 11336 2264
rect 11388 2252 11394 2304
rect 12158 2292 12164 2304
rect 12119 2264 12164 2292
rect 12158 2252 12164 2264
rect 12216 2252 12222 2304
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 12360 2292 12388 2459
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 12492 2468 14197 2496
rect 12492 2456 12498 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 15197 2499 15255 2505
rect 15197 2465 15209 2499
rect 15243 2496 15255 2499
rect 15286 2496 15292 2508
rect 15243 2468 15292 2496
rect 15243 2465 15255 2468
rect 15197 2459 15255 2465
rect 15286 2456 15292 2468
rect 15344 2456 15350 2508
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 12452 2400 13277 2428
rect 12452 2372 12480 2400
rect 13265 2397 13277 2400
rect 13311 2428 13323 2431
rect 13906 2428 13912 2440
rect 13311 2400 13912 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 13906 2388 13912 2400
rect 13964 2428 13970 2440
rect 14369 2431 14427 2437
rect 14369 2428 14381 2431
rect 13964 2400 14381 2428
rect 13964 2388 13970 2400
rect 14369 2397 14381 2400
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 12434 2320 12440 2372
rect 12492 2320 12498 2372
rect 12621 2363 12679 2369
rect 12621 2329 12633 2363
rect 12667 2360 12679 2363
rect 12802 2360 12808 2372
rect 12667 2332 12808 2360
rect 12667 2329 12679 2332
rect 12621 2323 12679 2329
rect 12802 2320 12808 2332
rect 12860 2320 12866 2372
rect 13722 2320 13728 2372
rect 13780 2360 13786 2372
rect 14274 2360 14280 2372
rect 13780 2332 14280 2360
rect 13780 2320 13786 2332
rect 14274 2320 14280 2332
rect 14332 2320 14338 2372
rect 13814 2292 13820 2304
rect 12308 2264 12388 2292
rect 13775 2264 13820 2292
rect 12308 2252 12314 2264
rect 13814 2252 13820 2264
rect 13872 2252 13878 2304
rect 13906 2252 13912 2304
rect 13964 2292 13970 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 13964 2264 15025 2292
rect 13964 2252 13970 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 7926 2048 7932 2100
rect 7984 2088 7990 2100
rect 8938 2088 8944 2100
rect 7984 2060 8944 2088
rect 7984 2048 7990 2060
rect 8938 2048 8944 2060
rect 8996 2048 9002 2100
rect 10226 2048 10232 2100
rect 10284 2088 10290 2100
rect 13906 2088 13912 2100
rect 10284 2060 13912 2088
rect 10284 2048 10290 2060
rect 13906 2048 13912 2060
rect 13964 2048 13970 2100
rect 8570 1980 8576 2032
rect 8628 2020 8634 2032
rect 9122 2020 9128 2032
rect 8628 1992 9128 2020
rect 8628 1980 8634 1992
rect 9122 1980 9128 1992
rect 9180 1980 9186 2032
rect 9306 1980 9312 2032
rect 9364 2020 9370 2032
rect 12250 2020 12256 2032
rect 9364 1992 12256 2020
rect 9364 1980 9370 1992
rect 12250 1980 12256 1992
rect 12308 1980 12314 2032
rect 12526 1980 12532 2032
rect 12584 2020 12590 2032
rect 13354 2020 13360 2032
rect 12584 1992 13360 2020
rect 12584 1980 12590 1992
rect 13354 1980 13360 1992
rect 13412 1980 13418 2032
rect 4338 1912 4344 1964
rect 4396 1952 4402 1964
rect 16022 1952 16028 1964
rect 4396 1924 16028 1952
rect 4396 1912 4402 1924
rect 16022 1912 16028 1924
rect 16080 1912 16086 1964
rect 6914 1844 6920 1896
rect 6972 1884 6978 1896
rect 8110 1884 8116 1896
rect 6972 1856 8116 1884
rect 6972 1844 6978 1856
rect 8110 1844 8116 1856
rect 8168 1844 8174 1896
rect 10318 1844 10324 1896
rect 10376 1884 10382 1896
rect 13630 1884 13636 1896
rect 10376 1856 13636 1884
rect 10376 1844 10382 1856
rect 13630 1844 13636 1856
rect 13688 1844 13694 1896
rect 2958 1776 2964 1828
rect 3016 1816 3022 1828
rect 9306 1816 9312 1828
rect 3016 1788 9312 1816
rect 3016 1776 3022 1788
rect 9306 1776 9312 1788
rect 9364 1776 9370 1828
rect 9766 1776 9772 1828
rect 9824 1816 9830 1828
rect 14826 1816 14832 1828
rect 9824 1788 14832 1816
rect 9824 1776 9830 1788
rect 14826 1776 14832 1788
rect 14884 1776 14890 1828
rect 1854 1708 1860 1760
rect 1912 1748 1918 1760
rect 13814 1748 13820 1760
rect 1912 1720 13820 1748
rect 1912 1708 1918 1720
rect 13814 1708 13820 1720
rect 13872 1708 13878 1760
rect 1394 1640 1400 1692
rect 1452 1680 1458 1692
rect 9030 1680 9036 1692
rect 1452 1652 9036 1680
rect 1452 1640 1458 1652
rect 9030 1640 9036 1652
rect 9088 1640 9094 1692
rect 4982 1572 4988 1624
rect 5040 1612 5046 1624
rect 12158 1612 12164 1624
rect 5040 1584 12164 1612
rect 5040 1572 5046 1584
rect 12158 1572 12164 1584
rect 12216 1572 12222 1624
rect 8202 1504 8208 1556
rect 8260 1544 8266 1556
rect 11422 1544 11428 1556
rect 8260 1516 11428 1544
rect 8260 1504 8266 1516
rect 11422 1504 11428 1516
rect 11480 1504 11486 1556
rect 3142 1232 3148 1284
rect 3200 1272 3206 1284
rect 5074 1272 5080 1284
rect 3200 1244 5080 1272
rect 3200 1232 3206 1244
rect 5074 1232 5080 1244
rect 5132 1232 5138 1284
rect 3510 960 3516 1012
rect 3568 1000 3574 1012
rect 7282 1000 7288 1012
rect 3568 972 7288 1000
rect 3568 960 3574 972
rect 7282 960 7288 972
rect 7340 960 7346 1012
<< via1 >>
rect 7564 18436 7616 18488
rect 9404 18436 9456 18488
rect 11428 18096 11480 18148
rect 12072 18096 12124 18148
rect 9680 18028 9732 18080
rect 14464 18028 14516 18080
rect 16028 18028 16080 18080
rect 4068 17960 4120 18012
rect 13912 17960 13964 18012
rect 7932 17892 7984 17944
rect 8852 17892 8904 17944
rect 8944 17892 8996 17944
rect 12808 17892 12860 17944
rect 5172 17824 5224 17876
rect 9128 17824 9180 17876
rect 7840 17756 7892 17808
rect 13176 17756 13228 17808
rect 6920 17688 6972 17740
rect 14280 17688 14332 17740
rect 5448 17620 5500 17672
rect 12716 17620 12768 17672
rect 3516 17552 3568 17604
rect 9864 17552 9916 17604
rect 5724 17484 5776 17536
rect 9312 17484 9364 17536
rect 10232 17484 10284 17536
rect 11796 17484 11848 17536
rect 14372 17484 14424 17536
rect 3447 17382 3499 17434
rect 3511 17382 3563 17434
rect 3575 17382 3627 17434
rect 3639 17382 3691 17434
rect 8378 17382 8430 17434
rect 8442 17382 8494 17434
rect 8506 17382 8558 17434
rect 8570 17382 8622 17434
rect 13308 17382 13360 17434
rect 13372 17382 13424 17434
rect 13436 17382 13488 17434
rect 13500 17382 13552 17434
rect 6184 17280 6236 17332
rect 2412 17212 2464 17264
rect 756 17144 808 17196
rect 1492 17119 1544 17128
rect 1492 17085 1501 17119
rect 1501 17085 1535 17119
rect 1535 17085 1544 17119
rect 1492 17076 1544 17085
rect 2136 17144 2188 17196
rect 3792 17212 3844 17264
rect 6368 17212 6420 17264
rect 3148 17144 3200 17196
rect 4988 17187 5040 17196
rect 4988 17153 4997 17187
rect 4997 17153 5031 17187
rect 5031 17153 5040 17187
rect 4988 17144 5040 17153
rect 7472 17187 7524 17196
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 7472 17144 7524 17153
rect 7656 17212 7708 17264
rect 8944 17212 8996 17264
rect 9404 17212 9456 17264
rect 8024 17144 8076 17196
rect 2688 17076 2740 17128
rect 3240 17076 3292 17128
rect 4068 17119 4120 17128
rect 4068 17085 4077 17119
rect 4077 17085 4111 17119
rect 4111 17085 4120 17119
rect 4068 17076 4120 17085
rect 5540 17076 5592 17128
rect 8852 17076 8904 17128
rect 9496 17119 9548 17128
rect 9496 17085 9505 17119
rect 9505 17085 9539 17119
rect 9539 17085 9548 17119
rect 9496 17076 9548 17085
rect 10048 17076 10100 17128
rect 10416 17076 10468 17128
rect 12532 17076 12584 17128
rect 13084 17076 13136 17128
rect 1860 17008 1912 17060
rect 2964 17008 3016 17060
rect 6276 17008 6328 17060
rect 7932 17008 7984 17060
rect 8484 17051 8536 17060
rect 8484 17017 8493 17051
rect 8493 17017 8527 17051
rect 8527 17017 8536 17051
rect 8484 17008 8536 17017
rect 8760 17008 8812 17060
rect 9588 17008 9640 17060
rect 11428 17008 11480 17060
rect 11704 17008 11756 17060
rect 3332 16983 3384 16992
rect 3332 16949 3341 16983
rect 3341 16949 3375 16983
rect 3375 16949 3384 16983
rect 3332 16940 3384 16949
rect 5632 16983 5684 16992
rect 5632 16949 5641 16983
rect 5641 16949 5675 16983
rect 5675 16949 5684 16983
rect 5632 16940 5684 16949
rect 5724 16940 5776 16992
rect 7748 16940 7800 16992
rect 9772 16940 9824 16992
rect 10140 16940 10192 16992
rect 11152 16940 11204 16992
rect 11888 16940 11940 16992
rect 12900 16940 12952 16992
rect 5912 16838 5964 16890
rect 5976 16838 6028 16890
rect 6040 16838 6092 16890
rect 6104 16838 6156 16890
rect 10843 16838 10895 16890
rect 10907 16838 10959 16890
rect 10971 16838 11023 16890
rect 11035 16838 11087 16890
rect 2780 16736 2832 16788
rect 1676 16711 1728 16720
rect 1676 16677 1685 16711
rect 1685 16677 1719 16711
rect 1719 16677 1728 16711
rect 1676 16668 1728 16677
rect 4620 16736 4672 16788
rect 5448 16779 5500 16788
rect 5448 16745 5457 16779
rect 5457 16745 5491 16779
rect 5491 16745 5500 16779
rect 5448 16736 5500 16745
rect 6276 16779 6328 16788
rect 6276 16745 6285 16779
rect 6285 16745 6319 16779
rect 6319 16745 6328 16779
rect 6276 16736 6328 16745
rect 7840 16779 7892 16788
rect 7840 16745 7849 16779
rect 7849 16745 7883 16779
rect 7883 16745 7892 16779
rect 7840 16736 7892 16745
rect 8116 16736 8168 16788
rect 8300 16736 8352 16788
rect 8852 16736 8904 16788
rect 3332 16668 3384 16720
rect 1584 16600 1636 16652
rect 2596 16600 2648 16652
rect 1124 16532 1176 16584
rect 1492 16532 1544 16584
rect 3976 16600 4028 16652
rect 4528 16668 4580 16720
rect 4252 16600 4304 16652
rect 5356 16643 5408 16652
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 5356 16600 5408 16609
rect 7656 16668 7708 16720
rect 9036 16668 9088 16720
rect 9312 16668 9364 16720
rect 1584 16464 1636 16516
rect 3240 16464 3292 16516
rect 3884 16464 3936 16516
rect 5080 16464 5132 16516
rect 6644 16532 6696 16584
rect 7196 16532 7248 16584
rect 7656 16532 7708 16584
rect 7748 16532 7800 16584
rect 8852 16600 8904 16652
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 8208 16464 8260 16516
rect 9772 16464 9824 16516
rect 9864 16507 9916 16516
rect 9864 16473 9873 16507
rect 9873 16473 9907 16507
rect 9907 16473 9916 16507
rect 10140 16532 10192 16584
rect 11428 16736 11480 16788
rect 12256 16736 12308 16788
rect 14280 16779 14332 16788
rect 14280 16745 14289 16779
rect 14289 16745 14323 16779
rect 14323 16745 14332 16779
rect 14280 16736 14332 16745
rect 12164 16668 12216 16720
rect 11520 16600 11572 16652
rect 11888 16643 11940 16652
rect 11888 16609 11897 16643
rect 11897 16609 11931 16643
rect 11931 16609 11940 16643
rect 11888 16600 11940 16609
rect 12072 16600 12124 16652
rect 12440 16600 12492 16652
rect 14096 16643 14148 16652
rect 14096 16609 14105 16643
rect 14105 16609 14139 16643
rect 14139 16609 14148 16643
rect 14096 16600 14148 16609
rect 9864 16464 9916 16473
rect 12808 16507 12860 16516
rect 12808 16473 12817 16507
rect 12817 16473 12851 16507
rect 12851 16473 12860 16507
rect 12808 16464 12860 16473
rect 3792 16396 3844 16448
rect 6368 16396 6420 16448
rect 7840 16396 7892 16448
rect 8024 16396 8076 16448
rect 8668 16396 8720 16448
rect 11428 16396 11480 16448
rect 3447 16294 3499 16346
rect 3511 16294 3563 16346
rect 3575 16294 3627 16346
rect 3639 16294 3691 16346
rect 8378 16294 8430 16346
rect 8442 16294 8494 16346
rect 8506 16294 8558 16346
rect 8570 16294 8622 16346
rect 13308 16294 13360 16346
rect 13372 16294 13424 16346
rect 13436 16294 13488 16346
rect 13500 16294 13552 16346
rect 1860 16192 1912 16244
rect 4068 16192 4120 16244
rect 4712 16192 4764 16244
rect 4804 16192 4856 16244
rect 9864 16192 9916 16244
rect 9956 16192 10008 16244
rect 11244 16192 11296 16244
rect 12348 16192 12400 16244
rect 5816 16124 5868 16176
rect 1400 16056 1452 16108
rect 1768 16056 1820 16108
rect 5540 16056 5592 16108
rect 5632 16056 5684 16108
rect 6644 16124 6696 16176
rect 6828 16167 6880 16176
rect 6828 16133 6837 16167
rect 6837 16133 6871 16167
rect 6871 16133 6880 16167
rect 6828 16124 6880 16133
rect 6920 16124 6972 16176
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 7564 16056 7616 16108
rect 7932 16056 7984 16108
rect 8484 16056 8536 16108
rect 112 15988 164 16040
rect 1308 15988 1360 16040
rect 2412 16031 2464 16040
rect 388 15920 440 15972
rect 2412 15997 2444 16031
rect 2444 15997 2464 16031
rect 2412 15988 2464 15997
rect 4436 15988 4488 16040
rect 7196 16031 7248 16040
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 7748 15988 7800 16040
rect 8300 15988 8352 16040
rect 3608 15963 3660 15972
rect 3608 15929 3617 15963
rect 3617 15929 3651 15963
rect 3651 15929 3660 15963
rect 3608 15920 3660 15929
rect 4712 15963 4764 15972
rect 4712 15929 4721 15963
rect 4721 15929 4755 15963
rect 4755 15929 4764 15963
rect 4712 15920 4764 15929
rect 6184 15920 6236 15972
rect 7564 15920 7616 15972
rect 9128 16056 9180 16108
rect 10784 16124 10836 16176
rect 12900 16124 12952 16176
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 5172 15852 5224 15904
rect 7380 15852 7432 15904
rect 8392 15895 8444 15904
rect 8392 15861 8401 15895
rect 8401 15861 8435 15895
rect 8435 15861 8444 15895
rect 8392 15852 8444 15861
rect 9128 15920 9180 15972
rect 10692 16056 10744 16108
rect 10232 15988 10284 16040
rect 11336 15988 11388 16040
rect 12348 15988 12400 16040
rect 8760 15852 8812 15904
rect 9496 15852 9548 15904
rect 11888 15920 11940 15972
rect 12072 15920 12124 15972
rect 11428 15852 11480 15904
rect 5912 15750 5964 15802
rect 5976 15750 6028 15802
rect 6040 15750 6092 15802
rect 6104 15750 6156 15802
rect 10843 15750 10895 15802
rect 10907 15750 10959 15802
rect 10971 15750 11023 15802
rect 11035 15750 11087 15802
rect 3056 15648 3108 15700
rect 4528 15648 4580 15700
rect 7288 15648 7340 15700
rect 8116 15691 8168 15700
rect 8116 15657 8125 15691
rect 8125 15657 8159 15691
rect 8159 15657 8168 15691
rect 8116 15648 8168 15657
rect 6828 15580 6880 15632
rect 8208 15580 8260 15632
rect 9772 15580 9824 15632
rect 12256 15648 12308 15700
rect 11244 15580 11296 15632
rect 1492 15512 1544 15564
rect 3240 15555 3292 15564
rect 3240 15521 3249 15555
rect 3249 15521 3283 15555
rect 3283 15521 3292 15555
rect 3240 15512 3292 15521
rect 8024 15555 8076 15564
rect 2044 15444 2096 15496
rect 4344 15444 4396 15496
rect 5724 15444 5776 15496
rect 8024 15521 8033 15555
rect 8033 15521 8067 15555
rect 8067 15521 8076 15555
rect 8024 15512 8076 15521
rect 8484 15512 8536 15564
rect 9312 15512 9364 15564
rect 10232 15512 10284 15564
rect 10600 15512 10652 15564
rect 11428 15512 11480 15564
rect 11796 15512 11848 15564
rect 12256 15512 12308 15564
rect 2688 15376 2740 15428
rect 4988 15376 5040 15428
rect 5632 15376 5684 15428
rect 8116 15444 8168 15496
rect 8300 15444 8352 15496
rect 8668 15444 8720 15496
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 10692 15444 10744 15496
rect 11704 15444 11756 15496
rect 12900 15444 12952 15496
rect 14004 15444 14056 15496
rect 2320 15308 2372 15360
rect 4160 15308 4212 15360
rect 5356 15308 5408 15360
rect 8392 15376 8444 15428
rect 9220 15376 9272 15428
rect 11796 15419 11848 15428
rect 11796 15385 11805 15419
rect 11805 15385 11839 15419
rect 11839 15385 11848 15419
rect 11796 15376 11848 15385
rect 6920 15308 6972 15360
rect 7196 15308 7248 15360
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 7840 15308 7892 15360
rect 9772 15308 9824 15360
rect 3447 15206 3499 15258
rect 3511 15206 3563 15258
rect 3575 15206 3627 15258
rect 3639 15206 3691 15258
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 13308 15206 13360 15258
rect 13372 15206 13424 15258
rect 13436 15206 13488 15258
rect 13500 15206 13552 15258
rect 4804 15104 4856 15156
rect 3424 15036 3476 15088
rect 5264 15104 5316 15156
rect 3056 14968 3108 15020
rect 4160 15011 4212 15020
rect 4160 14977 4169 15011
rect 4169 14977 4203 15011
rect 4203 14977 4212 15011
rect 4160 14968 4212 14977
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 1860 14900 1912 14952
rect 3792 14900 3844 14952
rect 4988 14900 5040 14952
rect 8668 15147 8720 15156
rect 8668 15113 8677 15147
rect 8677 15113 8711 15147
rect 8711 15113 8720 15147
rect 8668 15104 8720 15113
rect 9128 15104 9180 15156
rect 9956 15104 10008 15156
rect 10876 15104 10928 15156
rect 8024 15036 8076 15088
rect 11060 15079 11112 15088
rect 11060 15045 11069 15079
rect 11069 15045 11103 15079
rect 11103 15045 11112 15079
rect 11060 15036 11112 15045
rect 6552 14968 6604 15020
rect 3240 14832 3292 14884
rect 4160 14832 4212 14884
rect 6736 14900 6788 14952
rect 8116 14968 8168 15020
rect 9220 15011 9272 15020
rect 9220 14977 9229 15011
rect 9229 14977 9263 15011
rect 9263 14977 9272 15011
rect 9220 14968 9272 14977
rect 9496 14968 9548 15020
rect 11520 15011 11572 15020
rect 11520 14977 11529 15011
rect 11529 14977 11563 15011
rect 11563 14977 11572 15011
rect 11520 14968 11572 14977
rect 11796 14968 11848 15020
rect 7564 14900 7616 14952
rect 12440 14900 12492 14952
rect 8300 14832 8352 14884
rect 8392 14832 8444 14884
rect 9956 14832 10008 14884
rect 10508 14832 10560 14884
rect 5448 14764 5500 14816
rect 8116 14764 8168 14816
rect 8668 14764 8720 14816
rect 9312 14764 9364 14816
rect 10140 14764 10192 14816
rect 10600 14764 10652 14816
rect 11704 14764 11756 14816
rect 12440 14807 12492 14816
rect 12440 14773 12449 14807
rect 12449 14773 12483 14807
rect 12483 14773 12492 14807
rect 14372 14807 14424 14816
rect 12440 14764 12492 14773
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 5912 14662 5964 14714
rect 5976 14662 6028 14714
rect 6040 14662 6092 14714
rect 6104 14662 6156 14714
rect 10843 14662 10895 14714
rect 10907 14662 10959 14714
rect 10971 14662 11023 14714
rect 11035 14662 11087 14714
rect 2780 14492 2832 14544
rect 6644 14560 6696 14612
rect 7472 14560 7524 14612
rect 7564 14560 7616 14612
rect 9588 14560 9640 14612
rect 4804 14467 4856 14476
rect 3424 14399 3476 14408
rect 3424 14365 3433 14399
rect 3433 14365 3467 14399
rect 3467 14365 3476 14399
rect 3424 14356 3476 14365
rect 4804 14433 4813 14467
rect 4813 14433 4847 14467
rect 4847 14433 4856 14467
rect 4804 14424 4856 14433
rect 4896 14467 4948 14476
rect 4896 14433 4905 14467
rect 4905 14433 4939 14467
rect 4939 14433 4948 14467
rect 5540 14492 5592 14544
rect 6276 14492 6328 14544
rect 6828 14492 6880 14544
rect 13268 14560 13320 14612
rect 4896 14424 4948 14433
rect 7564 14424 7616 14476
rect 7748 14467 7800 14476
rect 7748 14433 7782 14467
rect 7782 14433 7800 14467
rect 7748 14424 7800 14433
rect 8300 14424 8352 14476
rect 4712 14288 4764 14340
rect 5540 14356 5592 14408
rect 5632 14399 5684 14408
rect 5632 14365 5641 14399
rect 5641 14365 5675 14399
rect 5675 14365 5684 14399
rect 5632 14356 5684 14365
rect 6828 14356 6880 14408
rect 9588 14424 9640 14476
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 11152 14424 11204 14476
rect 11796 14424 11848 14476
rect 12716 14424 12768 14476
rect 13636 14424 13688 14476
rect 9864 14356 9916 14408
rect 10140 14399 10192 14408
rect 10140 14365 10149 14399
rect 10149 14365 10183 14399
rect 10183 14365 10192 14399
rect 10140 14356 10192 14365
rect 1676 14220 1728 14272
rect 4252 14220 4304 14272
rect 4436 14263 4488 14272
rect 4436 14229 4445 14263
rect 4445 14229 4479 14263
rect 4479 14229 4488 14263
rect 4436 14220 4488 14229
rect 8668 14288 8720 14340
rect 8944 14288 8996 14340
rect 9220 14288 9272 14340
rect 10968 14356 11020 14408
rect 10692 14288 10744 14340
rect 8760 14220 8812 14272
rect 9404 14220 9456 14272
rect 9864 14220 9916 14272
rect 11704 14220 11756 14272
rect 15016 14220 15068 14272
rect 3447 14118 3499 14170
rect 3511 14118 3563 14170
rect 3575 14118 3627 14170
rect 3639 14118 3691 14170
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 13308 14118 13360 14170
rect 13372 14118 13424 14170
rect 13436 14118 13488 14170
rect 13500 14118 13552 14170
rect 3332 14016 3384 14068
rect 4804 14016 4856 14068
rect 5172 14016 5224 14068
rect 6276 14059 6328 14068
rect 6276 14025 6285 14059
rect 6285 14025 6319 14059
rect 6319 14025 6328 14059
rect 6276 14016 6328 14025
rect 7564 14016 7616 14068
rect 7932 13948 7984 14000
rect 10140 14016 10192 14068
rect 10692 14016 10744 14068
rect 11060 14016 11112 14068
rect 4252 13880 4304 13932
rect 4528 13880 4580 13932
rect 6828 13923 6880 13932
rect 6828 13889 6837 13923
rect 6837 13889 6871 13923
rect 6871 13889 6880 13923
rect 6828 13880 6880 13889
rect 8116 13880 8168 13932
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 2504 13812 2556 13864
rect 4988 13812 5040 13864
rect 6736 13812 6788 13864
rect 7472 13812 7524 13864
rect 8668 13855 8720 13864
rect 5264 13744 5316 13796
rect 6368 13744 6420 13796
rect 6828 13744 6880 13796
rect 8668 13821 8677 13855
rect 8677 13821 8711 13855
rect 8711 13821 8720 13855
rect 8668 13812 8720 13821
rect 9680 13880 9732 13932
rect 9956 13880 10008 13932
rect 14924 13948 14976 14000
rect 13268 13880 13320 13932
rect 8116 13744 8168 13796
rect 12348 13812 12400 13864
rect 12716 13812 12768 13864
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 14188 13812 14240 13864
rect 14464 13812 14516 13864
rect 10324 13744 10376 13796
rect 10876 13787 10928 13796
rect 10876 13753 10885 13787
rect 10885 13753 10919 13787
rect 10919 13753 10928 13787
rect 10876 13744 10928 13753
rect 10968 13744 11020 13796
rect 2964 13676 3016 13728
rect 7656 13676 7708 13728
rect 8392 13676 8444 13728
rect 9588 13676 9640 13728
rect 9772 13676 9824 13728
rect 11152 13676 11204 13728
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 15292 13676 15344 13728
rect 15752 13676 15804 13728
rect 5912 13574 5964 13626
rect 5976 13574 6028 13626
rect 6040 13574 6092 13626
rect 6104 13574 6156 13626
rect 10843 13574 10895 13626
rect 10907 13574 10959 13626
rect 10971 13574 11023 13626
rect 11035 13574 11087 13626
rect 1676 13472 1728 13524
rect 2688 13336 2740 13388
rect 2964 13472 3016 13524
rect 4804 13472 4856 13524
rect 6736 13472 6788 13524
rect 8392 13515 8444 13524
rect 8392 13481 8401 13515
rect 8401 13481 8435 13515
rect 8435 13481 8444 13515
rect 8392 13472 8444 13481
rect 8668 13472 8720 13524
rect 9588 13472 9640 13524
rect 10692 13472 10744 13524
rect 11704 13472 11756 13524
rect 13084 13515 13136 13524
rect 13084 13481 13093 13515
rect 13093 13481 13127 13515
rect 13127 13481 13136 13515
rect 13084 13472 13136 13481
rect 13176 13515 13228 13524
rect 13176 13481 13185 13515
rect 13185 13481 13219 13515
rect 13219 13481 13228 13515
rect 13176 13472 13228 13481
rect 3332 13404 3384 13456
rect 2228 13311 2280 13320
rect 2228 13277 2237 13311
rect 2237 13277 2271 13311
rect 2271 13277 2280 13311
rect 2228 13268 2280 13277
rect 2780 13268 2832 13320
rect 3148 13132 3200 13184
rect 5448 13404 5500 13456
rect 5540 13404 5592 13456
rect 6276 13404 6328 13456
rect 6920 13404 6972 13456
rect 3792 13336 3844 13388
rect 5816 13336 5868 13388
rect 6828 13336 6880 13388
rect 7288 13336 7340 13388
rect 7656 13336 7708 13388
rect 9404 13379 9456 13388
rect 8024 13268 8076 13320
rect 9128 13268 9180 13320
rect 9404 13345 9413 13379
rect 9413 13345 9447 13379
rect 9447 13345 9456 13379
rect 9404 13336 9456 13345
rect 9680 13404 9732 13456
rect 9772 13336 9824 13388
rect 10140 13404 10192 13456
rect 5632 13200 5684 13252
rect 7472 13200 7524 13252
rect 7104 13132 7156 13184
rect 7564 13175 7616 13184
rect 7564 13141 7573 13175
rect 7573 13141 7607 13175
rect 7607 13141 7616 13175
rect 7564 13132 7616 13141
rect 9312 13200 9364 13252
rect 10968 13336 11020 13388
rect 10968 13200 11020 13252
rect 11704 13336 11756 13388
rect 12532 13336 12584 13388
rect 13912 13379 13964 13388
rect 11796 13268 11848 13320
rect 12256 13268 12308 13320
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 13912 13345 13921 13379
rect 13921 13345 13955 13379
rect 13955 13345 13964 13379
rect 13912 13336 13964 13345
rect 14464 13268 14516 13320
rect 15384 13268 15436 13320
rect 9404 13132 9456 13184
rect 9680 13132 9732 13184
rect 3447 13030 3499 13082
rect 3511 13030 3563 13082
rect 3575 13030 3627 13082
rect 3639 13030 3691 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 13308 13030 13360 13082
rect 13372 13030 13424 13082
rect 13436 13030 13488 13082
rect 13500 13030 13552 13082
rect 6276 12971 6328 12980
rect 6276 12937 6285 12971
rect 6285 12937 6319 12971
rect 6319 12937 6328 12971
rect 6276 12928 6328 12937
rect 6552 12860 6604 12912
rect 6644 12792 6696 12844
rect 8024 12928 8076 12980
rect 9864 12860 9916 12912
rect 10140 12860 10192 12912
rect 10968 12860 11020 12912
rect 8668 12835 8720 12844
rect 8668 12801 8677 12835
rect 8677 12801 8711 12835
rect 8711 12801 8720 12835
rect 8668 12792 8720 12801
rect 9680 12792 9732 12844
rect 13268 12860 13320 12912
rect 11704 12835 11756 12844
rect 3700 12724 3752 12776
rect 3148 12656 3200 12708
rect 3792 12656 3844 12708
rect 5172 12699 5224 12708
rect 2228 12631 2280 12640
rect 2228 12597 2237 12631
rect 2237 12597 2271 12631
rect 2271 12597 2280 12631
rect 2228 12588 2280 12597
rect 5172 12665 5206 12699
rect 5206 12665 5224 12699
rect 5172 12656 5224 12665
rect 5264 12588 5316 12640
rect 6920 12724 6972 12776
rect 8116 12724 8168 12776
rect 8576 12724 8628 12776
rect 10048 12724 10100 12776
rect 7656 12656 7708 12708
rect 7748 12588 7800 12640
rect 7932 12656 7984 12708
rect 9496 12656 9548 12708
rect 9680 12656 9732 12708
rect 10784 12656 10836 12708
rect 10140 12588 10192 12640
rect 10600 12588 10652 12640
rect 10692 12588 10744 12640
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 12256 12792 12308 12844
rect 13636 12792 13688 12844
rect 11796 12724 11848 12776
rect 14832 12767 14884 12776
rect 14832 12733 14841 12767
rect 14841 12733 14875 12767
rect 14875 12733 14884 12767
rect 14832 12724 14884 12733
rect 12716 12656 12768 12708
rect 13176 12656 13228 12708
rect 15752 12656 15804 12708
rect 12624 12588 12676 12640
rect 14280 12588 14332 12640
rect 15016 12631 15068 12640
rect 15016 12597 15025 12631
rect 15025 12597 15059 12631
rect 15059 12597 15068 12631
rect 15016 12588 15068 12597
rect 5912 12486 5964 12538
rect 5976 12486 6028 12538
rect 6040 12486 6092 12538
rect 6104 12486 6156 12538
rect 10843 12486 10895 12538
rect 10907 12486 10959 12538
rect 10971 12486 11023 12538
rect 11035 12486 11087 12538
rect 2780 12427 2832 12436
rect 2780 12393 2789 12427
rect 2789 12393 2823 12427
rect 2823 12393 2832 12427
rect 3148 12427 3200 12436
rect 2780 12384 2832 12393
rect 3148 12393 3157 12427
rect 3157 12393 3191 12427
rect 3191 12393 3200 12427
rect 3148 12384 3200 12393
rect 5540 12316 5592 12368
rect 5632 12316 5684 12368
rect 6368 12384 6420 12436
rect 8852 12384 8904 12436
rect 9128 12384 9180 12436
rect 9312 12384 9364 12436
rect 9588 12384 9640 12436
rect 11520 12384 11572 12436
rect 12348 12384 12400 12436
rect 12532 12427 12584 12436
rect 12532 12393 12541 12427
rect 12541 12393 12575 12427
rect 12575 12393 12584 12427
rect 12532 12384 12584 12393
rect 7380 12316 7432 12368
rect 7656 12359 7708 12368
rect 7656 12325 7690 12359
rect 7690 12325 7708 12359
rect 7656 12316 7708 12325
rect 4712 12291 4764 12300
rect 4712 12257 4721 12291
rect 4721 12257 4755 12291
rect 4755 12257 4764 12291
rect 4712 12248 4764 12257
rect 6368 12248 6420 12300
rect 7196 12248 7248 12300
rect 9772 12316 9824 12368
rect 10876 12316 10928 12368
rect 11060 12316 11112 12368
rect 7932 12248 7984 12300
rect 8576 12248 8628 12300
rect 9404 12291 9456 12300
rect 9404 12257 9413 12291
rect 9413 12257 9447 12291
rect 9447 12257 9456 12291
rect 9404 12248 9456 12257
rect 3240 12180 3292 12232
rect 4160 12180 4212 12232
rect 4896 12223 4948 12232
rect 4896 12189 4905 12223
rect 4905 12189 4939 12223
rect 4939 12189 4948 12223
rect 4896 12180 4948 12189
rect 5080 12112 5132 12164
rect 2872 12044 2924 12096
rect 4344 12087 4396 12096
rect 4344 12053 4353 12087
rect 4353 12053 4387 12087
rect 4387 12053 4396 12087
rect 4344 12044 4396 12053
rect 4712 12044 4764 12096
rect 5172 12044 5224 12096
rect 6552 12180 6604 12232
rect 6736 12180 6788 12232
rect 6920 12155 6972 12164
rect 6920 12121 6929 12155
rect 6929 12121 6963 12155
rect 6963 12121 6972 12155
rect 6920 12112 6972 12121
rect 6644 12044 6696 12096
rect 6828 12044 6880 12096
rect 9496 12180 9548 12232
rect 9956 12180 10008 12232
rect 11704 12248 11756 12300
rect 11888 12248 11940 12300
rect 8668 12112 8720 12164
rect 9864 12112 9916 12164
rect 9128 12044 9180 12096
rect 9772 12044 9824 12096
rect 10232 12044 10284 12096
rect 10416 12180 10468 12232
rect 10508 12112 10560 12164
rect 10784 12112 10836 12164
rect 10968 12180 11020 12232
rect 11520 12180 11572 12232
rect 11612 12112 11664 12164
rect 15384 12180 15436 12232
rect 11520 12044 11572 12096
rect 12440 12044 12492 12096
rect 13084 12112 13136 12164
rect 12808 12044 12860 12096
rect 14096 12044 14148 12096
rect 3447 11942 3499 11994
rect 3511 11942 3563 11994
rect 3575 11942 3627 11994
rect 3639 11942 3691 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 13308 11942 13360 11994
rect 13372 11942 13424 11994
rect 13436 11942 13488 11994
rect 13500 11942 13552 11994
rect 1768 11840 1820 11892
rect 2964 11840 3016 11892
rect 3148 11840 3200 11892
rect 3332 11840 3384 11892
rect 3792 11704 3844 11756
rect 5632 11840 5684 11892
rect 6552 11840 6604 11892
rect 10232 11840 10284 11892
rect 4436 11772 4488 11824
rect 8576 11772 8628 11824
rect 9036 11772 9088 11824
rect 11704 11840 11756 11892
rect 12900 11840 12952 11892
rect 4344 11747 4396 11756
rect 4344 11713 4353 11747
rect 4353 11713 4387 11747
rect 4387 11713 4396 11747
rect 4344 11704 4396 11713
rect 6828 11704 6880 11756
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 8484 11704 8536 11756
rect 8852 11704 8904 11756
rect 1676 11636 1728 11688
rect 2872 11679 2924 11688
rect 2872 11645 2881 11679
rect 2881 11645 2915 11679
rect 2915 11645 2924 11679
rect 2872 11636 2924 11645
rect 4896 11679 4948 11688
rect 4896 11645 4905 11679
rect 4905 11645 4939 11679
rect 4939 11645 4948 11679
rect 4896 11636 4948 11645
rect 5540 11636 5592 11688
rect 8944 11636 8996 11688
rect 9588 11679 9640 11688
rect 9588 11645 9597 11679
rect 9597 11645 9631 11679
rect 9631 11645 9640 11679
rect 9588 11636 9640 11645
rect 4252 11568 4304 11620
rect 5172 11611 5224 11620
rect 5172 11577 5206 11611
rect 5206 11577 5224 11611
rect 5172 11568 5224 11577
rect 3148 11500 3200 11552
rect 7288 11568 7340 11620
rect 7564 11568 7616 11620
rect 9496 11568 9548 11620
rect 10048 11704 10100 11756
rect 10876 11772 10928 11824
rect 10600 11704 10652 11756
rect 10968 11568 11020 11620
rect 11336 11772 11388 11824
rect 11520 11772 11572 11824
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 15108 11704 15160 11756
rect 11244 11636 11296 11688
rect 11520 11636 11572 11688
rect 12532 11636 12584 11688
rect 13268 11636 13320 11688
rect 13728 11636 13780 11688
rect 13820 11636 13872 11688
rect 13912 11568 13964 11620
rect 16396 11568 16448 11620
rect 6920 11500 6972 11552
rect 8852 11500 8904 11552
rect 9220 11543 9272 11552
rect 9220 11509 9229 11543
rect 9229 11509 9263 11543
rect 9263 11509 9272 11543
rect 9220 11500 9272 11509
rect 9772 11500 9824 11552
rect 10232 11500 10284 11552
rect 10508 11500 10560 11552
rect 11244 11500 11296 11552
rect 12716 11500 12768 11552
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 6104 11398 6156 11450
rect 10843 11398 10895 11450
rect 10907 11398 10959 11450
rect 10971 11398 11023 11450
rect 11035 11398 11087 11450
rect 1400 11296 1452 11348
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 5356 11296 5408 11348
rect 5448 11296 5500 11348
rect 7840 11296 7892 11348
rect 8208 11296 8260 11348
rect 9496 11296 9548 11348
rect 9956 11296 10008 11348
rect 10416 11296 10468 11348
rect 10508 11296 10560 11348
rect 11336 11339 11388 11348
rect 11336 11305 11345 11339
rect 11345 11305 11379 11339
rect 11379 11305 11388 11339
rect 11336 11296 11388 11305
rect 11796 11296 11848 11348
rect 13636 11296 13688 11348
rect 4436 11228 4488 11280
rect 1584 11160 1636 11212
rect 1952 11203 2004 11212
rect 1952 11169 1961 11203
rect 1961 11169 1995 11203
rect 1995 11169 2004 11203
rect 1952 11160 2004 11169
rect 2412 11160 2464 11212
rect 4620 11160 4672 11212
rect 5816 11203 5868 11212
rect 1492 11092 1544 11144
rect 2872 11092 2924 11144
rect 4804 11092 4856 11144
rect 5264 11135 5316 11144
rect 2596 11024 2648 11076
rect 4436 11024 4488 11076
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 5264 11092 5316 11101
rect 5448 11092 5500 11144
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 5908 11160 5960 11212
rect 6920 11160 6972 11212
rect 7472 11160 7524 11212
rect 9220 11228 9272 11280
rect 7380 11092 7432 11144
rect 8852 11092 8904 11144
rect 9220 11092 9272 11144
rect 10968 11160 11020 11212
rect 11060 11160 11112 11212
rect 11704 11228 11756 11280
rect 12624 11228 12676 11280
rect 12716 11228 12768 11280
rect 13176 11228 13228 11280
rect 13728 11228 13780 11280
rect 13084 11160 13136 11212
rect 10600 11092 10652 11144
rect 11796 11092 11848 11144
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 5816 11024 5868 11076
rect 9312 11024 9364 11076
rect 10968 11024 11020 11076
rect 11612 11024 11664 11076
rect 12900 11024 12952 11076
rect 13544 11024 13596 11076
rect 14372 11024 14424 11076
rect 2688 10956 2740 11008
rect 7012 10956 7064 11008
rect 7196 10999 7248 11008
rect 7196 10965 7205 10999
rect 7205 10965 7239 10999
rect 7239 10965 7248 10999
rect 7196 10956 7248 10965
rect 7288 10956 7340 11008
rect 11704 10956 11756 11008
rect 12440 10956 12492 11008
rect 12624 10956 12676 11008
rect 3447 10854 3499 10906
rect 3511 10854 3563 10906
rect 3575 10854 3627 10906
rect 3639 10854 3691 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 13308 10854 13360 10906
rect 13372 10854 13424 10906
rect 13436 10854 13488 10906
rect 13500 10854 13552 10906
rect 3240 10752 3292 10804
rect 2504 10684 2556 10736
rect 3056 10684 3108 10736
rect 2136 10616 2188 10668
rect 5172 10752 5224 10804
rect 5632 10752 5684 10804
rect 6460 10752 6512 10804
rect 7288 10752 7340 10804
rect 7564 10752 7616 10804
rect 9404 10752 9456 10804
rect 11060 10752 11112 10804
rect 4804 10616 4856 10668
rect 15200 10752 15252 10804
rect 11704 10727 11756 10736
rect 7472 10659 7524 10668
rect 1860 10523 1912 10532
rect 1860 10489 1869 10523
rect 1869 10489 1903 10523
rect 1903 10489 1912 10523
rect 1860 10480 1912 10489
rect 4896 10591 4948 10600
rect 2596 10480 2648 10532
rect 4620 10480 4672 10532
rect 4896 10557 4905 10591
rect 4905 10557 4939 10591
rect 4939 10557 4948 10591
rect 4896 10548 4948 10557
rect 5540 10548 5592 10600
rect 5080 10480 5132 10532
rect 5448 10480 5500 10532
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 7012 10548 7064 10600
rect 7380 10548 7432 10600
rect 8208 10591 8260 10600
rect 8208 10557 8217 10591
rect 8217 10557 8251 10591
rect 8251 10557 8260 10591
rect 8208 10548 8260 10557
rect 10784 10616 10836 10668
rect 10968 10659 11020 10668
rect 10968 10625 10977 10659
rect 10977 10625 11011 10659
rect 11011 10625 11020 10659
rect 10968 10616 11020 10625
rect 11704 10693 11713 10727
rect 11713 10693 11747 10727
rect 11747 10693 11756 10727
rect 11704 10684 11756 10693
rect 11612 10616 11664 10668
rect 13084 10616 13136 10668
rect 11704 10548 11756 10600
rect 2780 10412 2832 10464
rect 9312 10480 9364 10532
rect 7104 10412 7156 10464
rect 8852 10412 8904 10464
rect 10416 10412 10468 10464
rect 10508 10412 10560 10464
rect 12348 10480 12400 10532
rect 13084 10480 13136 10532
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 13820 10684 13872 10736
rect 13820 10548 13872 10600
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14004 10548 14056 10557
rect 16764 10548 16816 10600
rect 12440 10412 12492 10421
rect 14188 10412 14240 10464
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 6104 10310 6156 10362
rect 10843 10310 10895 10362
rect 10907 10310 10959 10362
rect 10971 10310 11023 10362
rect 11035 10310 11087 10362
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 2780 10208 2832 10217
rect 3240 10208 3292 10260
rect 3976 10208 4028 10260
rect 4252 10251 4304 10260
rect 4252 10217 4261 10251
rect 4261 10217 4295 10251
rect 4295 10217 4304 10251
rect 4252 10208 4304 10217
rect 4344 10208 4396 10260
rect 4896 10208 4948 10260
rect 5448 10208 5500 10260
rect 4436 10140 4488 10192
rect 4620 10183 4672 10192
rect 4620 10149 4629 10183
rect 4629 10149 4663 10183
rect 4663 10149 4672 10183
rect 4620 10140 4672 10149
rect 4804 10140 4856 10192
rect 7196 10208 7248 10260
rect 8024 10208 8076 10260
rect 11428 10208 11480 10260
rect 12072 10208 12124 10260
rect 2780 10072 2832 10124
rect 6828 10072 6880 10124
rect 7380 10072 7432 10124
rect 7564 10115 7616 10124
rect 7564 10081 7598 10115
rect 7598 10081 7616 10115
rect 7564 10072 7616 10081
rect 8024 10072 8076 10124
rect 9312 10115 9364 10124
rect 9312 10081 9321 10115
rect 9321 10081 9355 10115
rect 9355 10081 9364 10115
rect 9312 10072 9364 10081
rect 9772 10140 9824 10192
rect 10232 10140 10284 10192
rect 10416 10140 10468 10192
rect 10692 10140 10744 10192
rect 12900 10140 12952 10192
rect 13728 10208 13780 10260
rect 15568 10140 15620 10192
rect 3884 10004 3936 10056
rect 5080 10004 5132 10056
rect 2596 9868 2648 9920
rect 5264 9936 5316 9988
rect 5080 9868 5132 9920
rect 5448 10047 5500 10056
rect 5448 10013 5457 10047
rect 5457 10013 5491 10047
rect 5491 10013 5500 10047
rect 11244 10072 11296 10124
rect 5448 10004 5500 10013
rect 7656 9868 7708 9920
rect 9496 9936 9548 9988
rect 11060 10004 11112 10056
rect 11704 10072 11756 10124
rect 13912 10072 13964 10124
rect 14556 10072 14608 10124
rect 14648 10072 14700 10124
rect 14924 10072 14976 10124
rect 10416 9936 10468 9988
rect 11612 10004 11664 10056
rect 12072 10004 12124 10056
rect 12624 10004 12676 10056
rect 12900 10004 12952 10056
rect 13820 10047 13872 10056
rect 13820 10013 13829 10047
rect 13829 10013 13863 10047
rect 13863 10013 13872 10047
rect 13820 10004 13872 10013
rect 15476 10004 15528 10056
rect 14648 9979 14700 9988
rect 9404 9868 9456 9920
rect 11704 9868 11756 9920
rect 14648 9945 14657 9979
rect 14657 9945 14691 9979
rect 14691 9945 14700 9979
rect 14648 9936 14700 9945
rect 15292 9868 15344 9920
rect 3447 9766 3499 9818
rect 3511 9766 3563 9818
rect 3575 9766 3627 9818
rect 3639 9766 3691 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 13308 9766 13360 9818
rect 13372 9766 13424 9818
rect 13436 9766 13488 9818
rect 13500 9766 13552 9818
rect 2136 9639 2188 9648
rect 2136 9605 2145 9639
rect 2145 9605 2179 9639
rect 2179 9605 2188 9639
rect 2136 9596 2188 9605
rect 3700 9596 3752 9648
rect 2596 9571 2648 9580
rect 2596 9537 2605 9571
rect 2605 9537 2639 9571
rect 2639 9537 2648 9571
rect 2596 9528 2648 9537
rect 4896 9664 4948 9716
rect 5172 9707 5224 9716
rect 5172 9673 5181 9707
rect 5181 9673 5215 9707
rect 5215 9673 5224 9707
rect 5172 9664 5224 9673
rect 5264 9664 5316 9716
rect 9220 9664 9272 9716
rect 9404 9664 9456 9716
rect 10232 9664 10284 9716
rect 11336 9664 11388 9716
rect 11612 9664 11664 9716
rect 12164 9664 12216 9716
rect 13820 9664 13872 9716
rect 14004 9664 14056 9716
rect 14188 9664 14240 9716
rect 2872 9460 2924 9512
rect 2964 9460 3016 9512
rect 3332 9460 3384 9512
rect 2504 9435 2556 9444
rect 2504 9401 2513 9435
rect 2513 9401 2547 9435
rect 2547 9401 2556 9435
rect 2504 9392 2556 9401
rect 4896 9528 4948 9580
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 8116 9528 8168 9580
rect 9220 9528 9272 9580
rect 9404 9528 9456 9580
rect 3884 9392 3936 9444
rect 5540 9435 5592 9444
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 5172 9324 5224 9376
rect 5540 9401 5574 9435
rect 5574 9401 5592 9435
rect 5540 9392 5592 9401
rect 5816 9460 5868 9512
rect 8208 9460 8260 9512
rect 6276 9392 6328 9444
rect 7840 9392 7892 9444
rect 8300 9392 8352 9444
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 12348 9596 12400 9648
rect 12716 9596 12768 9648
rect 12808 9596 12860 9648
rect 13728 9596 13780 9648
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 10600 9528 10652 9580
rect 12624 9528 12676 9580
rect 9128 9460 9180 9469
rect 11152 9460 11204 9512
rect 11428 9460 11480 9512
rect 12256 9460 12308 9512
rect 12716 9460 12768 9512
rect 10692 9392 10744 9444
rect 12808 9435 12860 9444
rect 12808 9401 12817 9435
rect 12817 9401 12851 9435
rect 12851 9401 12860 9435
rect 12808 9392 12860 9401
rect 13084 9528 13136 9580
rect 13912 9460 13964 9512
rect 13084 9392 13136 9444
rect 6920 9324 6972 9376
rect 7564 9324 7616 9376
rect 9680 9324 9732 9376
rect 10324 9367 10376 9376
rect 10324 9333 10333 9367
rect 10333 9333 10367 9367
rect 10367 9333 10376 9367
rect 10324 9324 10376 9333
rect 11336 9324 11388 9376
rect 11520 9324 11572 9376
rect 11796 9324 11848 9376
rect 12256 9324 12308 9376
rect 14188 9324 14240 9376
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 6104 9222 6156 9274
rect 10843 9222 10895 9274
rect 10907 9222 10959 9274
rect 10971 9222 11023 9274
rect 11035 9222 11087 9274
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 3332 9120 3384 9172
rect 11336 9163 11388 9172
rect 11336 9129 11345 9163
rect 11345 9129 11379 9163
rect 11379 9129 11388 9163
rect 11336 9120 11388 9129
rect 13176 9120 13228 9172
rect 1308 9052 1360 9104
rect 5632 9052 5684 9104
rect 7564 9052 7616 9104
rect 7656 9052 7708 9104
rect 7840 9052 7892 9104
rect 8024 9052 8076 9104
rect 8392 9052 8444 9104
rect 2596 8984 2648 9036
rect 4620 9027 4672 9036
rect 1768 8916 1820 8968
rect 2688 8916 2740 8968
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 4804 8984 4856 9036
rect 5080 8984 5132 9036
rect 8668 9052 8720 9104
rect 8852 9052 8904 9104
rect 9128 9052 9180 9104
rect 10140 9095 10192 9104
rect 10140 9061 10149 9095
rect 10149 9061 10183 9095
rect 10183 9061 10192 9095
rect 10140 9052 10192 9061
rect 10324 9052 10376 9104
rect 14924 9120 14976 9172
rect 13820 9052 13872 9104
rect 4436 8916 4488 8968
rect 4528 8916 4580 8968
rect 4988 8916 5040 8968
rect 5172 8916 5224 8968
rect 8300 8959 8352 8968
rect 8300 8925 8309 8959
rect 8309 8925 8343 8959
rect 8343 8925 8352 8959
rect 8300 8916 8352 8925
rect 9404 8984 9456 9036
rect 9864 8984 9916 9036
rect 11244 9027 11296 9036
rect 3332 8848 3384 8900
rect 7472 8848 7524 8900
rect 7748 8891 7800 8900
rect 7748 8857 7757 8891
rect 7757 8857 7791 8891
rect 7791 8857 7800 8891
rect 7748 8848 7800 8857
rect 7840 8848 7892 8900
rect 9220 8916 9272 8968
rect 10416 8916 10468 8968
rect 11244 8993 11253 9027
rect 11253 8993 11287 9027
rect 11287 8993 11296 9027
rect 11244 8984 11296 8993
rect 12440 9027 12492 9036
rect 12440 8993 12449 9027
rect 12449 8993 12483 9027
rect 12483 8993 12492 9027
rect 12440 8984 12492 8993
rect 13176 8984 13228 9036
rect 14464 9027 14516 9036
rect 14464 8993 14473 9027
rect 14473 8993 14507 9027
rect 14507 8993 14516 9027
rect 14464 8984 14516 8993
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 12164 8916 12216 8968
rect 9496 8848 9548 8900
rect 1952 8780 2004 8832
rect 2320 8780 2372 8832
rect 2964 8780 3016 8832
rect 4252 8823 4304 8832
rect 4252 8789 4261 8823
rect 4261 8789 4295 8823
rect 4295 8789 4304 8823
rect 4252 8780 4304 8789
rect 4436 8780 4488 8832
rect 6920 8780 6972 8832
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 8852 8780 8904 8832
rect 9680 8823 9732 8832
rect 9680 8789 9689 8823
rect 9689 8789 9723 8823
rect 9723 8789 9732 8823
rect 9680 8780 9732 8789
rect 10784 8848 10836 8900
rect 12808 8916 12860 8968
rect 12992 8916 13044 8968
rect 13728 8916 13780 8968
rect 10600 8780 10652 8832
rect 10968 8780 11020 8832
rect 11704 8780 11756 8832
rect 12440 8780 12492 8832
rect 13820 8780 13872 8832
rect 3447 8678 3499 8730
rect 3511 8678 3563 8730
rect 3575 8678 3627 8730
rect 3639 8678 3691 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 13308 8678 13360 8730
rect 13372 8678 13424 8730
rect 13436 8678 13488 8730
rect 13500 8678 13552 8730
rect 2412 8576 2464 8628
rect 4068 8576 4120 8628
rect 9588 8576 9640 8628
rect 9864 8576 9916 8628
rect 11244 8576 11296 8628
rect 13636 8619 13688 8628
rect 13636 8585 13645 8619
rect 13645 8585 13679 8619
rect 13679 8585 13688 8619
rect 13636 8576 13688 8585
rect 4620 8508 4672 8560
rect 6276 8551 6328 8560
rect 6276 8517 6285 8551
rect 6285 8517 6319 8551
rect 6319 8517 6328 8551
rect 6276 8508 6328 8517
rect 7840 8508 7892 8560
rect 9496 8508 9548 8560
rect 11428 8508 11480 8560
rect 3608 8440 3660 8492
rect 3884 8372 3936 8424
rect 4068 8415 4120 8424
rect 4068 8381 4077 8415
rect 4077 8381 4111 8415
rect 4111 8381 4120 8415
rect 4068 8372 4120 8381
rect 4620 8372 4672 8424
rect 4804 8372 4856 8424
rect 8116 8440 8168 8492
rect 9404 8440 9456 8492
rect 10048 8440 10100 8492
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 11244 8440 11296 8492
rect 12164 8508 12216 8560
rect 12624 8440 12676 8492
rect 12808 8440 12860 8492
rect 13360 8508 13412 8560
rect 13728 8440 13780 8492
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 6276 8372 6328 8424
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 6920 8372 6972 8424
rect 9220 8372 9272 8424
rect 10232 8415 10284 8424
rect 10232 8381 10241 8415
rect 10241 8381 10275 8415
rect 10275 8381 10284 8415
rect 10232 8372 10284 8381
rect 1216 8304 1268 8356
rect 4344 8304 4396 8356
rect 1124 8236 1176 8288
rect 1584 8236 1636 8288
rect 2320 8236 2372 8288
rect 2688 8236 2740 8288
rect 3700 8236 3752 8288
rect 3884 8236 3936 8288
rect 4896 8236 4948 8288
rect 7196 8304 7248 8356
rect 7012 8236 7064 8288
rect 7380 8236 7432 8288
rect 8116 8236 8168 8288
rect 8300 8236 8352 8288
rect 9496 8304 9548 8356
rect 10784 8372 10836 8424
rect 10416 8304 10468 8356
rect 10968 8304 11020 8356
rect 11520 8304 11572 8356
rect 9404 8236 9456 8288
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 13452 8372 13504 8424
rect 12624 8304 12676 8356
rect 13912 8372 13964 8424
rect 14556 8372 14608 8424
rect 14924 8372 14976 8424
rect 13728 8304 13780 8356
rect 14280 8236 14332 8288
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 6104 8134 6156 8186
rect 10843 8134 10895 8186
rect 10907 8134 10959 8186
rect 10971 8134 11023 8186
rect 11035 8134 11087 8186
rect 1216 8032 1268 8084
rect 4252 8032 4304 8084
rect 4436 8032 4488 8084
rect 8300 8032 8352 8084
rect 8944 8032 8996 8084
rect 9588 8032 9640 8084
rect 9864 8032 9916 8084
rect 2688 7964 2740 8016
rect 11428 8032 11480 8084
rect 11520 8032 11572 8084
rect 13084 8032 13136 8084
rect 13360 8032 13412 8084
rect 13452 8032 13504 8084
rect 3884 7896 3936 7948
rect 4344 7939 4396 7948
rect 4344 7905 4378 7939
rect 4378 7905 4396 7939
rect 4344 7896 4396 7905
rect 4896 7896 4948 7948
rect 7840 7896 7892 7948
rect 3240 7871 3292 7880
rect 3240 7837 3249 7871
rect 3249 7837 3283 7871
rect 3283 7837 3292 7871
rect 3240 7828 3292 7837
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 3516 7760 3568 7812
rect 3884 7760 3936 7812
rect 2228 7692 2280 7744
rect 5448 7735 5500 7744
rect 5448 7701 5457 7735
rect 5457 7701 5491 7735
rect 5491 7701 5500 7735
rect 7104 7760 7156 7812
rect 5448 7692 5500 7701
rect 7564 7692 7616 7744
rect 7656 7692 7708 7744
rect 9128 7896 9180 7948
rect 9404 7896 9456 7948
rect 11704 7964 11756 8016
rect 8944 7828 8996 7880
rect 10968 7828 11020 7880
rect 11428 7871 11480 7880
rect 11428 7837 11437 7871
rect 11437 7837 11471 7871
rect 11471 7837 11480 7871
rect 11428 7828 11480 7837
rect 12072 7896 12124 7948
rect 12256 7896 12308 7948
rect 12440 7939 12492 7948
rect 12440 7905 12449 7939
rect 12449 7905 12483 7939
rect 12483 7905 12492 7939
rect 12440 7896 12492 7905
rect 12716 7964 12768 8016
rect 12532 7871 12584 7880
rect 12164 7760 12216 7812
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 12808 7828 12860 7880
rect 13176 7896 13228 7948
rect 14188 7828 14240 7880
rect 13452 7760 13504 7812
rect 13544 7760 13596 7812
rect 14924 7760 14976 7812
rect 9036 7692 9088 7744
rect 9680 7692 9732 7744
rect 10232 7692 10284 7744
rect 10600 7692 10652 7744
rect 11704 7692 11756 7744
rect 12256 7692 12308 7744
rect 12532 7692 12584 7744
rect 12808 7692 12860 7744
rect 13636 7692 13688 7744
rect 3447 7590 3499 7642
rect 3511 7590 3563 7642
rect 3575 7590 3627 7642
rect 3639 7590 3691 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 13308 7590 13360 7642
rect 13372 7590 13424 7642
rect 13436 7590 13488 7642
rect 13500 7590 13552 7642
rect 1676 7488 1728 7540
rect 1492 7352 1544 7404
rect 2320 7395 2372 7404
rect 2320 7361 2329 7395
rect 2329 7361 2363 7395
rect 2363 7361 2372 7395
rect 2320 7352 2372 7361
rect 4344 7488 4396 7540
rect 6276 7531 6328 7540
rect 6276 7497 6285 7531
rect 6285 7497 6319 7531
rect 6319 7497 6328 7531
rect 6276 7488 6328 7497
rect 4712 7420 4764 7472
rect 7472 7488 7524 7540
rect 7564 7488 7616 7540
rect 2228 7327 2280 7336
rect 2228 7293 2237 7327
rect 2237 7293 2271 7327
rect 2271 7293 2280 7327
rect 2228 7284 2280 7293
rect 3056 7327 3108 7336
rect 3056 7293 3065 7327
rect 3065 7293 3099 7327
rect 3099 7293 3108 7327
rect 3056 7284 3108 7293
rect 4068 7284 4120 7336
rect 4896 7327 4948 7336
rect 4896 7293 4905 7327
rect 4905 7293 4939 7327
rect 4939 7293 4948 7327
rect 4896 7284 4948 7293
rect 8116 7420 8168 7472
rect 9864 7420 9916 7472
rect 6276 7352 6328 7404
rect 6000 7284 6052 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 8484 7352 8536 7404
rect 10140 7352 10192 7404
rect 10416 7352 10468 7404
rect 1492 7148 1544 7200
rect 3884 7148 3936 7200
rect 6276 7148 6328 7200
rect 8576 7216 8628 7268
rect 9496 7284 9548 7336
rect 10232 7284 10284 7336
rect 9036 7216 9088 7268
rect 9128 7216 9180 7268
rect 8208 7148 8260 7200
rect 9864 7148 9916 7200
rect 11060 7488 11112 7540
rect 11336 7488 11388 7540
rect 11704 7488 11756 7540
rect 12992 7488 13044 7540
rect 10968 7420 11020 7472
rect 11152 7420 11204 7472
rect 12716 7420 12768 7472
rect 14004 7420 14056 7472
rect 11704 7352 11756 7404
rect 12072 7352 12124 7404
rect 12532 7352 12584 7404
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 14924 7284 14976 7336
rect 11152 7148 11204 7200
rect 12348 7148 12400 7200
rect 12716 7148 12768 7200
rect 12900 7148 12952 7200
rect 13636 7191 13688 7200
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 14832 7148 14884 7200
rect 14924 7148 14976 7200
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 6104 7046 6156 7098
rect 10843 7046 10895 7098
rect 10907 7046 10959 7098
rect 10971 7046 11023 7098
rect 11035 7046 11087 7098
rect 7012 6944 7064 6996
rect 8392 6944 8444 6996
rect 8576 6944 8628 6996
rect 8944 6987 8996 6996
rect 8944 6953 8953 6987
rect 8953 6953 8987 6987
rect 8987 6953 8996 6987
rect 8944 6944 8996 6953
rect 9128 6944 9180 6996
rect 10048 6987 10100 6996
rect 10048 6953 10057 6987
rect 10057 6953 10091 6987
rect 10091 6953 10100 6987
rect 10048 6944 10100 6953
rect 2320 6876 2372 6928
rect 4344 6876 4396 6928
rect 9772 6876 9824 6928
rect 10140 6919 10192 6928
rect 10140 6885 10149 6919
rect 10149 6885 10183 6919
rect 10183 6885 10192 6919
rect 10140 6876 10192 6885
rect 10416 6944 10468 6996
rect 12256 6944 12308 6996
rect 12348 6944 12400 6996
rect 12808 6944 12860 6996
rect 11612 6876 11664 6928
rect 13728 6876 13780 6928
rect 1492 6740 1544 6792
rect 1860 6740 1912 6792
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 3976 6808 4028 6860
rect 5080 6851 5132 6860
rect 5080 6817 5089 6851
rect 5089 6817 5123 6851
rect 5123 6817 5132 6851
rect 5080 6808 5132 6817
rect 7656 6808 7708 6860
rect 7840 6851 7892 6860
rect 7840 6817 7874 6851
rect 7874 6817 7892 6851
rect 7840 6808 7892 6817
rect 8392 6808 8444 6860
rect 8944 6808 8996 6860
rect 4712 6740 4764 6792
rect 4896 6740 4948 6792
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 9404 6740 9456 6792
rect 9680 6740 9732 6792
rect 8668 6672 8720 6724
rect 10416 6808 10468 6860
rect 10968 6808 11020 6860
rect 11704 6808 11756 6860
rect 14464 6851 14516 6860
rect 10140 6740 10192 6792
rect 10508 6740 10560 6792
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 11612 6740 11664 6792
rect 12808 6740 12860 6792
rect 14464 6817 14473 6851
rect 14473 6817 14507 6851
rect 14507 6817 14516 6851
rect 14464 6808 14516 6817
rect 14648 6808 14700 6860
rect 1492 6604 1544 6656
rect 4712 6604 4764 6656
rect 5264 6604 5316 6656
rect 5448 6604 5500 6656
rect 9220 6604 9272 6656
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 11060 6672 11112 6724
rect 11152 6672 11204 6724
rect 9680 6604 9732 6613
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 3240 6400 3292 6452
rect 4160 6400 4212 6452
rect 2136 6332 2188 6384
rect 2228 6239 2280 6248
rect 2228 6205 2237 6239
rect 2237 6205 2271 6239
rect 2271 6205 2280 6239
rect 3056 6239 3108 6248
rect 2228 6196 2280 6205
rect 3056 6205 3065 6239
rect 3065 6205 3099 6239
rect 3099 6205 3108 6239
rect 3056 6196 3108 6205
rect 8208 6400 8260 6452
rect 9036 6400 9088 6452
rect 6276 6375 6328 6384
rect 6276 6341 6285 6375
rect 6285 6341 6319 6375
rect 6319 6341 6328 6375
rect 6276 6332 6328 6341
rect 9772 6400 9824 6452
rect 10324 6400 10376 6452
rect 12440 6443 12492 6452
rect 12440 6409 12449 6443
rect 12449 6409 12483 6443
rect 12483 6409 12492 6443
rect 12440 6400 12492 6409
rect 4896 6307 4948 6316
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 7840 6264 7892 6316
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 7564 6196 7616 6248
rect 10232 6264 10284 6316
rect 12532 6264 12584 6316
rect 12716 6332 12768 6384
rect 14280 6307 14332 6316
rect 14280 6273 14289 6307
rect 14289 6273 14323 6307
rect 14323 6273 14332 6307
rect 14280 6264 14332 6273
rect 10324 6196 10376 6248
rect 10600 6196 10652 6248
rect 10968 6239 11020 6248
rect 10968 6205 10977 6239
rect 10977 6205 11011 6239
rect 11011 6205 11020 6239
rect 10968 6196 11020 6205
rect 12440 6196 12492 6248
rect 13084 6196 13136 6248
rect 15476 6196 15528 6248
rect 5448 6128 5500 6180
rect 5540 6128 5592 6180
rect 6460 6128 6512 6180
rect 8116 6128 8168 6180
rect 9496 6128 9548 6180
rect 1308 6060 1360 6112
rect 3884 6060 3936 6112
rect 4160 6060 4212 6112
rect 7564 6060 7616 6112
rect 7656 6060 7708 6112
rect 8208 6103 8260 6112
rect 8208 6069 8217 6103
rect 8217 6069 8251 6103
rect 8251 6069 8260 6103
rect 8208 6060 8260 6069
rect 8576 6060 8628 6112
rect 10692 6060 10744 6112
rect 13360 6128 13412 6180
rect 15108 6128 15160 6180
rect 12716 6060 12768 6112
rect 13636 6103 13688 6112
rect 13636 6069 13645 6103
rect 13645 6069 13679 6103
rect 13679 6069 13688 6103
rect 13636 6060 13688 6069
rect 13820 6060 13872 6112
rect 14188 6060 14240 6112
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 2228 5788 2280 5840
rect 5540 5788 5592 5840
rect 5632 5788 5684 5840
rect 7288 5788 7340 5840
rect 8576 5788 8628 5840
rect 10048 5856 10100 5908
rect 11336 5856 11388 5908
rect 11888 5899 11940 5908
rect 11888 5865 11897 5899
rect 11897 5865 11931 5899
rect 11931 5865 11940 5899
rect 11888 5856 11940 5865
rect 12532 5856 12584 5908
rect 12716 5899 12768 5908
rect 12716 5865 12725 5899
rect 12725 5865 12759 5899
rect 12759 5865 12768 5899
rect 12716 5856 12768 5865
rect 12900 5856 12952 5908
rect 9772 5788 9824 5840
rect 2136 5763 2188 5772
rect 2136 5729 2145 5763
rect 2145 5729 2179 5763
rect 2179 5729 2188 5763
rect 2136 5720 2188 5729
rect 4620 5720 4672 5772
rect 5172 5652 5224 5704
rect 6736 5720 6788 5772
rect 7196 5720 7248 5772
rect 8852 5720 8904 5772
rect 6828 5652 6880 5704
rect 3884 5584 3936 5636
rect 5080 5584 5132 5636
rect 8300 5584 8352 5636
rect 8852 5584 8904 5636
rect 9312 5584 9364 5636
rect 1400 5516 1452 5568
rect 1860 5516 1912 5568
rect 2412 5516 2464 5568
rect 4068 5516 4120 5568
rect 5448 5516 5500 5568
rect 7564 5516 7616 5568
rect 10508 5720 10560 5772
rect 11060 5788 11112 5840
rect 12164 5788 12216 5840
rect 10784 5720 10836 5772
rect 11612 5720 11664 5772
rect 12440 5720 12492 5772
rect 13912 5720 13964 5772
rect 12164 5695 12216 5704
rect 11060 5627 11112 5636
rect 11060 5593 11069 5627
rect 11069 5593 11103 5627
rect 11103 5593 11112 5627
rect 11060 5584 11112 5593
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 12992 5652 13044 5704
rect 13360 5652 13412 5704
rect 15108 5720 15160 5772
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 14188 5584 14240 5636
rect 10416 5516 10468 5568
rect 11152 5516 11204 5568
rect 13912 5559 13964 5568
rect 13912 5525 13921 5559
rect 13921 5525 13955 5559
rect 13955 5525 13964 5559
rect 13912 5516 13964 5525
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 3240 5312 3292 5364
rect 4344 5312 4396 5364
rect 3056 5244 3108 5296
rect 4620 5244 4672 5296
rect 6644 5244 6696 5296
rect 6828 5244 6880 5296
rect 8116 5312 8168 5364
rect 10232 5312 10284 5364
rect 11060 5312 11112 5364
rect 11520 5312 11572 5364
rect 11888 5312 11940 5364
rect 12348 5312 12400 5364
rect 13636 5355 13688 5364
rect 13636 5321 13645 5355
rect 13645 5321 13679 5355
rect 13679 5321 13688 5355
rect 13636 5312 13688 5321
rect 8668 5244 8720 5296
rect 11428 5244 11480 5296
rect 12624 5244 12676 5296
rect 2504 5219 2556 5228
rect 2504 5185 2513 5219
rect 2513 5185 2547 5219
rect 2547 5185 2556 5219
rect 2504 5176 2556 5185
rect 2320 5015 2372 5024
rect 2320 4981 2329 5015
rect 2329 4981 2363 5015
rect 2363 4981 2372 5015
rect 9956 5176 10008 5228
rect 10508 5176 10560 5228
rect 11060 5219 11112 5228
rect 4896 5151 4948 5160
rect 4896 5117 4905 5151
rect 4905 5117 4939 5151
rect 4939 5117 4948 5151
rect 4896 5108 4948 5117
rect 3424 5040 3476 5092
rect 5448 5108 5500 5160
rect 6736 5108 6788 5160
rect 6920 5108 6972 5160
rect 7104 5151 7156 5160
rect 7104 5117 7138 5151
rect 7138 5117 7156 5151
rect 7104 5108 7156 5117
rect 7656 5108 7708 5160
rect 8944 5151 8996 5160
rect 8944 5117 8978 5151
rect 8978 5117 8996 5151
rect 8944 5108 8996 5117
rect 10600 5108 10652 5160
rect 11060 5185 11069 5219
rect 11069 5185 11103 5219
rect 11103 5185 11112 5219
rect 11060 5176 11112 5185
rect 12164 5176 12216 5228
rect 12992 5219 13044 5228
rect 12992 5185 13001 5219
rect 13001 5185 13035 5219
rect 13035 5185 13044 5219
rect 12992 5176 13044 5185
rect 13452 5219 13504 5228
rect 13452 5185 13461 5219
rect 13461 5185 13495 5219
rect 13495 5185 13504 5219
rect 14188 5219 14240 5228
rect 13452 5176 13504 5185
rect 11244 5108 11296 5160
rect 11612 5108 11664 5160
rect 13820 5108 13872 5160
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 14924 5108 14976 5160
rect 5632 5040 5684 5092
rect 8116 5040 8168 5092
rect 9128 5040 9180 5092
rect 9496 5040 9548 5092
rect 10968 5083 11020 5092
rect 6276 5015 6328 5024
rect 2320 4972 2372 4981
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 6920 4972 6972 5024
rect 8576 4972 8628 5024
rect 9220 4972 9272 5024
rect 9312 4972 9364 5024
rect 10048 4972 10100 5024
rect 10140 4972 10192 5024
rect 10968 5049 10977 5083
rect 10977 5049 11011 5083
rect 11011 5049 11020 5083
rect 10968 5040 11020 5049
rect 11796 5040 11848 5092
rect 13268 5040 13320 5092
rect 13636 5040 13688 5092
rect 12440 4972 12492 5024
rect 13820 4972 13872 5024
rect 14648 4972 14700 5024
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 3056 4768 3108 4820
rect 10048 4811 10100 4820
rect 2412 4743 2464 4752
rect 2412 4709 2446 4743
rect 2446 4709 2464 4743
rect 2412 4700 2464 4709
rect 2688 4700 2740 4752
rect 4344 4700 4396 4752
rect 6828 4700 6880 4752
rect 7012 4700 7064 4752
rect 7656 4700 7708 4752
rect 7748 4700 7800 4752
rect 8852 4700 8904 4752
rect 9404 4700 9456 4752
rect 1860 4632 1912 4684
rect 2872 4632 2924 4684
rect 2964 4632 3016 4684
rect 3792 4632 3844 4684
rect 5356 4632 5408 4684
rect 5540 4675 5592 4684
rect 5540 4641 5574 4675
rect 5574 4641 5592 4675
rect 5540 4632 5592 4641
rect 7380 4675 7432 4684
rect 7380 4641 7414 4675
rect 7414 4641 7432 4675
rect 7380 4632 7432 4641
rect 8208 4632 8260 4684
rect 9588 4700 9640 4752
rect 10048 4777 10057 4811
rect 10057 4777 10091 4811
rect 10091 4777 10100 4811
rect 10048 4768 10100 4777
rect 11244 4768 11296 4820
rect 11336 4768 11388 4820
rect 9956 4700 10008 4752
rect 11060 4700 11112 4752
rect 11888 4700 11940 4752
rect 12440 4743 12492 4752
rect 12440 4709 12449 4743
rect 12449 4709 12483 4743
rect 12483 4709 12492 4743
rect 12440 4700 12492 4709
rect 12716 4700 12768 4752
rect 13176 4768 13228 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 4620 4496 4672 4548
rect 2412 4428 2464 4480
rect 4344 4428 4396 4480
rect 5080 4564 5132 4616
rect 6736 4564 6788 4616
rect 8852 4564 8904 4616
rect 10968 4632 11020 4684
rect 11244 4675 11296 4684
rect 11244 4641 11253 4675
rect 11253 4641 11287 4675
rect 11287 4641 11296 4675
rect 11244 4632 11296 4641
rect 11520 4632 11572 4684
rect 11796 4632 11848 4684
rect 9864 4564 9916 4616
rect 10048 4564 10100 4616
rect 10784 4564 10836 4616
rect 11612 4564 11664 4616
rect 11704 4564 11756 4616
rect 8300 4496 8352 4548
rect 8484 4539 8536 4548
rect 8484 4505 8493 4539
rect 8493 4505 8527 4539
rect 8527 4505 8536 4539
rect 8484 4496 8536 4505
rect 8668 4496 8720 4548
rect 12992 4496 13044 4548
rect 14188 4564 14240 4616
rect 14648 4539 14700 4548
rect 14648 4505 14657 4539
rect 14657 4505 14691 4539
rect 14691 4505 14700 4539
rect 14648 4496 14700 4505
rect 5080 4428 5132 4480
rect 7380 4428 7432 4480
rect 7472 4428 7524 4480
rect 9680 4471 9732 4480
rect 9680 4437 9689 4471
rect 9689 4437 9723 4471
rect 9723 4437 9732 4471
rect 9680 4428 9732 4437
rect 10324 4428 10376 4480
rect 10968 4428 11020 4480
rect 11888 4428 11940 4480
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 2872 4224 2924 4276
rect 2504 4131 2556 4140
rect 2504 4097 2513 4131
rect 2513 4097 2547 4131
rect 2547 4097 2556 4131
rect 2504 4088 2556 4097
rect 4896 4224 4948 4276
rect 5080 4224 5132 4276
rect 7012 4224 7064 4276
rect 7104 4224 7156 4276
rect 4252 4156 4304 4208
rect 4620 4156 4672 4208
rect 7840 4224 7892 4276
rect 9220 4224 9272 4276
rect 9312 4224 9364 4276
rect 10232 4224 10284 4276
rect 11244 4224 11296 4276
rect 11428 4224 11480 4276
rect 4160 4088 4212 4140
rect 8116 4156 8168 4208
rect 8576 4156 8628 4208
rect 9312 4131 9364 4140
rect 4896 4063 4948 4072
rect 4252 3952 4304 4004
rect 2136 3884 2188 3936
rect 4160 3884 4212 3936
rect 4896 4029 4905 4063
rect 4905 4029 4939 4063
rect 4939 4029 4948 4063
rect 4896 4020 4948 4029
rect 6736 4020 6788 4072
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 5172 3995 5224 4004
rect 5172 3961 5206 3995
rect 5206 3961 5224 3995
rect 8668 4020 8720 4072
rect 9772 4156 9824 4208
rect 12164 4224 12216 4276
rect 13636 4224 13688 4276
rect 10048 4088 10100 4140
rect 11336 4088 11388 4140
rect 11888 4088 11940 4140
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 13084 4088 13136 4140
rect 14464 4156 14516 4208
rect 10232 4063 10284 4072
rect 5172 3952 5224 3961
rect 5448 3884 5500 3936
rect 5540 3884 5592 3936
rect 6920 3952 6972 4004
rect 7012 3952 7064 4004
rect 7472 3952 7524 4004
rect 8116 3952 8168 4004
rect 8484 3952 8536 4004
rect 9680 3952 9732 4004
rect 10232 4029 10241 4063
rect 10241 4029 10275 4063
rect 10275 4029 10284 4063
rect 10232 4020 10284 4029
rect 10692 4020 10744 4072
rect 12440 4020 12492 4072
rect 13268 4020 13320 4072
rect 15200 4020 15252 4072
rect 10784 3952 10836 4004
rect 11060 3952 11112 4004
rect 9036 3927 9088 3936
rect 9036 3893 9045 3927
rect 9045 3893 9079 3927
rect 9079 3893 9088 3927
rect 9036 3884 9088 3893
rect 9220 3884 9272 3936
rect 9496 3884 9548 3936
rect 10048 3884 10100 3936
rect 11244 3884 11296 3936
rect 11612 3952 11664 4004
rect 11796 3884 11848 3936
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 13268 3884 13320 3936
rect 14464 3884 14516 3936
rect 14648 3884 14700 3936
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 1952 3723 2004 3732
rect 1952 3689 1961 3723
rect 1961 3689 1995 3723
rect 1995 3689 2004 3723
rect 1952 3680 2004 3689
rect 2136 3680 2188 3732
rect 3240 3723 3292 3732
rect 3240 3689 3249 3723
rect 3249 3689 3283 3723
rect 3283 3689 3292 3723
rect 3240 3680 3292 3689
rect 4252 3680 4304 3732
rect 4436 3680 4488 3732
rect 4988 3723 5040 3732
rect 4988 3689 4997 3723
rect 4997 3689 5031 3723
rect 5031 3689 5040 3723
rect 4988 3680 5040 3689
rect 5448 3680 5500 3732
rect 2688 3612 2740 3664
rect 8484 3612 8536 3664
rect 8852 3680 8904 3732
rect 9680 3680 9732 3732
rect 9956 3680 10008 3732
rect 11244 3723 11296 3732
rect 11244 3689 11253 3723
rect 11253 3689 11287 3723
rect 11287 3689 11296 3723
rect 11244 3680 11296 3689
rect 12072 3723 12124 3732
rect 12072 3689 12081 3723
rect 12081 3689 12115 3723
rect 12115 3689 12124 3723
rect 12072 3680 12124 3689
rect 13268 3680 13320 3732
rect 13636 3723 13688 3732
rect 13636 3689 13645 3723
rect 13645 3689 13679 3723
rect 13679 3689 13688 3723
rect 13636 3680 13688 3689
rect 3240 3476 3292 3528
rect 6276 3544 6328 3596
rect 6736 3544 6788 3596
rect 6920 3544 6972 3596
rect 7564 3587 7616 3596
rect 7564 3553 7573 3587
rect 7573 3553 7607 3587
rect 7607 3553 7616 3587
rect 7564 3544 7616 3553
rect 7656 3544 7708 3596
rect 9128 3544 9180 3596
rect 9496 3544 9548 3596
rect 13912 3680 13964 3732
rect 13820 3612 13872 3664
rect 14188 3612 14240 3664
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 5448 3476 5500 3528
rect 2780 3451 2832 3460
rect 2780 3417 2789 3451
rect 2789 3417 2823 3451
rect 2823 3417 2832 3451
rect 2780 3408 2832 3417
rect 3148 3408 3200 3460
rect 5632 3408 5684 3460
rect 6828 3408 6880 3460
rect 756 3340 808 3392
rect 1492 3340 1544 3392
rect 4160 3340 4212 3392
rect 7104 3383 7156 3392
rect 7104 3349 7113 3383
rect 7113 3349 7147 3383
rect 7147 3349 7156 3383
rect 7104 3340 7156 3349
rect 10048 3476 10100 3528
rect 10416 3544 10468 3596
rect 11152 3544 11204 3596
rect 11244 3544 11296 3596
rect 14096 3544 14148 3596
rect 10784 3476 10836 3528
rect 10876 3476 10928 3528
rect 11704 3476 11756 3528
rect 11888 3476 11940 3528
rect 9220 3340 9272 3392
rect 10692 3408 10744 3460
rect 10048 3340 10100 3392
rect 11428 3340 11480 3392
rect 12256 3408 12308 3460
rect 13268 3451 13320 3460
rect 13268 3417 13277 3451
rect 13277 3417 13311 3451
rect 13311 3417 13320 3451
rect 13268 3408 13320 3417
rect 13820 3408 13872 3460
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 2320 3136 2372 3188
rect 4252 3136 4304 3188
rect 3240 3068 3292 3120
rect 1124 3000 1176 3052
rect 2504 3000 2556 3052
rect 3148 3043 3200 3052
rect 3148 3009 3157 3043
rect 3157 3009 3191 3043
rect 3191 3009 3200 3043
rect 3148 3000 3200 3009
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 4068 2975 4120 2984
rect 4068 2941 4077 2975
rect 4077 2941 4111 2975
rect 4111 2941 4120 2975
rect 4068 2932 4120 2941
rect 5540 3136 5592 3188
rect 7196 3136 7248 3188
rect 8116 3136 8168 3188
rect 4896 3068 4948 3120
rect 4436 3000 4488 3052
rect 4620 3000 4672 3052
rect 6276 3000 6328 3052
rect 6552 3000 6604 3052
rect 6736 3000 6788 3052
rect 5632 2932 5684 2984
rect 388 2796 440 2848
rect 1400 2796 1452 2848
rect 3056 2796 3108 2848
rect 5724 2864 5776 2916
rect 6368 2864 6420 2916
rect 5540 2796 5592 2848
rect 5632 2796 5684 2848
rect 7564 2932 7616 2984
rect 13084 3136 13136 3188
rect 13728 3136 13780 3188
rect 8668 3111 8720 3120
rect 8668 3077 8677 3111
rect 8677 3077 8711 3111
rect 8711 3077 8720 3111
rect 8668 3068 8720 3077
rect 9772 3111 9824 3120
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 9772 3077 9781 3111
rect 9781 3077 9815 3111
rect 9815 3077 9824 3111
rect 9772 3068 9824 3077
rect 10048 3068 10100 3120
rect 10416 3000 10468 3052
rect 10784 3068 10836 3120
rect 11796 3068 11848 3120
rect 10968 3000 11020 3052
rect 13820 3000 13872 3052
rect 14096 3043 14148 3052
rect 14096 3009 14105 3043
rect 14105 3009 14139 3043
rect 14139 3009 14148 3043
rect 14096 3000 14148 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 8392 2932 8444 2984
rect 10048 2932 10100 2984
rect 7012 2864 7064 2916
rect 7196 2864 7248 2916
rect 7840 2864 7892 2916
rect 8116 2864 8168 2916
rect 9220 2864 9272 2916
rect 11520 2932 11572 2984
rect 11796 2932 11848 2984
rect 10968 2864 11020 2916
rect 8852 2796 8904 2848
rect 8944 2796 8996 2848
rect 9864 2839 9916 2848
rect 9864 2805 9873 2839
rect 9873 2805 9907 2839
rect 9907 2805 9916 2839
rect 9864 2796 9916 2805
rect 10048 2796 10100 2848
rect 12992 2864 13044 2916
rect 13912 2932 13964 2984
rect 15108 2864 15160 2916
rect 11428 2839 11480 2848
rect 11428 2805 11437 2839
rect 11437 2805 11471 2839
rect 11471 2805 11480 2839
rect 11428 2796 11480 2805
rect 12440 2839 12492 2848
rect 12440 2805 12449 2839
rect 12449 2805 12483 2839
rect 12483 2805 12492 2839
rect 12900 2839 12952 2848
rect 12440 2796 12492 2805
rect 12900 2805 12909 2839
rect 12909 2805 12943 2839
rect 12943 2805 12952 2839
rect 12900 2796 12952 2805
rect 13636 2796 13688 2848
rect 14096 2796 14148 2848
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 5724 2592 5776 2644
rect 6460 2592 6512 2644
rect 8024 2592 8076 2644
rect 4436 2524 4488 2576
rect 5448 2524 5500 2576
rect 5540 2524 5592 2576
rect 9680 2592 9732 2644
rect 10140 2635 10192 2644
rect 10140 2601 10149 2635
rect 10149 2601 10183 2635
rect 10183 2601 10192 2635
rect 10140 2592 10192 2601
rect 10324 2592 10376 2644
rect 11428 2635 11480 2644
rect 11428 2601 11437 2635
rect 11437 2601 11471 2635
rect 11471 2601 11480 2635
rect 11428 2592 11480 2601
rect 12256 2592 12308 2644
rect 12440 2592 12492 2644
rect 14188 2592 14240 2644
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 2872 2456 2924 2508
rect 3976 2456 4028 2508
rect 4620 2456 4672 2508
rect 4344 2431 4396 2440
rect 112 2252 164 2304
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 7012 2252 7064 2304
rect 7656 2456 7708 2508
rect 9036 2456 9088 2508
rect 9496 2499 9548 2508
rect 9496 2465 9505 2499
rect 9505 2465 9539 2499
rect 9539 2465 9548 2499
rect 9496 2456 9548 2465
rect 10692 2524 10744 2576
rect 12164 2524 12216 2576
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 8116 2388 8168 2440
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 7380 2320 7432 2372
rect 9312 2388 9364 2440
rect 11336 2388 11388 2440
rect 10416 2320 10468 2372
rect 12716 2524 12768 2576
rect 12992 2567 13044 2576
rect 12992 2533 13001 2567
rect 13001 2533 13035 2567
rect 13035 2533 13044 2567
rect 12992 2524 13044 2533
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9772 2295 9824 2304
rect 9312 2252 9364 2261
rect 9772 2261 9781 2295
rect 9781 2261 9815 2295
rect 9815 2261 9824 2295
rect 9772 2252 9824 2261
rect 11336 2252 11388 2304
rect 12164 2295 12216 2304
rect 12164 2261 12173 2295
rect 12173 2261 12207 2295
rect 12207 2261 12216 2295
rect 12164 2252 12216 2261
rect 12256 2252 12308 2304
rect 12440 2456 12492 2508
rect 15292 2456 15344 2508
rect 13912 2388 13964 2440
rect 12440 2320 12492 2372
rect 12808 2320 12860 2372
rect 13728 2320 13780 2372
rect 14280 2320 14332 2372
rect 13820 2295 13872 2304
rect 13820 2261 13829 2295
rect 13829 2261 13863 2295
rect 13863 2261 13872 2295
rect 13820 2252 13872 2261
rect 13912 2252 13964 2304
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 7932 2048 7984 2100
rect 8944 2048 8996 2100
rect 10232 2048 10284 2100
rect 13912 2048 13964 2100
rect 8576 1980 8628 2032
rect 9128 1980 9180 2032
rect 9312 1980 9364 2032
rect 12256 1980 12308 2032
rect 12532 1980 12584 2032
rect 13360 1980 13412 2032
rect 4344 1912 4396 1964
rect 16028 1912 16080 1964
rect 6920 1844 6972 1896
rect 8116 1844 8168 1896
rect 10324 1844 10376 1896
rect 13636 1844 13688 1896
rect 2964 1776 3016 1828
rect 9312 1776 9364 1828
rect 9772 1776 9824 1828
rect 14832 1776 14884 1828
rect 1860 1708 1912 1760
rect 13820 1708 13872 1760
rect 1400 1640 1452 1692
rect 9036 1640 9088 1692
rect 4988 1572 5040 1624
rect 12164 1572 12216 1624
rect 8208 1504 8260 1556
rect 11428 1504 11480 1556
rect 3148 1232 3200 1284
rect 5080 1232 5132 1284
rect 3516 960 3568 1012
rect 7288 960 7340 1012
<< metal2 >>
rect 110 19520 166 20000
rect 386 19520 442 20000
rect 754 19520 810 20000
rect 1122 19520 1178 20000
rect 1398 19520 1454 20000
rect 1766 19520 1822 20000
rect 2134 19520 2190 20000
rect 2410 19520 2466 20000
rect 2778 19520 2834 20000
rect 3146 19520 3202 20000
rect 3514 19520 3570 20000
rect 3790 19520 3846 20000
rect 4158 19520 4214 20000
rect 4526 19520 4582 20000
rect 4802 19520 4858 20000
rect 5170 19520 5226 20000
rect 5538 19520 5594 20000
rect 5814 19520 5870 20000
rect 6182 19520 6238 20000
rect 6550 19520 6606 20000
rect 6918 19520 6974 20000
rect 7194 19520 7250 20000
rect 7562 19520 7618 20000
rect 7930 19520 7986 20000
rect 8206 19520 8262 20000
rect 8574 19520 8630 20000
rect 8942 19520 8998 20000
rect 9218 19520 9274 20000
rect 9586 19520 9642 20000
rect 9954 19520 10010 20000
rect 10322 19520 10378 20000
rect 10598 19520 10654 20000
rect 10966 19520 11022 20000
rect 11334 19530 11390 20000
rect 11334 19520 11468 19530
rect 11610 19520 11666 20000
rect 11978 19520 12034 20000
rect 12346 19520 12402 20000
rect 12622 19520 12678 20000
rect 12990 19520 13046 20000
rect 13358 19520 13414 20000
rect 13726 19520 13782 20000
rect 14002 19520 14058 20000
rect 14370 19520 14426 20000
rect 14738 19520 14794 20000
rect 15014 19520 15070 20000
rect 15382 19520 15438 20000
rect 15750 19520 15806 20000
rect 16026 19520 16082 20000
rect 16394 19520 16450 20000
rect 16762 19520 16818 20000
rect 124 16046 152 19520
rect 112 16040 164 16046
rect 112 15982 164 15988
rect 400 15978 428 19520
rect 768 17202 796 19520
rect 756 17196 808 17202
rect 756 17138 808 17144
rect 1136 16590 1164 19520
rect 1124 16584 1176 16590
rect 1124 16526 1176 16532
rect 1412 16114 1440 19520
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 1504 17134 1532 19343
rect 1674 18456 1730 18465
rect 1674 18391 1730 18400
rect 1492 17128 1544 17134
rect 1492 17070 1544 17076
rect 1688 16726 1716 18391
rect 1676 16720 1728 16726
rect 1676 16662 1728 16668
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1492 16584 1544 16590
rect 1492 16526 1544 16532
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 388 15972 440 15978
rect 388 15914 440 15920
rect 1320 15065 1348 15982
rect 1504 15688 1532 16526
rect 1596 16522 1624 16594
rect 1584 16516 1636 16522
rect 1584 16458 1636 16464
rect 1780 16114 1808 19520
rect 2148 17202 2176 19520
rect 2424 17270 2452 19520
rect 2412 17264 2464 17270
rect 2412 17206 2464 17212
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 1860 17060 1912 17066
rect 1860 17002 1912 17008
rect 1872 16250 1900 17002
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 1860 16244 1912 16250
rect 1860 16186 1912 16192
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 2412 16040 2464 16046
rect 2412 15982 2464 15988
rect 1412 15660 1532 15688
rect 1306 15056 1362 15065
rect 1306 14991 1362 15000
rect 1412 12889 1440 15660
rect 1492 15564 1544 15570
rect 1492 15506 1544 15512
rect 1398 12880 1454 12889
rect 1398 12815 1454 12824
rect 1412 11354 1440 12815
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1504 11234 1532 15506
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1596 11354 1624 13806
rect 1688 13530 1716 14214
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1780 11898 1808 14894
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1412 11206 1532 11234
rect 1584 11212 1636 11218
rect 1308 9104 1360 9110
rect 1308 9046 1360 9052
rect 1214 8392 1270 8401
rect 1214 8327 1216 8336
rect 1268 8327 1270 8336
rect 1216 8298 1268 8304
rect 1124 8288 1176 8294
rect 1124 8230 1176 8236
rect 1214 8256 1270 8265
rect 756 3392 808 3398
rect 756 3334 808 3340
rect 388 2848 440 2854
rect 388 2790 440 2796
rect 112 2304 164 2310
rect 112 2246 164 2252
rect 124 480 152 2246
rect 400 480 428 2790
rect 768 480 796 3334
rect 1136 3058 1164 8230
rect 1214 8191 1270 8200
rect 1228 8090 1256 8191
rect 1216 8084 1268 8090
rect 1216 8026 1268 8032
rect 1320 6118 1348 9046
rect 1412 7290 1440 11206
rect 1584 11154 1636 11160
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1504 7410 1532 11086
rect 1596 8294 1624 11154
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1582 8120 1638 8129
rect 1688 8106 1716 11630
rect 1872 10690 1900 14894
rect 1950 11248 2006 11257
rect 1950 11183 1952 11192
rect 2004 11183 2006 11192
rect 1952 11154 2004 11160
rect 1780 10662 1900 10690
rect 1780 10282 1808 10662
rect 1860 10532 1912 10538
rect 1860 10474 1912 10480
rect 1872 10441 1900 10474
rect 1858 10432 1914 10441
rect 1858 10367 1914 10376
rect 1780 10254 1900 10282
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1780 8129 1808 8910
rect 1638 8078 1716 8106
rect 1766 8120 1822 8129
rect 1582 8055 1638 8064
rect 1766 8055 1822 8064
rect 1582 7984 1638 7993
rect 1766 7984 1822 7993
rect 1638 7942 1716 7970
rect 1582 7919 1638 7928
rect 1688 7546 1716 7942
rect 1766 7919 1822 7928
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1412 7262 1624 7290
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6798 1532 7142
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1308 6112 1360 6118
rect 1308 6054 1360 6060
rect 1400 5568 1452 5574
rect 1400 5510 1452 5516
rect 1124 3052 1176 3058
rect 1124 2994 1176 3000
rect 1122 2952 1178 2961
rect 1122 2887 1178 2896
rect 1136 480 1164 2887
rect 1412 2854 1440 5510
rect 1504 3398 1532 6598
rect 1596 3738 1624 7262
rect 1780 4570 1808 7919
rect 1872 7313 1900 10254
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1858 7304 1914 7313
rect 1858 7239 1914 7248
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1872 5574 1900 6734
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1858 4720 1914 4729
rect 1858 4655 1860 4664
rect 1912 4655 1914 4664
rect 1860 4626 1912 4632
rect 1780 4542 1900 4570
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1766 3632 1822 3641
rect 1766 3567 1822 3576
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1490 3224 1546 3233
rect 1490 3159 1546 3168
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1412 1698 1440 2450
rect 1400 1692 1452 1698
rect 1400 1634 1452 1640
rect 1504 1578 1532 3159
rect 1412 1550 1532 1578
rect 1412 480 1440 1550
rect 1780 480 1808 3567
rect 1872 1766 1900 4542
rect 1964 3738 1992 8774
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1860 1760 1912 1766
rect 1860 1702 1912 1708
rect 2056 1465 2084 15438
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2228 13320 2280 13326
rect 2226 13288 2228 13297
rect 2280 13288 2282 13297
rect 2226 13223 2282 13232
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2240 12209 2268 12582
rect 2226 12200 2282 12209
rect 2226 12135 2282 12144
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2148 9654 2176 10610
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2332 8838 2360 15302
rect 2424 14521 2452 15982
rect 2410 14512 2466 14521
rect 2410 14447 2466 14456
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2424 8786 2452 11154
rect 2516 10742 2544 13806
rect 2608 12753 2636 16594
rect 2700 15609 2728 17070
rect 2792 16794 2820 19520
rect 3054 17368 3110 17377
rect 3054 17303 3110 17312
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2778 16416 2834 16425
rect 2778 16351 2834 16360
rect 2686 15600 2742 15609
rect 2686 15535 2742 15544
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 2700 14362 2728 15370
rect 2792 14550 2820 16351
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 2700 14334 2912 14362
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2594 12744 2650 12753
rect 2594 12679 2650 12688
rect 2596 11076 2648 11082
rect 2596 11018 2648 11024
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2608 10538 2636 11018
rect 2700 11014 2728 13330
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2792 12442 2820 13262
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2884 12186 2912 14334
rect 2976 13734 3004 17002
rect 3068 15706 3096 17303
rect 3160 17202 3188 19520
rect 3528 17610 3556 19520
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 3421 17436 3717 17456
rect 3477 17434 3501 17436
rect 3557 17434 3581 17436
rect 3637 17434 3661 17436
rect 3499 17382 3501 17434
rect 3563 17382 3575 17434
rect 3637 17382 3639 17434
rect 3477 17380 3501 17382
rect 3557 17380 3581 17382
rect 3637 17380 3661 17382
rect 3421 17360 3717 17380
rect 3804 17270 3832 19520
rect 4068 18012 4120 18018
rect 4068 17954 4120 17960
rect 3792 17264 3844 17270
rect 3792 17206 3844 17212
rect 3148 17196 3200 17202
rect 3148 17138 3200 17144
rect 4080 17134 4108 17954
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3252 16522 3280 17070
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3344 16833 3372 16934
rect 3330 16824 3386 16833
rect 3330 16759 3386 16768
rect 3332 16720 3384 16726
rect 3332 16662 3384 16668
rect 3240 16516 3292 16522
rect 3240 16458 3292 16464
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 3252 15570 3280 16458
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 2976 12481 3004 13466
rect 2962 12472 3018 12481
rect 2962 12407 3018 12416
rect 2792 12158 2912 12186
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2792 10554 2820 12158
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11694 2912 12038
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2596 10532 2648 10538
rect 2596 10474 2648 10480
rect 2700 10526 2820 10554
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2608 9586 2636 9862
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2502 9480 2558 9489
rect 2502 9415 2504 9424
rect 2556 9415 2558 9424
rect 2504 9386 2556 9392
rect 2700 9058 2728 10526
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 10266 2820 10406
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2792 9178 2820 10066
rect 2884 10033 2912 11086
rect 2870 10024 2926 10033
rect 2870 9959 2926 9968
rect 2976 9518 3004 11834
rect 3068 11393 3096 14962
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 3146 13832 3202 13841
rect 3146 13767 3202 13776
rect 3160 13190 3188 13767
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3160 12442 3188 12650
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3252 12322 3280 14826
rect 3344 14074 3372 16662
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3421 16348 3717 16368
rect 3477 16346 3501 16348
rect 3557 16346 3581 16348
rect 3637 16346 3661 16348
rect 3499 16294 3501 16346
rect 3563 16294 3575 16346
rect 3637 16294 3639 16346
rect 3477 16292 3501 16294
rect 3557 16292 3581 16294
rect 3637 16292 3661 16294
rect 3421 16272 3717 16292
rect 3608 15972 3660 15978
rect 3608 15914 3660 15920
rect 3620 15473 3648 15914
rect 3606 15464 3662 15473
rect 3606 15399 3662 15408
rect 3421 15260 3717 15280
rect 3477 15258 3501 15260
rect 3557 15258 3581 15260
rect 3637 15258 3661 15260
rect 3499 15206 3501 15258
rect 3563 15206 3575 15258
rect 3637 15206 3639 15258
rect 3477 15204 3501 15206
rect 3557 15204 3581 15206
rect 3637 15204 3661 15206
rect 3421 15184 3717 15204
rect 3424 15088 3476 15094
rect 3424 15030 3476 15036
rect 3436 14414 3464 15030
rect 3804 14958 3832 16390
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3421 14172 3717 14192
rect 3477 14170 3501 14172
rect 3557 14170 3581 14172
rect 3637 14170 3661 14172
rect 3499 14118 3501 14170
rect 3563 14118 3575 14170
rect 3637 14118 3639 14170
rect 3477 14116 3501 14118
rect 3557 14116 3581 14118
rect 3637 14116 3661 14118
rect 3421 14096 3717 14116
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3332 13456 3384 13462
rect 3332 13398 3384 13404
rect 3160 12294 3280 12322
rect 3160 11898 3188 12294
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3054 11384 3110 11393
rect 3054 11319 3110 11328
rect 3056 10736 3108 10742
rect 3056 10678 3108 10684
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2596 9036 2648 9042
rect 2700 9030 2820 9058
rect 2596 8978 2648 8984
rect 2424 8758 2544 8786
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2134 7848 2190 7857
rect 2134 7783 2190 7792
rect 2148 6882 2176 7783
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2240 7342 2268 7686
rect 2332 7410 2360 8230
rect 2424 7426 2452 8570
rect 2516 7585 2544 8758
rect 2502 7576 2558 7585
rect 2502 7511 2558 7520
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2415 7398 2452 7426
rect 2228 7336 2280 7342
rect 2415 7290 2443 7398
rect 2228 7278 2280 7284
rect 2332 7262 2443 7290
rect 2332 6934 2360 7262
rect 2320 6928 2372 6934
rect 2148 6854 2268 6882
rect 2320 6870 2372 6876
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2148 6390 2176 6734
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2148 5778 2176 6326
rect 2240 6254 2268 6854
rect 2228 6248 2280 6254
rect 2608 6225 2636 8978
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2700 8294 2728 8910
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2686 8120 2742 8129
rect 2686 8055 2742 8064
rect 2700 8022 2728 8055
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2792 7834 2820 9030
rect 2700 7806 2820 7834
rect 2228 6190 2280 6196
rect 2594 6216 2650 6225
rect 2240 5846 2268 6190
rect 2594 6151 2650 6160
rect 2228 5840 2280 5846
rect 2228 5782 2280 5788
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2134 4584 2190 4593
rect 2134 4519 2190 4528
rect 2148 4026 2176 4519
rect 2148 3998 2268 4026
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2148 3738 2176 3878
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 2240 1850 2268 3998
rect 2332 3194 2360 4966
rect 2424 4758 2452 5510
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2412 4480 2464 4486
rect 2412 4422 2464 4428
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2148 1822 2268 1850
rect 2042 1456 2098 1465
rect 2042 1391 2098 1400
rect 2148 480 2176 1822
rect 2424 480 2452 4422
rect 2516 4146 2544 5170
rect 2700 5080 2728 7806
rect 2778 7712 2834 7721
rect 2778 7647 2834 7656
rect 2608 5052 2728 5080
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2502 4040 2558 4049
rect 2502 3975 2558 3984
rect 2516 3058 2544 3975
rect 2608 3505 2636 5052
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2700 3670 2728 4694
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2594 3496 2650 3505
rect 2792 3466 2820 7647
rect 2884 6905 2912 9454
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 9217 3004 9318
rect 2962 9208 3018 9217
rect 2962 9143 3018 9152
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2976 7721 3004 8774
rect 2962 7712 3018 7721
rect 2962 7647 3018 7656
rect 3068 7562 3096 10678
rect 2976 7534 3096 7562
rect 2870 6896 2926 6905
rect 2870 6831 2926 6840
rect 2976 5409 3004 7534
rect 3054 7440 3110 7449
rect 3160 7426 3188 11494
rect 3252 10810 3280 12174
rect 3344 11898 3372 13398
rect 3804 13394 3832 14894
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3421 13084 3717 13104
rect 3477 13082 3501 13084
rect 3557 13082 3581 13084
rect 3637 13082 3661 13084
rect 3499 13030 3501 13082
rect 3563 13030 3575 13082
rect 3637 13030 3639 13082
rect 3477 13028 3501 13030
rect 3557 13028 3581 13030
rect 3637 13028 3661 13030
rect 3421 13008 3717 13028
rect 3804 12866 3832 13330
rect 3712 12838 3832 12866
rect 3712 12782 3740 12838
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3792 12708 3844 12714
rect 3792 12650 3844 12656
rect 3421 11996 3717 12016
rect 3477 11994 3501 11996
rect 3557 11994 3581 11996
rect 3637 11994 3661 11996
rect 3499 11942 3501 11994
rect 3563 11942 3575 11994
rect 3637 11942 3639 11994
rect 3477 11940 3501 11942
rect 3557 11940 3581 11942
rect 3637 11940 3661 11942
rect 3421 11920 3717 11940
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3804 11762 3832 12650
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3421 10908 3717 10928
rect 3477 10906 3501 10908
rect 3557 10906 3581 10908
rect 3637 10906 3661 10908
rect 3499 10854 3501 10906
rect 3563 10854 3575 10906
rect 3637 10854 3639 10906
rect 3477 10852 3501 10854
rect 3557 10852 3581 10854
rect 3637 10852 3661 10854
rect 3421 10832 3717 10852
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3896 10282 3924 16458
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3804 10254 3924 10282
rect 3988 10266 4016 16594
rect 4172 16425 4200 19520
rect 4540 16726 4568 19520
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4528 16720 4580 16726
rect 4528 16662 4580 16668
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4158 16416 4214 16425
rect 4158 16351 4214 16360
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 3976 10260 4028 10266
rect 3252 7970 3280 10202
rect 3421 9820 3717 9840
rect 3477 9818 3501 9820
rect 3557 9818 3581 9820
rect 3637 9818 3661 9820
rect 3499 9766 3501 9818
rect 3563 9766 3575 9818
rect 3637 9766 3639 9818
rect 3477 9764 3501 9766
rect 3557 9764 3581 9766
rect 3637 9764 3661 9766
rect 3421 9744 3717 9764
rect 3700 9648 3752 9654
rect 3804 9636 3832 10254
rect 3976 10202 4028 10208
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3752 9608 3832 9636
rect 3700 9590 3752 9596
rect 3332 9512 3384 9518
rect 3384 9460 3832 9466
rect 3332 9454 3832 9460
rect 3344 9438 3832 9454
rect 3896 9450 3924 9998
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 9178 3372 9318
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3344 8072 3372 8842
rect 3421 8732 3717 8752
rect 3477 8730 3501 8732
rect 3557 8730 3581 8732
rect 3637 8730 3661 8732
rect 3499 8678 3501 8730
rect 3563 8678 3575 8730
rect 3637 8678 3639 8730
rect 3477 8676 3501 8678
rect 3557 8676 3581 8678
rect 3637 8676 3661 8678
rect 3421 8656 3717 8676
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3620 8401 3648 8434
rect 3606 8392 3662 8401
rect 3606 8327 3662 8336
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3344 8044 3464 8072
rect 3252 7942 3372 7970
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3110 7398 3188 7426
rect 3054 7375 3110 7384
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3068 6254 3096 7278
rect 3252 6458 3280 7822
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 2962 5400 3018 5409
rect 2962 5335 3018 5344
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 3068 4826 3096 5238
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2884 4282 2912 4626
rect 2976 4457 3004 4626
rect 2962 4448 3018 4457
rect 2962 4383 3018 4392
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 3252 3738 3280 5306
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3344 3618 3372 7942
rect 3436 7857 3464 8044
rect 3514 7984 3570 7993
rect 3514 7919 3570 7928
rect 3422 7848 3478 7857
rect 3528 7818 3556 7919
rect 3712 7857 3740 8230
rect 3698 7848 3754 7857
rect 3422 7783 3478 7792
rect 3516 7812 3568 7818
rect 3698 7783 3754 7792
rect 3516 7754 3568 7760
rect 3421 7644 3717 7664
rect 3477 7642 3501 7644
rect 3557 7642 3581 7644
rect 3637 7642 3661 7644
rect 3499 7590 3501 7642
rect 3563 7590 3575 7642
rect 3637 7590 3639 7642
rect 3477 7588 3501 7590
rect 3557 7588 3581 7590
rect 3637 7588 3661 7590
rect 3421 7568 3717 7588
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 3422 5128 3478 5137
rect 3422 5063 3424 5072
rect 3476 5063 3478 5072
rect 3424 5034 3476 5040
rect 3804 4690 3832 9438
rect 3884 9444 3936 9450
rect 4080 9432 4108 16186
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4172 15026 4200 15302
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4160 14884 4212 14890
rect 4160 14826 4212 14832
rect 4172 12238 4200 14826
rect 4264 14385 4292 16594
rect 4436 16040 4488 16046
rect 4436 15982 4488 15988
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4250 14376 4306 14385
rect 4250 14311 4306 14320
rect 4252 14272 4304 14278
rect 4356 14260 4384 15438
rect 4448 14278 4476 15982
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4304 14232 4384 14260
rect 4436 14272 4488 14278
rect 4252 14214 4304 14220
rect 4436 14214 4488 14220
rect 4540 13938 4568 15642
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4264 13841 4292 13874
rect 4250 13832 4306 13841
rect 4250 13767 4306 13776
rect 4540 13025 4568 13874
rect 4632 13138 4660 16730
rect 4710 16280 4766 16289
rect 4816 16250 4844 19520
rect 5184 17882 5212 19520
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 4986 17232 5042 17241
rect 4986 17167 4988 17176
rect 5040 17167 5042 17176
rect 4988 17138 5040 17144
rect 5460 16794 5488 17614
rect 5552 17134 5580 19520
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5736 16998 5764 17478
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5354 16688 5410 16697
rect 5354 16623 5356 16632
rect 5408 16623 5410 16632
rect 5356 16594 5408 16600
rect 5080 16516 5132 16522
rect 5080 16458 5132 16464
rect 4710 16215 4712 16224
rect 4764 16215 4766 16224
rect 4804 16244 4856 16250
rect 4712 16186 4764 16192
rect 4804 16186 4856 16192
rect 4894 16144 4950 16153
rect 4894 16079 4950 16088
rect 4712 15972 4764 15978
rect 4712 15914 4764 15920
rect 4724 14346 4752 15914
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4816 15162 4844 15846
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4908 14482 4936 16079
rect 4988 15428 5040 15434
rect 4988 15370 5040 15376
rect 5000 14958 5028 15370
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4712 14340 4764 14346
rect 4712 14282 4764 14288
rect 4816 14074 4844 14418
rect 4894 14376 4950 14385
rect 4894 14311 4950 14320
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4908 13954 4936 14311
rect 4816 13926 4936 13954
rect 4816 13530 4844 13926
rect 5000 13870 5028 14894
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4632 13110 5028 13138
rect 4526 13016 4582 13025
rect 4526 12951 4582 12960
rect 4710 12336 4766 12345
rect 4540 12280 4710 12288
rect 4540 12260 4712 12280
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4172 11744 4200 12174
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 11937 4384 12038
rect 4342 11928 4398 11937
rect 4342 11863 4398 11872
rect 4436 11824 4488 11830
rect 4436 11766 4488 11772
rect 4344 11756 4396 11762
rect 4172 11716 4344 11744
rect 4344 11698 4396 11704
rect 4342 11656 4398 11665
rect 4252 11620 4304 11626
rect 4342 11591 4398 11600
rect 4252 11562 4304 11568
rect 4264 10266 4292 11562
rect 4356 10266 4384 11591
rect 4448 11286 4476 11766
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4448 10198 4476 11018
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 3884 9386 3936 9392
rect 3988 9404 4108 9432
rect 3882 8528 3938 8537
rect 3882 8463 3938 8472
rect 3896 8430 3924 8463
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 7954 3924 8230
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3896 7206 3924 7754
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3988 6866 4016 9404
rect 4540 8974 4568 12260
rect 4764 12271 4766 12280
rect 4712 12242 4764 12248
rect 4896 12232 4948 12238
rect 4618 12200 4674 12209
rect 4618 12135 4674 12144
rect 4816 12192 4896 12220
rect 4632 11218 4660 12135
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4632 10198 4660 10474
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4436 8968 4488 8974
rect 4528 8968 4580 8974
rect 4436 8910 4488 8916
rect 4526 8936 4528 8945
rect 4580 8936 4582 8945
rect 4448 8838 4476 8910
rect 4526 8871 4582 8880
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4080 8430 4108 8570
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4158 8392 4214 8401
rect 4158 8327 4214 8336
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4080 7342 4108 7822
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3896 5642 3924 6054
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 3882 5536 3938 5545
rect 3882 5471 3938 5480
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3896 3618 3924 5471
rect 2976 3590 3372 3618
rect 3804 3590 3924 3618
rect 2594 3431 2650 3440
rect 2780 3460 2832 3466
rect 2780 3402 2832 3408
rect 2778 3088 2834 3097
rect 2504 3052 2556 3058
rect 2778 3023 2834 3032
rect 2504 2994 2556 3000
rect 2792 480 2820 3023
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2884 513 2912 2450
rect 2976 1834 3004 3590
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3148 3460 3200 3466
rect 3148 3402 3200 3408
rect 3160 3058 3188 3402
rect 3252 3126 3280 3470
rect 3421 3292 3717 3312
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 3068 2553 3096 2790
rect 3054 2544 3110 2553
rect 3054 2479 3110 2488
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3421 2128 3717 2148
rect 2964 1828 3016 1834
rect 2964 1770 3016 1776
rect 3148 1284 3200 1290
rect 3148 1226 3200 1232
rect 2870 504 2926 513
rect 110 0 166 480
rect 386 0 442 480
rect 754 0 810 480
rect 1122 0 1178 480
rect 1398 0 1454 480
rect 1766 0 1822 480
rect 2134 0 2190 480
rect 2410 0 2466 480
rect 2778 0 2834 480
rect 3160 480 3188 1226
rect 3516 1012 3568 1018
rect 3516 954 3568 960
rect 3528 480 3556 954
rect 3804 480 3832 3590
rect 3988 2514 4016 6802
rect 4172 6458 4200 8327
rect 4264 8090 4292 8774
rect 4342 8664 4398 8673
rect 4342 8599 4398 8608
rect 4356 8362 4384 8599
rect 4632 8566 4660 8978
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4434 8120 4490 8129
rect 4252 8084 4304 8090
rect 4434 8055 4436 8064
rect 4252 8026 4304 8032
rect 4488 8055 4490 8064
rect 4436 8026 4488 8032
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4250 7848 4306 7857
rect 4250 7783 4306 7792
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4172 6118 4200 6394
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 2990 4108 5510
rect 4264 5137 4292 7783
rect 4356 7546 4384 7890
rect 4632 7721 4660 8366
rect 4618 7712 4674 7721
rect 4618 7647 4674 7656
rect 4618 7576 4674 7585
rect 4344 7540 4396 7546
rect 4618 7511 4674 7520
rect 4344 7482 4396 7488
rect 4356 6934 4384 7482
rect 4344 6928 4396 6934
rect 4344 6870 4396 6876
rect 4434 6896 4490 6905
rect 4434 6831 4490 6840
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4250 5128 4306 5137
rect 4250 5063 4306 5072
rect 4264 4214 4292 5063
rect 4356 4758 4384 5306
rect 4344 4752 4396 4758
rect 4344 4694 4396 4700
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4321 4384 4422
rect 4342 4312 4398 4321
rect 4342 4247 4398 4256
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4172 3942 4200 4082
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4264 3738 4292 3946
rect 4448 3890 4476 6831
rect 4526 5808 4582 5817
rect 4632 5778 4660 7511
rect 4724 7478 4752 12038
rect 4816 11150 4844 12192
rect 4896 12174 4948 12180
rect 4896 11688 4948 11694
rect 4894 11656 4896 11665
rect 4948 11656 4950 11665
rect 4894 11591 4950 11600
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4816 10674 4844 11086
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4816 10198 4844 10610
rect 4908 10606 4936 11591
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4908 10266 4936 10542
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4802 10024 4858 10033
rect 4802 9959 4858 9968
rect 4816 9042 4844 9959
rect 4908 9722 4936 10202
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 4896 9580 4948 9586
rect 5000 9568 5028 13110
rect 5092 12288 5120 16458
rect 5644 16114 5672 16934
rect 5828 16561 5856 19520
rect 6196 17338 6224 19520
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 6368 17264 6420 17270
rect 6368 17206 6420 17212
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 5886 16892 6182 16912
rect 5942 16890 5966 16892
rect 6022 16890 6046 16892
rect 6102 16890 6126 16892
rect 5964 16838 5966 16890
rect 6028 16838 6040 16890
rect 6102 16838 6104 16890
rect 5942 16836 5966 16838
rect 6022 16836 6046 16838
rect 6102 16836 6126 16838
rect 5886 16816 6182 16836
rect 6288 16794 6316 17002
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 5814 16552 5870 16561
rect 5814 16487 5870 16496
rect 6380 16454 6408 17206
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 14074 5212 15846
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5276 13802 5304 15098
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 5170 13016 5226 13025
rect 5170 12951 5226 12960
rect 5184 12714 5212 12951
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5092 12260 5212 12288
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 5092 10538 5120 12106
rect 5184 12102 5212 12260
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 5184 10810 5212 11562
rect 5276 11150 5304 12582
rect 5368 11354 5396 15302
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5460 13462 5488 14758
rect 5552 14550 5580 16050
rect 5724 15496 5776 15502
rect 5722 15464 5724 15473
rect 5776 15464 5778 15473
rect 5632 15428 5684 15434
rect 5722 15399 5778 15408
rect 5632 15370 5684 15376
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5644 14414 5672 15370
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5552 13462 5580 14350
rect 5630 13832 5686 13841
rect 5630 13767 5686 13776
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5644 13258 5672 13767
rect 5828 13394 5856 16118
rect 6196 16068 6408 16096
rect 6196 15978 6224 16068
rect 6184 15972 6236 15978
rect 6184 15914 6236 15920
rect 5886 15804 6182 15824
rect 5942 15802 5966 15804
rect 6022 15802 6046 15804
rect 6102 15802 6126 15804
rect 5964 15750 5966 15802
rect 6028 15750 6040 15802
rect 6102 15750 6104 15802
rect 5942 15748 5966 15750
rect 6022 15748 6046 15750
rect 6102 15748 6126 15750
rect 5886 15728 6182 15748
rect 6380 14929 6408 16068
rect 6564 16017 6592 19520
rect 6932 17746 6960 19520
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 7208 16590 7236 19520
rect 7576 18494 7604 19520
rect 7564 18488 7616 18494
rect 7564 18430 7616 18436
rect 7944 17950 7972 19520
rect 7932 17944 7984 17950
rect 7932 17886 7984 17892
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7656 17264 7708 17270
rect 7656 17206 7708 17212
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 6656 16182 6684 16526
rect 7010 16280 7066 16289
rect 7010 16215 7066 16224
rect 6644 16176 6696 16182
rect 6828 16176 6880 16182
rect 6644 16118 6696 16124
rect 6826 16144 6828 16153
rect 6920 16176 6972 16182
rect 6880 16144 6882 16153
rect 6550 16008 6606 16017
rect 6550 15943 6606 15952
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6366 14920 6422 14929
rect 6366 14855 6422 14864
rect 5886 14716 6182 14736
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6126 14716
rect 5964 14662 5966 14714
rect 6028 14662 6040 14714
rect 6102 14662 6104 14714
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6126 14662
rect 5886 14640 6182 14660
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 6288 14074 6316 14486
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 5886 13628 6182 13648
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6126 13628
rect 5964 13574 5966 13626
rect 6028 13574 6040 13626
rect 6102 13574 6104 13626
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6126 13574
rect 5886 13552 6182 13572
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5632 13252 5684 13258
rect 5632 13194 5684 13200
rect 5644 12374 5672 13194
rect 6288 12986 6316 13398
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 5886 12540 6182 12560
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6126 12540
rect 5964 12486 5966 12538
rect 6028 12486 6040 12538
rect 6102 12486 6104 12538
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6126 12486
rect 5886 12464 6182 12484
rect 6380 12442 6408 13738
rect 6564 12918 6592 14962
rect 6656 14793 6684 16118
rect 6920 16118 6972 16124
rect 6826 16079 6882 16088
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6642 14784 6698 14793
rect 6642 14719 6698 14728
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6656 13410 6684 14554
rect 6748 14396 6776 14894
rect 6840 14550 6868 15574
rect 6932 15473 6960 16118
rect 6918 15464 6974 15473
rect 6918 15399 6974 15408
rect 6932 15366 6960 15399
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6828 14408 6880 14414
rect 6748 14368 6828 14396
rect 6828 14350 6880 14356
rect 6840 13938 6868 14350
rect 6828 13932 6880 13938
rect 7024 13920 7052 16215
rect 7194 16144 7250 16153
rect 7380 16108 7432 16114
rect 7194 16079 7250 16088
rect 7208 16046 7236 16079
rect 7300 16068 7380 16096
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7300 15706 7328 16068
rect 7380 16050 7432 16056
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7208 15144 7236 15302
rect 7208 15116 7328 15144
rect 7194 15056 7250 15065
rect 7194 14991 7250 15000
rect 7024 13892 7144 13920
rect 6828 13874 6880 13880
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6748 13530 6776 13806
rect 6840 13802 6868 13874
rect 6828 13796 6880 13802
rect 6828 13738 6880 13744
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6656 13382 6776 13410
rect 6840 13394 6868 13738
rect 7116 13569 7144 13892
rect 7102 13560 7158 13569
rect 7102 13495 7158 13504
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6564 12753 6592 12854
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6550 12744 6606 12753
rect 6550 12679 6606 12688
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5632 12368 5684 12374
rect 5632 12310 5684 12316
rect 5552 11937 5580 12310
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 5538 11928 5594 11937
rect 6380 11914 6408 12242
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 5538 11863 5594 11872
rect 5632 11892 5684 11898
rect 6380 11886 6500 11914
rect 6564 11898 6592 12174
rect 6656 12102 6684 12786
rect 6748 12238 6776 13382
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6932 13297 6960 13398
rect 6918 13288 6974 13297
rect 6918 13223 6974 13232
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6932 12170 6960 12718
rect 7116 12481 7144 13126
rect 7102 12472 7158 12481
rect 7102 12407 7158 12416
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 5632 11834 5684 11840
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5460 11150 5488 11290
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5092 10062 5120 10474
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5080 9920 5132 9926
rect 5078 9888 5080 9897
rect 5132 9888 5134 9897
rect 5078 9823 5134 9832
rect 5184 9722 5212 10746
rect 5552 10606 5580 11630
rect 5644 10810 5672 11834
rect 6366 11792 6422 11801
rect 6366 11727 6422 11736
rect 5814 11656 5870 11665
rect 5814 11591 5870 11600
rect 5828 11218 5856 11591
rect 6274 11520 6330 11529
rect 5886 11452 6182 11472
rect 6274 11455 6330 11464
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6126 11452
rect 5964 11398 5966 11450
rect 6028 11398 6040 11450
rect 6102 11398 6104 11450
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6126 11398
rect 5886 11376 6182 11396
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5908 11212 5960 11218
rect 6288 11200 6316 11455
rect 5960 11172 6316 11200
rect 5908 11154 5960 11160
rect 5814 11112 5870 11121
rect 5814 11047 5816 11056
rect 5868 11047 5870 11056
rect 5816 11018 5868 11024
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5460 10418 5488 10474
rect 5368 10390 5488 10418
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5276 9722 5304 9930
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 4948 9540 5028 9568
rect 4896 9522 4948 9528
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 4804 8424 4856 8430
rect 4908 8412 4936 9522
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 4988 8968 5040 8974
rect 4986 8936 4988 8945
rect 5040 8936 5042 8945
rect 4986 8871 5042 8880
rect 4856 8384 4936 8412
rect 4804 8366 4856 8372
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4724 6798 4752 7414
rect 4816 7324 4844 8366
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4908 7954 4936 8230
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4896 7336 4948 7342
rect 4816 7296 4896 7324
rect 4896 7278 4948 7284
rect 4908 6798 4936 7278
rect 5092 6866 5120 8978
rect 5184 8974 5212 9318
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5368 7936 5396 10390
rect 5886 10364 6182 10384
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6126 10364
rect 5964 10310 5966 10362
rect 6028 10310 6040 10362
rect 6102 10310 6104 10362
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6126 10310
rect 5886 10288 6182 10308
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5460 10062 5488 10202
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5538 9888 5594 9897
rect 5538 9823 5594 9832
rect 5552 9450 5580 9823
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5630 9208 5686 9217
rect 5630 9143 5686 9152
rect 5644 9110 5672 9143
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5722 9072 5778 9081
rect 5722 9007 5778 9016
rect 5276 7908 5396 7936
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4526 5743 4582 5752
rect 4620 5772 4672 5778
rect 4356 3862 4476 3890
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4172 3058 4200 3334
rect 4252 3188 4304 3194
rect 4356 3176 4384 3862
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4448 3233 4476 3674
rect 4304 3148 4384 3176
rect 4434 3224 4490 3233
rect 4434 3159 4490 3168
rect 4252 3130 4304 3136
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4448 2582 4476 2994
rect 4436 2576 4488 2582
rect 4436 2518 4488 2524
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4158 2000 4214 2009
rect 4356 1970 4384 2382
rect 4158 1935 4214 1944
rect 4344 1964 4396 1970
rect 4172 480 4200 1935
rect 4344 1906 4396 1912
rect 4540 480 4568 5743
rect 4620 5714 4672 5720
rect 4632 5302 4660 5714
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4632 4457 4660 4490
rect 4618 4448 4674 4457
rect 4618 4383 4674 4392
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4632 3058 4660 4150
rect 4724 3380 4752 6598
rect 4908 6322 4936 6734
rect 5276 6662 5304 7908
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 6662 5488 7686
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5262 6352 5318 6361
rect 4896 6316 4948 6322
rect 5262 6287 5318 6296
rect 4896 6258 4948 6264
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 5092 5545 5120 5578
rect 5078 5536 5134 5545
rect 5078 5471 5134 5480
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4908 4570 4936 5102
rect 5080 4616 5132 4622
rect 4908 4564 5080 4570
rect 4908 4558 5132 4564
rect 4908 4542 5120 4558
rect 4908 4282 4936 4542
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4986 4312 5042 4321
rect 4896 4276 4948 4282
rect 5092 4282 5120 4422
rect 4986 4247 5042 4256
rect 5080 4276 5132 4282
rect 4896 4218 4948 4224
rect 4908 4078 4936 4218
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4908 3618 4936 4014
rect 5000 3738 5028 4247
rect 5080 4218 5132 4224
rect 5078 4176 5134 4185
rect 5078 4111 5134 4120
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4908 3590 5028 3618
rect 4724 3352 4844 3380
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4618 2816 4674 2825
rect 4618 2751 4674 2760
rect 4632 2514 4660 2751
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4816 480 4844 3352
rect 4896 3120 4948 3126
rect 5000 3074 5028 3590
rect 4948 3068 5028 3074
rect 4896 3062 5028 3068
rect 4908 3046 5028 3062
rect 5000 2825 5028 3046
rect 4986 2816 5042 2825
rect 4986 2751 5042 2760
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5000 1630 5028 2382
rect 4988 1624 5040 1630
rect 4988 1566 5040 1572
rect 5092 1290 5120 4111
rect 5184 4010 5212 5646
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5184 3534 5212 3946
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5276 3210 5304 6287
rect 5460 6186 5488 6598
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5552 5846 5580 6122
rect 5736 5930 5764 9007
rect 5828 8673 5856 9454
rect 6276 9444 6328 9450
rect 6276 9386 6328 9392
rect 5886 9276 6182 9296
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6126 9276
rect 5964 9222 5966 9274
rect 6028 9222 6040 9274
rect 6102 9222 6104 9274
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6126 9222
rect 5886 9200 6182 9220
rect 5814 8664 5870 8673
rect 5814 8599 5870 8608
rect 6288 8566 6316 9386
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 5886 8188 6182 8208
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6126 8188
rect 5964 8134 5966 8186
rect 6028 8134 6040 8186
rect 6102 8134 6104 8186
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6126 8134
rect 5886 8112 6182 8132
rect 5908 7880 5960 7886
rect 5960 7840 6040 7868
rect 5908 7822 5960 7828
rect 6012 7342 6040 7840
rect 6288 7546 6316 8366
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6288 7410 6316 7482
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 5886 7100 6182 7120
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6126 7100
rect 5964 7046 5966 7098
rect 6028 7046 6040 7098
rect 6102 7046 6104 7098
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6126 7046
rect 5886 7024 6182 7044
rect 6288 6769 6316 7142
rect 6274 6760 6330 6769
rect 6274 6695 6330 6704
rect 6288 6390 6316 6695
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 5736 5902 5856 5930
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5460 5166 5488 5510
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5644 5098 5672 5782
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5368 4321 5396 4626
rect 5354 4312 5410 4321
rect 5354 4247 5410 4256
rect 5552 3942 5580 4626
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5460 3738 5488 3878
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5184 3182 5304 3210
rect 5080 1284 5132 1290
rect 5080 1226 5132 1232
rect 5184 480 5212 3182
rect 5460 2582 5488 3470
rect 5552 3194 5580 3878
rect 5644 3466 5672 5034
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5630 3224 5686 3233
rect 5540 3188 5592 3194
rect 5630 3159 5686 3168
rect 5540 3130 5592 3136
rect 5644 2990 5672 3159
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5552 2582 5580 2790
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 5644 1442 5672 2790
rect 5736 2650 5764 2858
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5552 1414 5672 1442
rect 5552 480 5580 1414
rect 5828 480 5856 5902
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 5886 3836 6182 3856
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 6288 3602 6316 4966
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 6288 2632 6316 2994
rect 6380 2922 6408 11727
rect 6472 10810 6500 11886
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6840 11762 6868 12038
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 11218 6960 11494
rect 7010 11384 7066 11393
rect 7010 11319 7066 11328
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7024 11014 7052 11319
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6642 10704 6698 10713
rect 6642 10639 6698 10648
rect 6550 10024 6606 10033
rect 6550 9959 6606 9968
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 6368 2916 6420 2922
rect 6368 2858 6420 2864
rect 6472 2650 6500 6122
rect 6564 3058 6592 9959
rect 6656 5302 6684 10639
rect 7024 10606 7052 10950
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6840 9586 6868 10066
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 8838 6960 9318
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6920 8424 6972 8430
rect 7024 8412 7052 10542
rect 7116 10470 7144 12407
rect 7208 12306 7236 14991
rect 7300 13394 7328 15116
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7286 13288 7342 13297
rect 7286 13223 7342 13232
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7300 11626 7328 13223
rect 7392 12374 7420 15846
rect 7484 14618 7512 17138
rect 7668 16726 7696 17206
rect 7748 16992 7800 16998
rect 7746 16960 7748 16969
rect 7800 16960 7802 16969
rect 7746 16895 7802 16904
rect 7746 16824 7802 16833
rect 7852 16794 7880 17750
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 7746 16759 7802 16768
rect 7840 16788 7892 16794
rect 7656 16720 7708 16726
rect 7656 16662 7708 16668
rect 7760 16590 7788 16759
rect 7840 16730 7892 16736
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7562 16280 7618 16289
rect 7562 16215 7618 16224
rect 7576 16114 7604 16215
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7576 14958 7604 15914
rect 7668 15473 7696 16526
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7746 16144 7802 16153
rect 7746 16079 7802 16088
rect 7760 16046 7788 16079
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7654 15464 7710 15473
rect 7654 15399 7710 15408
rect 7852 15366 7880 16390
rect 7944 16114 7972 17002
rect 8036 16454 8064 17138
rect 8114 16824 8170 16833
rect 8114 16759 8116 16768
rect 8168 16759 8170 16768
rect 8116 16730 8168 16736
rect 8220 16674 8248 19520
rect 8588 17626 8616 19520
rect 8956 17950 8984 19520
rect 8852 17944 8904 17950
rect 8850 17912 8852 17921
rect 8944 17944 8996 17950
rect 8904 17912 8906 17921
rect 8944 17886 8996 17892
rect 8850 17847 8906 17856
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 8758 17640 8814 17649
rect 8588 17598 8708 17626
rect 8352 17436 8648 17456
rect 8408 17434 8432 17436
rect 8488 17434 8512 17436
rect 8568 17434 8592 17436
rect 8430 17382 8432 17434
rect 8494 17382 8506 17434
rect 8568 17382 8570 17434
rect 8408 17380 8432 17382
rect 8488 17380 8512 17382
rect 8568 17380 8592 17382
rect 8352 17360 8648 17380
rect 8482 17096 8538 17105
rect 8482 17031 8484 17040
rect 8536 17031 8538 17040
rect 8484 17002 8536 17008
rect 8298 16824 8354 16833
rect 8298 16759 8300 16768
rect 8352 16759 8354 16768
rect 8300 16730 8352 16736
rect 8128 16646 8248 16674
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 8036 15688 8064 16390
rect 8128 16028 8156 16646
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8220 16425 8248 16458
rect 8680 16454 8708 17598
rect 8758 17575 8814 17584
rect 8772 17066 8800 17575
rect 8944 17264 8996 17270
rect 8944 17206 8996 17212
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 8864 16794 8892 17070
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8668 16448 8720 16454
rect 8206 16416 8262 16425
rect 8668 16390 8720 16396
rect 8206 16351 8262 16360
rect 8352 16348 8648 16368
rect 8408 16346 8432 16348
rect 8488 16346 8512 16348
rect 8568 16346 8592 16348
rect 8430 16294 8432 16346
rect 8494 16294 8506 16346
rect 8568 16294 8570 16346
rect 8408 16292 8432 16294
rect 8488 16292 8512 16294
rect 8568 16292 8592 16294
rect 8352 16272 8648 16292
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8300 16040 8352 16046
rect 8128 16000 8248 16028
rect 7944 15660 8064 15688
rect 8114 15736 8170 15745
rect 8114 15671 8116 15680
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7562 14784 7618 14793
rect 7562 14719 7618 14728
rect 7576 14618 7604 14719
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7484 13870 7512 14554
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7576 14074 7604 14418
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7668 13734 7696 15302
rect 7944 15065 7972 15660
rect 8168 15671 8170 15680
rect 8116 15642 8168 15648
rect 8220 15638 8248 16000
rect 8300 15982 8352 15988
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8036 15094 8064 15506
rect 8312 15502 8340 15982
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8024 15088 8076 15094
rect 7930 15056 7986 15065
rect 8024 15030 8076 15036
rect 8128 15026 8156 15438
rect 8404 15434 8432 15846
rect 8496 15570 8524 16050
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8392 15428 8444 15434
rect 8392 15370 8444 15376
rect 8352 15260 8648 15280
rect 8408 15258 8432 15260
rect 8488 15258 8512 15260
rect 8568 15258 8592 15260
rect 8430 15206 8432 15258
rect 8494 15206 8506 15258
rect 8568 15206 8570 15258
rect 8408 15204 8432 15206
rect 8488 15204 8512 15206
rect 8568 15204 8592 15206
rect 8352 15184 8648 15204
rect 8680 15162 8708 15438
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 7930 14991 7986 15000
rect 8116 15020 8168 15026
rect 7748 14476 7800 14482
rect 7944 14464 7972 14991
rect 8116 14962 8168 14968
rect 8390 14920 8446 14929
rect 8300 14884 8352 14890
rect 8390 14855 8392 14864
rect 8300 14826 8352 14832
rect 8444 14855 8446 14864
rect 8392 14826 8444 14832
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 7800 14436 7972 14464
rect 7748 14418 7800 14424
rect 7944 14006 7972 14436
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 8128 13938 8156 14758
rect 8312 14482 8340 14826
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8680 14521 8708 14758
rect 8666 14512 8722 14521
rect 8300 14476 8352 14482
rect 8666 14447 8722 14456
rect 8300 14418 8352 14424
rect 8668 14340 8720 14346
rect 8668 14282 8720 14288
rect 8352 14172 8648 14192
rect 8408 14170 8432 14172
rect 8488 14170 8512 14172
rect 8568 14170 8592 14172
rect 8430 14118 8432 14170
rect 8494 14118 8506 14170
rect 8568 14118 8570 14170
rect 8408 14116 8432 14118
rect 8488 14116 8512 14118
rect 8568 14116 8592 14118
rect 8352 14096 8648 14116
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8680 13870 8708 14282
rect 8772 14278 8800 15846
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7392 11150 7420 11698
rect 7484 11506 7512 13194
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7576 11626 7604 13126
rect 7668 12714 7696 13330
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8036 12986 8064 13262
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 8128 12782 8156 13738
rect 8392 13728 8444 13734
rect 8206 13696 8262 13705
rect 8392 13670 8444 13676
rect 8206 13631 8262 13640
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 7656 12708 7708 12714
rect 7932 12708 7984 12714
rect 7656 12650 7708 12656
rect 7852 12668 7932 12696
rect 7668 12374 7696 12650
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7564 11620 7616 11626
rect 7564 11562 7616 11568
rect 7484 11478 7604 11506
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7208 10266 7236 10950
rect 7300 10810 7328 10950
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7392 10606 7420 11086
rect 7484 10674 7512 11154
rect 7576 10810 7604 11478
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7392 10130 7420 10542
rect 7470 10432 7526 10441
rect 7470 10367 7526 10376
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7102 9344 7158 9353
rect 7102 9279 7158 9288
rect 6972 8384 7052 8412
rect 6920 8366 6972 8372
rect 6840 7342 6868 8366
rect 7012 8288 7064 8294
rect 7116 8276 7144 9279
rect 7484 9024 7512 10367
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 9382 7604 10066
rect 7656 9920 7708 9926
rect 7654 9888 7656 9897
rect 7708 9888 7710 9897
rect 7654 9823 7710 9832
rect 7654 9616 7710 9625
rect 7654 9551 7710 9560
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7562 9208 7618 9217
rect 7562 9143 7618 9152
rect 7576 9110 7604 9143
rect 7668 9110 7696 9551
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7392 8996 7512 9024
rect 7194 8936 7250 8945
rect 7194 8871 7250 8880
rect 7208 8378 7236 8871
rect 7392 8838 7420 8996
rect 7470 8936 7526 8945
rect 7760 8906 7788 12582
rect 7852 11354 7880 12668
rect 7932 12650 7984 12656
rect 7930 12336 7986 12345
rect 7930 12271 7932 12280
rect 7984 12271 7986 12280
rect 7932 12242 7984 12248
rect 7930 12200 7986 12209
rect 7930 12135 7986 12144
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7852 9450 7880 11290
rect 7944 10418 7972 12135
rect 8220 12084 8248 13631
rect 8404 13530 8432 13670
rect 8680 13530 8708 13806
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8352 13084 8648 13104
rect 8408 13082 8432 13084
rect 8488 13082 8512 13084
rect 8568 13082 8592 13084
rect 8430 13030 8432 13082
rect 8494 13030 8506 13082
rect 8568 13030 8570 13082
rect 8408 13028 8432 13030
rect 8488 13028 8512 13030
rect 8568 13028 8592 13030
rect 8352 13008 8648 13028
rect 8680 12850 8708 13466
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8588 12306 8616 12718
rect 8864 12628 8892 16594
rect 8956 14346 8984 17206
rect 9036 16720 9088 16726
rect 9036 16662 9088 16668
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 8942 14240 8998 14249
rect 8942 14175 8998 14184
rect 8772 12600 8892 12628
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8668 12164 8720 12170
rect 8588 12124 8668 12152
rect 8588 12084 8616 12124
rect 8668 12106 8720 12112
rect 8220 12073 8616 12084
rect 8206 12064 8616 12073
rect 8262 12056 8616 12064
rect 8206 11999 8262 12008
rect 8352 11996 8648 12016
rect 8408 11994 8432 11996
rect 8488 11994 8512 11996
rect 8568 11994 8592 11996
rect 8430 11942 8432 11994
rect 8494 11942 8506 11994
rect 8568 11942 8570 11994
rect 8408 11940 8432 11942
rect 8488 11940 8512 11942
rect 8568 11940 8592 11942
rect 8206 11928 8262 11937
rect 8352 11920 8648 11940
rect 8206 11863 8262 11872
rect 8220 11354 8248 11863
rect 8576 11824 8628 11830
rect 8576 11766 8628 11772
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8496 11665 8524 11698
rect 8482 11656 8538 11665
rect 8482 11591 8538 11600
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8588 10996 8616 11766
rect 8666 11656 8722 11665
rect 8666 11591 8722 11600
rect 8680 11121 8708 11591
rect 8666 11112 8722 11121
rect 8666 11047 8722 11056
rect 8588 10968 8708 10996
rect 8352 10908 8648 10928
rect 8408 10906 8432 10908
rect 8488 10906 8512 10908
rect 8568 10906 8592 10908
rect 8430 10854 8432 10906
rect 8494 10854 8506 10906
rect 8568 10854 8570 10906
rect 8408 10852 8432 10854
rect 8488 10852 8512 10854
rect 8568 10852 8592 10854
rect 8352 10832 8648 10852
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8220 10441 8248 10542
rect 7935 10390 7972 10418
rect 8206 10432 8262 10441
rect 7935 10180 7963 10390
rect 8206 10367 8262 10376
rect 8206 10296 8262 10305
rect 8024 10260 8076 10266
rect 8206 10231 8262 10240
rect 8024 10202 8076 10208
rect 7935 10152 7972 10180
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7852 8906 7880 9046
rect 7470 8871 7472 8880
rect 7524 8871 7526 8880
rect 7748 8900 7800 8906
rect 7472 8842 7524 8848
rect 7748 8842 7800 8848
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7208 8362 7420 8378
rect 7196 8356 7420 8362
rect 7248 8350 7420 8356
rect 7196 8298 7248 8304
rect 7392 8294 7420 8350
rect 7064 8248 7144 8276
rect 7012 8230 7064 8236
rect 7116 7818 7144 8248
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7470 8120 7526 8129
rect 7470 8055 7526 8064
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 7484 7546 7512 8055
rect 7852 7954 7880 8502
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7838 7712 7894 7721
rect 7576 7546 7604 7686
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 6828 7336 6880 7342
rect 7668 7324 7696 7686
rect 7838 7647 7894 7656
rect 6828 7278 6880 7284
rect 7576 7296 7696 7324
rect 6840 6254 6868 7278
rect 7010 7032 7066 7041
rect 7010 6967 7012 6976
rect 7064 6967 7066 6976
rect 7012 6938 7064 6944
rect 7576 6798 7604 7296
rect 7852 7177 7880 7647
rect 7838 7168 7894 7177
rect 7838 7103 7894 7112
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7576 6254 7604 6734
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6748 5166 6776 5714
rect 6840 5710 6868 6190
rect 7668 6118 7696 6802
rect 7852 6769 7880 6802
rect 7838 6760 7894 6769
rect 7838 6695 7894 6704
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7576 5930 7604 6054
rect 7852 5930 7880 6258
rect 7576 5902 7880 5930
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6642 4856 6698 4865
rect 6642 4791 6698 4800
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6656 2938 6684 4791
rect 6748 4622 6776 5102
rect 6840 4865 6868 5238
rect 6920 5160 6972 5166
rect 7104 5160 7156 5166
rect 6972 5120 7052 5148
rect 6920 5102 6972 5108
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6826 4856 6882 4865
rect 6826 4791 6882 4800
rect 6828 4752 6880 4758
rect 6932 4729 6960 4966
rect 7024 4758 7052 5120
rect 7104 5102 7156 5108
rect 7012 4752 7064 4758
rect 6828 4694 6880 4700
rect 6918 4720 6974 4729
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6748 4078 6776 4558
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6748 3058 6776 3538
rect 6840 3466 6868 4694
rect 7012 4694 7064 4700
rect 6918 4655 6974 4664
rect 7116 4282 7144 5102
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7024 4010 7052 4218
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 6932 3602 6960 3946
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 7116 3398 7144 4218
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7208 3194 7236 5714
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6564 2910 6684 2938
rect 7012 2916 7064 2922
rect 6196 2604 6316 2632
rect 6460 2644 6512 2650
rect 6196 480 6224 2604
rect 6460 2586 6512 2592
rect 6564 480 6592 2910
rect 7012 2858 7064 2864
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7024 2825 7052 2858
rect 7010 2816 7066 2825
rect 7010 2751 7066 2760
rect 7024 2310 7052 2751
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 6920 1896 6972 1902
rect 6920 1838 6972 1844
rect 6932 480 6960 1838
rect 7208 480 7236 2858
rect 7300 1018 7328 5782
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7838 5536 7894 5545
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7392 4486 7420 4626
rect 7380 4480 7432 4486
rect 7472 4480 7524 4486
rect 7380 4422 7432 4428
rect 7470 4448 7472 4457
rect 7524 4448 7526 4457
rect 7392 2378 7420 4422
rect 7470 4383 7526 4392
rect 7576 4185 7604 5510
rect 7838 5471 7894 5480
rect 7746 5400 7802 5409
rect 7746 5335 7802 5344
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7668 4758 7696 5102
rect 7760 4758 7788 5335
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7746 4312 7802 4321
rect 7852 4282 7880 5471
rect 7746 4247 7802 4256
rect 7840 4276 7892 4282
rect 7562 4176 7618 4185
rect 7562 4111 7618 4120
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7484 2446 7512 3946
rect 7562 3768 7618 3777
rect 7562 3703 7618 3712
rect 7576 3602 7604 3703
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 7576 2553 7604 2926
rect 7562 2544 7618 2553
rect 7668 2514 7696 3538
rect 7562 2479 7618 2488
rect 7656 2508 7708 2514
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 7288 1012 7340 1018
rect 7288 954 7340 960
rect 7576 480 7604 2479
rect 7656 2450 7708 2456
rect 7760 1986 7788 4247
rect 7840 4218 7892 4224
rect 7852 2922 7880 4218
rect 7944 3913 7972 10152
rect 8036 10130 8064 10202
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8022 9616 8078 9625
rect 8022 9551 8078 9560
rect 8116 9580 8168 9586
rect 8036 9110 8064 9551
rect 8116 9522 8168 9528
rect 8128 9353 8156 9522
rect 8220 9518 8248 10231
rect 8352 9820 8648 9840
rect 8408 9818 8432 9820
rect 8488 9818 8512 9820
rect 8568 9818 8592 9820
rect 8430 9766 8432 9818
rect 8494 9766 8506 9818
rect 8568 9766 8570 9818
rect 8408 9764 8432 9766
rect 8488 9764 8512 9766
rect 8568 9764 8592 9766
rect 8352 9744 8648 9764
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8114 9344 8170 9353
rect 8114 9279 8170 9288
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 8036 4729 8064 9046
rect 8312 8974 8340 9386
rect 8390 9344 8446 9353
rect 8680 9330 8708 10968
rect 8390 9279 8446 9288
rect 8588 9302 8708 9330
rect 8404 9110 8432 9279
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 8300 8968 8352 8974
rect 8588 8956 8616 9302
rect 8666 9208 8722 9217
rect 8666 9143 8722 9152
rect 8680 9110 8708 9143
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8588 8928 8708 8956
rect 8300 8910 8352 8916
rect 8352 8732 8648 8752
rect 8408 8730 8432 8732
rect 8488 8730 8512 8732
rect 8568 8730 8592 8732
rect 8430 8678 8432 8730
rect 8494 8678 8506 8730
rect 8568 8678 8570 8730
rect 8408 8676 8432 8678
rect 8488 8676 8512 8678
rect 8568 8676 8592 8678
rect 8352 8656 8648 8676
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8128 8294 8156 8434
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8128 7478 8156 8230
rect 8312 8090 8340 8230
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8206 7848 8262 7857
rect 8206 7783 8262 7792
rect 8220 7585 8248 7783
rect 8352 7644 8648 7664
rect 8408 7642 8432 7644
rect 8488 7642 8512 7644
rect 8568 7642 8592 7644
rect 8430 7590 8432 7642
rect 8494 7590 8506 7642
rect 8568 7590 8570 7642
rect 8408 7588 8432 7590
rect 8488 7588 8512 7590
rect 8568 7588 8592 7590
rect 8206 7576 8262 7585
rect 8352 7568 8648 7588
rect 8206 7511 8262 7520
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8220 6458 8248 7142
rect 8496 7041 8524 7346
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8482 7032 8538 7041
rect 8392 6996 8444 7002
rect 8588 7002 8616 7210
rect 8482 6967 8538 6976
rect 8576 6996 8628 7002
rect 8392 6938 8444 6944
rect 8576 6938 8628 6944
rect 8404 6866 8432 6938
rect 8680 6905 8708 8928
rect 8666 6896 8722 6905
rect 8392 6860 8444 6866
rect 8666 6831 8722 6840
rect 8392 6802 8444 6808
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8352 6480 8648 6500
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8116 6180 8168 6186
rect 8116 6122 8168 6128
rect 8128 5370 8156 6122
rect 8208 6112 8260 6118
rect 8206 6080 8208 6089
rect 8576 6112 8628 6118
rect 8260 6080 8262 6089
rect 8576 6054 8628 6060
rect 8206 6015 8262 6024
rect 8588 5846 8616 6054
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8300 5636 8352 5642
rect 8220 5596 8300 5624
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8022 4720 8078 4729
rect 8022 4655 8078 4664
rect 7930 3904 7986 3913
rect 7930 3839 7986 3848
rect 7840 2916 7892 2922
rect 7840 2858 7892 2864
rect 7944 2106 7972 3839
rect 8036 2650 8064 4655
rect 8128 4214 8156 5034
rect 8220 4690 8248 5596
rect 8300 5578 8352 5584
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8352 5392 8648 5412
rect 8680 5302 8708 6666
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8312 5086 8616 5114
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 8116 4004 8168 4010
rect 8220 3992 8248 4626
rect 8312 4554 8340 5086
rect 8588 5030 8616 5086
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8482 4856 8538 4865
rect 8482 4791 8538 4800
rect 8496 4554 8524 4791
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8352 4380 8648 4400
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8168 3964 8248 3992
rect 8484 4004 8536 4010
rect 8116 3946 8168 3952
rect 8484 3946 8536 3952
rect 8496 3670 8524 3946
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8588 3380 8616 4150
rect 8680 4078 8708 4490
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8588 3352 8708 3380
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8206 3224 8262 3233
rect 8116 3188 8168 3194
rect 8352 3216 8648 3236
rect 8206 3159 8262 3168
rect 8116 3130 8168 3136
rect 8128 2922 8156 3130
rect 8220 2972 8248 3159
rect 8680 3126 8708 3352
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 8392 2984 8444 2990
rect 8220 2944 8392 2972
rect 8392 2926 8444 2932
rect 8116 2916 8168 2922
rect 8116 2858 8168 2864
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 8574 2544 8630 2553
rect 8574 2479 8630 2488
rect 8588 2446 8616 2479
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8666 2408 8722 2417
rect 7932 2100 7984 2106
rect 7932 2042 7984 2048
rect 7760 1958 7972 1986
rect 7944 480 7972 1958
rect 8128 1902 8156 2382
rect 8772 2394 8800 12600
rect 8850 12472 8906 12481
rect 8850 12407 8852 12416
rect 8904 12407 8906 12416
rect 8852 12378 8904 12384
rect 8850 12064 8906 12073
rect 8850 11999 8906 12008
rect 8864 11762 8892 11999
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8956 11694 8984 14175
rect 9048 11830 9076 16662
rect 9140 16114 9168 17818
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 9140 15162 9168 15914
rect 9232 15434 9260 19520
rect 9404 18488 9456 18494
rect 9404 18430 9456 18436
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9324 16726 9352 17478
rect 9416 17270 9444 18430
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9312 16720 9364 16726
rect 9312 16662 9364 16668
rect 9324 15745 9352 16662
rect 9402 16416 9458 16425
rect 9402 16351 9458 16360
rect 9310 15736 9366 15745
rect 9310 15671 9366 15680
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9232 14346 9260 14962
rect 9324 14822 9352 15506
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9416 14362 9444 16351
rect 9508 16289 9536 17070
rect 9600 17066 9628 19520
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9588 17060 9640 17066
rect 9588 17002 9640 17008
rect 9692 16946 9720 18022
rect 9864 17604 9916 17610
rect 9864 17546 9916 17552
rect 9600 16918 9720 16946
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9600 16833 9628 16918
rect 9586 16824 9642 16833
rect 9586 16759 9642 16768
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9494 16280 9550 16289
rect 9494 16215 9550 16224
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9508 15337 9536 15846
rect 9494 15328 9550 15337
rect 9494 15263 9550 15272
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9324 14334 9444 14362
rect 9128 13320 9180 13326
rect 9232 13308 9260 14282
rect 9324 13705 9352 14334
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9416 13841 9444 14214
rect 9402 13832 9458 13841
rect 9402 13767 9458 13776
rect 9310 13696 9366 13705
rect 9310 13631 9366 13640
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9180 13280 9260 13308
rect 9128 13262 9180 13268
rect 9312 13252 9364 13258
rect 9232 13212 9312 13240
rect 9232 13161 9260 13212
rect 9312 13194 9364 13200
rect 9416 13190 9444 13330
rect 9404 13184 9456 13190
rect 9218 13152 9274 13161
rect 9404 13126 9456 13132
rect 9218 13087 9274 13096
rect 9508 12714 9536 14962
rect 9586 14784 9642 14793
rect 9586 14719 9642 14728
rect 9600 14618 9628 14719
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9600 14113 9628 14418
rect 9586 14104 9642 14113
rect 9586 14039 9642 14048
rect 9692 13938 9720 16594
rect 9784 16522 9812 16934
rect 9876 16522 9904 17546
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 9862 16280 9918 16289
rect 9968 16250 9996 19520
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 9862 16215 9864 16224
rect 9916 16215 9918 16224
rect 9956 16244 10008 16250
rect 9864 16186 9916 16192
rect 9956 16186 10008 16192
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 9784 15473 9812 15574
rect 9770 15464 9826 15473
rect 9770 15399 9826 15408
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9784 15042 9812 15302
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9968 15042 9996 15098
rect 9784 15014 9996 15042
rect 9954 14920 10010 14929
rect 9954 14855 9956 14864
rect 10008 14855 10010 14864
rect 9956 14826 10008 14832
rect 9770 14648 9826 14657
rect 9770 14583 9826 14592
rect 9784 14113 9812 14583
rect 10060 14482 10088 17070
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10152 16833 10180 16934
rect 10138 16824 10194 16833
rect 10138 16759 10194 16768
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10152 15745 10180 16526
rect 10244 16046 10272 17478
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10138 15736 10194 15745
rect 10138 15671 10194 15680
rect 10152 15502 10180 15671
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10140 14816 10192 14822
rect 10138 14784 10140 14793
rect 10192 14784 10194 14793
rect 10138 14719 10194 14728
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9876 14278 9904 14350
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9770 14104 9826 14113
rect 9770 14039 9826 14048
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9600 13530 9628 13670
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 9692 13297 9720 13398
rect 9784 13394 9812 13670
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9678 13288 9734 13297
rect 9678 13223 9734 13232
rect 9862 13288 9918 13297
rect 9862 13223 9918 13232
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9692 12850 9720 13126
rect 9876 12918 9904 13223
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9876 12753 9904 12854
rect 9862 12744 9918 12753
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9680 12708 9732 12714
rect 9862 12679 9918 12688
rect 9680 12650 9732 12656
rect 9310 12608 9366 12617
rect 9140 12566 9310 12594
rect 9140 12442 9168 12566
rect 9310 12543 9366 12552
rect 9310 12472 9366 12481
rect 9128 12436 9180 12442
rect 9310 12407 9312 12416
rect 9128 12378 9180 12384
rect 9364 12407 9366 12416
rect 9588 12436 9640 12442
rect 9312 12378 9364 12384
rect 9588 12378 9640 12384
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 11150 8892 11494
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8942 11112 8998 11121
rect 8942 11047 8998 11056
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8864 9110 8892 10406
rect 8852 9104 8904 9110
rect 8852 9046 8904 9052
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8864 5778 8892 8774
rect 8956 8129 8984 11047
rect 9034 10976 9090 10985
rect 9034 10911 9090 10920
rect 8942 8120 8998 8129
rect 8942 8055 8944 8064
rect 8996 8055 8998 8064
rect 8944 8026 8996 8032
rect 8956 7995 8984 8026
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8956 7002 8984 7822
rect 9048 7750 9076 10911
rect 9140 9518 9168 12038
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 11286 9260 11494
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9232 9722 9260 11086
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9324 10538 9352 11018
rect 9416 10810 9444 12242
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9508 11626 9536 12174
rect 9600 11694 9628 12378
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9600 11529 9628 11630
rect 9586 11520 9642 11529
rect 9586 11455 9642 11464
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9402 10568 9458 10577
rect 9312 10532 9364 10538
rect 9402 10503 9458 10512
rect 9312 10474 9364 10480
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9140 7954 9168 9046
rect 9232 8974 9260 9522
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9232 8265 9260 8366
rect 9218 8256 9274 8265
rect 9218 8191 9274 8200
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9048 7274 9076 7686
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 9128 7268 9180 7274
rect 9128 7210 9180 7216
rect 9140 7177 9168 7210
rect 9126 7168 9182 7177
rect 9126 7103 9182 7112
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8864 5012 8892 5578
rect 8956 5166 8984 6802
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9048 5409 9076 6394
rect 9034 5400 9090 5409
rect 9034 5335 9090 5344
rect 9140 5284 9168 6938
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 6089 9260 6598
rect 9218 6080 9274 6089
rect 9218 6015 9274 6024
rect 9324 5642 9352 10066
rect 9416 9926 9444 10503
rect 9508 9994 9536 11290
rect 9586 10568 9642 10577
rect 9586 10503 9642 10512
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9416 9586 9444 9658
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9600 9353 9628 10503
rect 9692 9382 9720 12650
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9968 12322 9996 13874
rect 10060 12782 10088 14418
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10152 14074 10180 14350
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10140 13456 10192 13462
rect 10138 13424 10140 13433
rect 10192 13424 10194 13433
rect 10138 13359 10194 13368
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10152 12646 10180 12854
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10138 12472 10194 12481
rect 10138 12407 10194 12416
rect 9784 12102 9812 12310
rect 9968 12294 10088 12322
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9770 11656 9826 11665
rect 9770 11591 9826 11600
rect 9784 11558 9812 11591
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 9680 9376 9732 9382
rect 9586 9344 9642 9353
rect 9680 9318 9732 9324
rect 9586 9279 9642 9288
rect 9784 9160 9812 10134
rect 9600 9132 9812 9160
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9416 8809 9444 8978
rect 9600 8922 9628 9132
rect 9876 9042 9904 12106
rect 9968 11937 9996 12174
rect 9954 11928 10010 11937
rect 9954 11863 10010 11872
rect 10060 11762 10088 12294
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10060 11529 10088 11698
rect 10046 11520 10102 11529
rect 10046 11455 10102 11464
rect 10152 11370 10180 12407
rect 10244 12288 10272 15506
rect 10336 13802 10364 19520
rect 10612 17252 10640 19520
rect 10690 17912 10746 17921
rect 10690 17847 10746 17856
rect 10520 17224 10640 17252
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10336 12617 10364 13738
rect 10322 12608 10378 12617
rect 10322 12543 10378 12552
rect 10428 12322 10456 17070
rect 10520 16969 10548 17224
rect 10598 17096 10654 17105
rect 10598 17031 10654 17040
rect 10506 16960 10562 16969
rect 10506 16895 10562 16904
rect 10520 14890 10548 16895
rect 10612 15570 10640 17031
rect 10704 16114 10732 17847
rect 10980 17105 11008 19520
rect 11348 19502 11468 19520
rect 11440 18154 11468 19502
rect 11428 18148 11480 18154
rect 11428 18090 11480 18096
rect 10966 17096 11022 17105
rect 10966 17031 11022 17040
rect 11428 17060 11480 17066
rect 11428 17002 11480 17008
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 10817 16892 11113 16912
rect 10873 16890 10897 16892
rect 10953 16890 10977 16892
rect 11033 16890 11057 16892
rect 10895 16838 10897 16890
rect 10959 16838 10971 16890
rect 11033 16838 11035 16890
rect 10873 16836 10897 16838
rect 10953 16836 10977 16838
rect 11033 16836 11057 16838
rect 10817 16816 11113 16836
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10796 15892 10824 16118
rect 10704 15864 10824 15892
rect 10704 15586 10732 15864
rect 10817 15804 11113 15824
rect 10873 15802 10897 15804
rect 10953 15802 10977 15804
rect 11033 15802 11057 15804
rect 10895 15750 10897 15802
rect 10959 15750 10971 15802
rect 11033 15750 11035 15802
rect 10873 15748 10897 15750
rect 10953 15748 10977 15750
rect 11033 15748 11057 15750
rect 10817 15728 11113 15748
rect 10600 15564 10652 15570
rect 10704 15558 10824 15586
rect 10600 15506 10652 15512
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 10520 13025 10548 14826
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 14249 10640 14758
rect 10704 14498 10732 15438
rect 10796 15201 10824 15558
rect 10782 15192 10838 15201
rect 10966 15192 11022 15201
rect 10782 15127 10838 15136
rect 10876 15156 10928 15162
rect 10928 15136 10966 15144
rect 10928 15127 11022 15136
rect 10928 15116 11008 15127
rect 10876 15098 10928 15104
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 11072 14929 11100 15030
rect 11058 14920 11114 14929
rect 11058 14855 11114 14864
rect 10817 14716 11113 14736
rect 10873 14714 10897 14716
rect 10953 14714 10977 14716
rect 11033 14714 11057 14716
rect 10895 14662 10897 14714
rect 10959 14662 10971 14714
rect 11033 14662 11035 14714
rect 10873 14660 10897 14662
rect 10953 14660 10977 14662
rect 11033 14660 11057 14662
rect 10817 14640 11113 14660
rect 11164 14600 11192 16934
rect 11440 16794 11468 17002
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11256 15638 11284 16186
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11244 15632 11296 15638
rect 11244 15574 11296 15580
rect 11072 14572 11192 14600
rect 10704 14470 11008 14498
rect 10980 14414 11008 14470
rect 10968 14408 11020 14414
rect 10690 14376 10746 14385
rect 10690 14311 10692 14320
rect 10744 14311 10746 14320
rect 10874 14376 10930 14385
rect 10968 14350 11020 14356
rect 10874 14311 10930 14320
rect 10692 14282 10744 14288
rect 10598 14240 10654 14249
rect 10598 14175 10654 14184
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10704 13530 10732 14010
rect 10888 13802 10916 14311
rect 10980 13802 11008 14350
rect 11072 14074 11100 14572
rect 11150 14512 11206 14521
rect 11150 14447 11152 14456
rect 11204 14447 11206 14456
rect 11152 14418 11204 14424
rect 11256 14249 11284 15574
rect 11242 14240 11298 14249
rect 11242 14175 11298 14184
rect 11060 14068 11112 14074
rect 11112 14028 11284 14056
rect 11060 14010 11112 14016
rect 10876 13796 10928 13802
rect 10876 13738 10928 13744
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 10817 13628 11113 13648
rect 10873 13626 10897 13628
rect 10953 13626 10977 13628
rect 11033 13626 11057 13628
rect 10895 13574 10897 13626
rect 10959 13574 10971 13626
rect 11033 13574 11035 13626
rect 10873 13572 10897 13574
rect 10953 13572 10977 13574
rect 11033 13572 11057 13574
rect 10817 13552 11113 13572
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10980 13258 11008 13330
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10506 13016 10562 13025
rect 10506 12951 10562 12960
rect 10612 12940 10824 12968
rect 10612 12730 10640 12940
rect 10520 12702 10640 12730
rect 10796 12714 10824 12940
rect 10980 12918 11008 13194
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 10784 12708 10836 12714
rect 10520 12481 10548 12702
rect 10784 12650 10836 12656
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10506 12472 10562 12481
rect 10506 12407 10562 12416
rect 10428 12294 10548 12322
rect 10244 12260 10364 12288
rect 10230 12200 10286 12209
rect 10230 12135 10286 12144
rect 10244 12102 10272 12135
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10244 11558 10272 11834
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 9968 11354 10180 11370
rect 9956 11348 10180 11354
rect 10008 11342 10180 11348
rect 10230 11384 10286 11393
rect 10230 11319 10286 11328
rect 9956 11290 10008 11296
rect 9954 10296 10010 10305
rect 9954 10231 10010 10240
rect 9968 9897 9996 10231
rect 10244 10198 10272 11319
rect 10232 10192 10284 10198
rect 10232 10134 10284 10140
rect 10336 10044 10364 12260
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10428 11354 10456 12174
rect 10520 12170 10548 12294
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10612 11762 10640 12582
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10704 11608 10732 12582
rect 10817 12540 11113 12560
rect 10873 12538 10897 12540
rect 10953 12538 10977 12540
rect 11033 12538 11057 12540
rect 10895 12486 10897 12538
rect 10959 12486 10971 12538
rect 11033 12486 11035 12538
rect 10873 12484 10897 12486
rect 10953 12484 10977 12486
rect 11033 12484 11057 12486
rect 10817 12464 11113 12484
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10796 11665 10824 12106
rect 10888 11830 10916 12310
rect 10968 12232 11020 12238
rect 11072 12209 11100 12310
rect 10968 12174 11020 12180
rect 11058 12200 11114 12209
rect 10980 11937 11008 12174
rect 11058 12135 11114 12144
rect 10966 11928 11022 11937
rect 10966 11863 11022 11872
rect 10876 11824 10928 11830
rect 10876 11766 10928 11772
rect 10612 11580 10732 11608
rect 10782 11656 10838 11665
rect 10968 11620 11020 11626
rect 10782 11591 10838 11600
rect 10888 11580 10968 11608
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10520 11354 10548 11494
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10612 11150 10640 11580
rect 10888 11540 10916 11580
rect 10968 11562 11020 11568
rect 10704 11512 10916 11540
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10428 10198 10456 10406
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10244 10016 10364 10044
rect 9954 9888 10010 9897
rect 9954 9823 10010 9832
rect 10244 9722 10272 10016
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 9864 9036 9916 9042
rect 9916 8996 9996 9024
rect 9864 8978 9916 8984
rect 9496 8900 9548 8906
rect 9600 8894 9812 8922
rect 9496 8842 9548 8848
rect 9402 8800 9458 8809
rect 9402 8735 9458 8744
rect 9508 8566 9536 8842
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9416 8378 9444 8434
rect 9416 8362 9536 8378
rect 9416 8356 9548 8362
rect 9416 8350 9496 8356
rect 9496 8298 9548 8304
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 7954 9444 8230
rect 9494 8120 9550 8129
rect 9600 8090 9628 8570
rect 9494 8055 9550 8064
rect 9588 8084 9640 8090
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9416 7154 9444 7890
rect 9508 7342 9536 8055
rect 9588 8026 9640 8032
rect 9692 7750 9720 8774
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9416 7126 9536 7154
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 9310 5536 9366 5545
rect 9310 5471 9366 5480
rect 9218 5400 9274 5409
rect 9218 5335 9274 5344
rect 9048 5256 9168 5284
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 8864 4984 8984 5012
rect 9048 5001 9076 5256
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 8864 4622 8892 4694
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8864 3738 8892 4558
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8956 3448 8984 4984
rect 9034 4992 9090 5001
rect 9034 4927 9090 4936
rect 9140 4457 9168 5034
rect 9232 5030 9260 5335
rect 9324 5030 9352 5471
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4604 9352 4966
rect 9416 4865 9444 6734
rect 9508 6186 9536 7126
rect 9784 7018 9812 8894
rect 9862 8800 9918 8809
rect 9862 8735 9918 8744
rect 9876 8634 9904 8735
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9876 8090 9904 8230
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9876 7206 9904 7414
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9784 6990 9904 7018
rect 9772 6928 9824 6934
rect 9678 6896 9734 6905
rect 9772 6870 9824 6876
rect 9678 6831 9734 6840
rect 9692 6798 9720 6831
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9586 6352 9642 6361
rect 9586 6287 9642 6296
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9600 5817 9628 6287
rect 9692 5953 9720 6598
rect 9784 6458 9812 6870
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9678 5944 9734 5953
rect 9678 5879 9734 5888
rect 9772 5840 9824 5846
rect 9586 5808 9642 5817
rect 9876 5817 9904 6990
rect 9772 5782 9824 5788
rect 9862 5808 9918 5817
rect 9586 5743 9642 5752
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9402 4856 9458 4865
rect 9402 4791 9458 4800
rect 9404 4752 9456 4758
rect 9508 4740 9536 5034
rect 9678 4856 9734 4865
rect 9600 4814 9678 4842
rect 9600 4758 9628 4814
rect 9678 4791 9734 4800
rect 9456 4712 9536 4740
rect 9588 4752 9640 4758
rect 9404 4694 9456 4700
rect 9588 4694 9640 4700
rect 9324 4576 9444 4604
rect 9126 4448 9182 4457
rect 9126 4383 9182 4392
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9232 3942 9260 4218
rect 9324 4146 9352 4218
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9416 4026 9444 4576
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9586 4176 9642 4185
rect 9586 4111 9642 4120
rect 9324 3998 9444 4026
rect 9036 3936 9088 3942
rect 9220 3936 9272 3942
rect 9088 3896 9168 3924
rect 9036 3878 9088 3884
rect 9140 3602 9168 3896
rect 9220 3878 9272 3884
rect 9324 3618 9352 3998
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9232 3590 9352 3618
rect 9508 3602 9536 3878
rect 9496 3596 9548 3602
rect 9232 3482 9260 3590
rect 9496 3538 9548 3544
rect 8936 3420 8984 3448
rect 9140 3454 9260 3482
rect 8850 3360 8906 3369
rect 8936 3346 8964 3420
rect 9034 3360 9090 3369
rect 8936 3318 9034 3346
rect 8850 3295 8906 3304
rect 9034 3295 9090 3304
rect 8864 2938 8892 3295
rect 8864 2910 8984 2938
rect 8956 2854 8984 2910
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 8864 2417 8892 2790
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 8722 2366 8800 2394
rect 8850 2408 8906 2417
rect 8666 2343 8722 2352
rect 8850 2343 8906 2352
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 9048 2145 9076 2450
rect 9034 2136 9090 2145
rect 8944 2100 8996 2106
rect 9034 2071 9090 2080
rect 8944 2042 8996 2048
rect 8576 2032 8628 2038
rect 8576 1974 8628 1980
rect 8116 1896 8168 1902
rect 8116 1838 8168 1844
rect 8208 1556 8260 1562
rect 8208 1498 8260 1504
rect 8220 480 8248 1498
rect 8588 480 8616 1974
rect 8956 480 8984 2042
rect 9048 1698 9076 2071
rect 9140 2038 9168 3454
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9494 3360 9550 3369
rect 9232 2922 9260 3334
rect 9494 3295 9550 3304
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 9218 2680 9274 2689
rect 9218 2615 9274 2624
rect 9128 2032 9180 2038
rect 9128 1974 9180 1980
rect 9036 1692 9088 1698
rect 9036 1634 9088 1640
rect 9232 480 9260 2615
rect 9324 2446 9352 2994
rect 9508 2514 9536 3295
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9324 2038 9352 2246
rect 9312 2032 9364 2038
rect 9312 1974 9364 1980
rect 9324 1834 9352 1974
rect 9312 1828 9364 1834
rect 9312 1770 9364 1776
rect 9600 480 9628 4111
rect 9692 4010 9720 4422
rect 9784 4214 9812 5782
rect 9862 5743 9918 5752
rect 9968 5234 9996 8996
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10060 7188 10088 8434
rect 10152 7410 10180 9046
rect 10244 8430 10272 9658
rect 10428 9586 10456 9930
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10336 9110 10364 9318
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10244 7342 10272 7686
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10060 7160 10272 7188
rect 10046 7032 10102 7041
rect 10046 6967 10048 6976
rect 10100 6967 10102 6976
rect 10048 6938 10100 6944
rect 10140 6928 10192 6934
rect 10138 6896 10140 6905
rect 10192 6896 10194 6905
rect 10138 6831 10194 6840
rect 10140 6792 10192 6798
rect 10244 6769 10272 7160
rect 10140 6734 10192 6740
rect 10230 6760 10286 6769
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10060 5681 10088 5850
rect 10046 5672 10102 5681
rect 10046 5607 10102 5616
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 10152 5114 10180 6734
rect 10230 6695 10286 6704
rect 10336 6633 10364 9046
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10428 8498 10456 8910
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10428 8129 10456 8298
rect 10414 8120 10470 8129
rect 10414 8055 10470 8064
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10428 7002 10456 7346
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10520 6882 10548 10406
rect 10704 10198 10732 11512
rect 10817 11452 11113 11472
rect 10873 11450 10897 11452
rect 10953 11450 10977 11452
rect 11033 11450 11057 11452
rect 10895 11398 10897 11450
rect 10959 11398 10971 11450
rect 11033 11398 11035 11450
rect 10873 11396 10897 11398
rect 10953 11396 10977 11398
rect 11033 11396 11057 11398
rect 10817 11376 11113 11396
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10980 11082 11008 11154
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10782 10840 10838 10849
rect 10782 10775 10838 10784
rect 10796 10674 10824 10775
rect 10980 10674 11008 11018
rect 11072 10810 11100 11154
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10817 10364 11113 10384
rect 10873 10362 10897 10364
rect 10953 10362 10977 10364
rect 11033 10362 11057 10364
rect 10895 10310 10897 10362
rect 10959 10310 10971 10362
rect 11033 10310 11035 10362
rect 10873 10308 10897 10310
rect 10953 10308 10977 10310
rect 11033 10308 11057 10310
rect 10817 10288 11113 10308
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 11072 9761 11100 9998
rect 11058 9752 11114 9761
rect 11058 9687 11114 9696
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10612 8838 10640 9522
rect 11164 9518 11192 13670
rect 11256 11694 11284 14028
rect 11348 12617 11376 15982
rect 11440 15910 11468 16390
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11334 12608 11390 12617
rect 11334 12543 11390 12552
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11244 11552 11296 11558
rect 11242 11520 11244 11529
rect 11296 11520 11298 11529
rect 11242 11455 11298 11464
rect 11242 11384 11298 11393
rect 11348 11354 11376 11766
rect 11242 11319 11298 11328
rect 11336 11348 11388 11354
rect 11256 10985 11284 11319
rect 11336 11290 11388 11296
rect 11242 10976 11298 10985
rect 11440 10962 11468 15506
rect 11532 15026 11560 16594
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11532 12442 11560 14962
rect 11624 12617 11652 19520
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 11716 16425 11744 17002
rect 11702 16416 11758 16425
rect 11702 16351 11758 16360
rect 11808 15570 11836 17478
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 16658 11928 16934
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11794 15464 11850 15473
rect 11716 14822 11744 15438
rect 11794 15399 11796 15408
rect 11848 15399 11850 15408
rect 11796 15370 11848 15376
rect 11794 15056 11850 15065
rect 11794 14991 11796 15000
rect 11848 14991 11850 15000
rect 11796 14962 11848 14968
rect 11704 14816 11756 14822
rect 11702 14784 11704 14793
rect 11756 14784 11758 14793
rect 11702 14719 11758 14728
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 13530 11744 14214
rect 11808 13977 11836 14418
rect 11794 13968 11850 13977
rect 11794 13903 11850 13912
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11716 12850 11744 13330
rect 11796 13320 11848 13326
rect 11794 13288 11796 13297
rect 11848 13288 11850 13297
rect 11794 13223 11850 13232
rect 11794 13152 11850 13161
rect 11794 13087 11850 13096
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11808 12782 11836 13087
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11610 12608 11666 12617
rect 11610 12543 11666 12552
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11518 12336 11574 12345
rect 11794 12336 11850 12345
rect 11518 12271 11574 12280
rect 11704 12300 11756 12306
rect 11532 12238 11560 12271
rect 11900 12306 11928 15914
rect 11992 12617 12020 19520
rect 12072 18148 12124 18154
rect 12072 18090 12124 18096
rect 12084 16658 12112 18090
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 12072 15972 12124 15978
rect 12072 15914 12124 15920
rect 11978 12608 12034 12617
rect 11978 12543 12034 12552
rect 11978 12472 12034 12481
rect 11978 12407 12034 12416
rect 11794 12271 11850 12280
rect 11888 12300 11940 12306
rect 11704 12242 11756 12248
rect 11520 12232 11572 12238
rect 11716 12209 11744 12242
rect 11520 12174 11572 12180
rect 11702 12200 11758 12209
rect 11612 12164 11664 12170
rect 11702 12135 11758 12144
rect 11612 12106 11664 12112
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11532 11830 11560 12038
rect 11520 11824 11572 11830
rect 11520 11766 11572 11772
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11242 10911 11298 10920
rect 11348 10934 11468 10962
rect 11244 10124 11296 10130
rect 11348 10112 11376 10934
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11296 10084 11376 10112
rect 11244 10066 11296 10072
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10598 8120 10654 8129
rect 10598 8055 10654 8064
rect 10612 7857 10640 8055
rect 10598 7848 10654 7857
rect 10598 7783 10654 7792
rect 10704 7800 10732 9386
rect 10817 9276 11113 9296
rect 10873 9274 10897 9276
rect 10953 9274 10977 9276
rect 11033 9274 11057 9276
rect 10895 9222 10897 9274
rect 10959 9222 10971 9274
rect 11033 9222 11035 9274
rect 10873 9220 10897 9222
rect 10953 9220 10977 9222
rect 11033 9220 11057 9222
rect 10817 9200 11113 9220
rect 11256 9160 11284 10066
rect 11334 9752 11390 9761
rect 11334 9687 11336 9696
rect 11388 9687 11390 9696
rect 11336 9658 11388 9664
rect 11440 9518 11468 10202
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11532 9382 11560 11630
rect 11624 11082 11652 12106
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11716 11286 11744 11834
rect 11808 11354 11836 12271
rect 11888 12242 11940 12248
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11716 10742 11744 10950
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11624 10062 11652 10610
rect 11704 10600 11756 10606
rect 11702 10568 11704 10577
rect 11756 10568 11758 10577
rect 11702 10503 11758 10512
rect 11702 10432 11758 10441
rect 11702 10367 11758 10376
rect 11716 10130 11744 10367
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11704 9920 11756 9926
rect 11702 9888 11704 9897
rect 11756 9888 11758 9897
rect 11702 9823 11758 9832
rect 11612 9716 11664 9722
rect 11808 9704 11836 11086
rect 11612 9658 11664 9664
rect 11716 9676 11836 9704
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11348 9178 11376 9318
rect 11164 9132 11284 9160
rect 11336 9172 11388 9178
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10796 8430 10824 8842
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10980 8362 11008 8774
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10817 8188 11113 8208
rect 10873 8186 10897 8188
rect 10953 8186 10977 8188
rect 11033 8186 11057 8188
rect 10895 8134 10897 8186
rect 10959 8134 10971 8186
rect 11033 8134 11035 8186
rect 10873 8132 10897 8134
rect 10953 8132 10977 8134
rect 11033 8132 11057 8134
rect 10817 8112 11113 8132
rect 11164 7970 11192 9132
rect 11336 9114 11388 9120
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11256 8634 11284 8978
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11428 8560 11480 8566
rect 11242 8528 11298 8537
rect 11532 8548 11560 8910
rect 11480 8520 11560 8548
rect 11428 8502 11480 8508
rect 11242 8463 11244 8472
rect 11296 8463 11298 8472
rect 11244 8434 11296 8440
rect 11426 8392 11482 8401
rect 11426 8327 11482 8336
rect 11520 8356 11572 8362
rect 11440 8090 11468 8327
rect 11520 8298 11572 8304
rect 11532 8090 11560 8298
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11072 7942 11192 7970
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10704 7772 10916 7800
rect 10600 7744 10652 7750
rect 10598 7712 10600 7721
rect 10652 7712 10654 7721
rect 10598 7647 10654 7656
rect 10782 7712 10838 7721
rect 10782 7647 10838 7656
rect 10796 7562 10824 7647
rect 10428 6866 10548 6882
rect 10416 6860 10548 6866
rect 10468 6854 10548 6860
rect 10612 7534 10824 7562
rect 10416 6802 10468 6808
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10322 6624 10378 6633
rect 10322 6559 10378 6568
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10244 5370 10272 6258
rect 10336 6254 10364 6394
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10520 6089 10548 6734
rect 10612 6254 10640 7534
rect 10888 7324 10916 7772
rect 10980 7478 11008 7822
rect 11072 7546 11100 7942
rect 11428 7880 11480 7886
rect 11150 7848 11206 7857
rect 11428 7822 11480 7828
rect 11150 7783 11206 7792
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11164 7478 11192 7783
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 10888 7296 11284 7324
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 10817 7100 11113 7120
rect 10873 7098 10897 7100
rect 10953 7098 10977 7100
rect 11033 7098 11057 7100
rect 10895 7046 10897 7098
rect 10959 7046 10971 7098
rect 11033 7046 11035 7098
rect 10873 7044 10897 7046
rect 10953 7044 10977 7046
rect 11033 7044 11057 7046
rect 10817 7024 11113 7044
rect 10968 6860 11020 6866
rect 11164 6848 11192 7142
rect 10968 6802 11020 6808
rect 11072 6820 11192 6848
rect 10980 6254 11008 6802
rect 11072 6730 11100 6820
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10692 6112 10744 6118
rect 10506 6080 10562 6089
rect 11164 6100 11192 6666
rect 10744 6072 11192 6100
rect 10692 6054 10744 6060
rect 10506 6015 10562 6024
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 11060 5840 11112 5846
rect 10966 5808 11022 5817
rect 10508 5772 10560 5778
rect 10784 5772 10836 5778
rect 10508 5714 10560 5720
rect 10704 5732 10784 5760
rect 10520 5681 10548 5714
rect 10506 5672 10562 5681
rect 10506 5607 10562 5616
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10152 5086 10272 5114
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 9862 4856 9918 4865
rect 10060 4826 10088 4966
rect 9862 4791 9918 4800
rect 10048 4820 10100 4826
rect 9876 4622 9904 4791
rect 10048 4762 10100 4768
rect 9956 4752 10008 4758
rect 9956 4694 10008 4700
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9968 3738 9996 4694
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10060 4146 10088 4558
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10048 3936 10100 3942
rect 10046 3904 10048 3913
rect 10100 3904 10102 3913
rect 10046 3839 10102 3848
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9692 3448 9720 3674
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 9692 3420 9812 3448
rect 9784 3380 9812 3420
rect 10060 3398 10088 3470
rect 10048 3392 10100 3398
rect 9678 3360 9734 3369
rect 9784 3352 9904 3380
rect 9678 3295 9734 3304
rect 9692 2650 9720 3295
rect 9772 3120 9824 3126
rect 9770 3088 9772 3097
rect 9824 3088 9826 3097
rect 9770 3023 9826 3032
rect 9876 2854 9904 3352
rect 10048 3334 10100 3340
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10060 2990 10088 3062
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 9864 2848 9916 2854
rect 10048 2848 10100 2854
rect 9864 2790 9916 2796
rect 10046 2816 10048 2825
rect 10100 2816 10102 2825
rect 10046 2751 10102 2760
rect 9954 2680 10010 2689
rect 9680 2644 9732 2650
rect 10152 2650 10180 4966
rect 10244 4282 10272 5086
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 10244 3913 10272 4014
rect 10230 3904 10286 3913
rect 10230 3839 10286 3848
rect 10230 3768 10286 3777
rect 10230 3703 10286 3712
rect 9954 2615 10010 2624
rect 10140 2644 10192 2650
rect 9680 2586 9732 2592
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9784 1834 9812 2246
rect 9772 1828 9824 1834
rect 9772 1770 9824 1776
rect 9968 480 9996 2615
rect 10140 2586 10192 2592
rect 10244 2106 10272 3703
rect 10336 2650 10364 4422
rect 10428 3777 10456 5510
rect 10520 5409 10548 5607
rect 10506 5400 10562 5409
rect 10506 5335 10562 5344
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10414 3768 10470 3777
rect 10414 3703 10470 3712
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10428 3058 10456 3538
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10520 2904 10548 5170
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10428 2876 10548 2904
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10428 2378 10456 2876
rect 10416 2372 10468 2378
rect 10416 2314 10468 2320
rect 10232 2100 10284 2106
rect 10232 2042 10284 2048
rect 10324 1896 10376 1902
rect 10324 1838 10376 1844
rect 10336 480 10364 1838
rect 10612 480 10640 5102
rect 10704 4078 10732 5732
rect 11060 5782 11112 5788
rect 10966 5743 11022 5752
rect 10784 5714 10836 5720
rect 10980 5098 11008 5743
rect 11072 5642 11100 5782
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11072 5234 11100 5306
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10817 4848 11113 4868
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10796 4010 10824 4558
rect 10980 4486 11008 4626
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 11072 4010 11100 4694
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 11164 3602 11192 5510
rect 11256 5166 11284 7296
rect 11348 6066 11376 7482
rect 11440 6798 11468 7822
rect 11624 6934 11652 9658
rect 11716 8838 11744 9676
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11716 7750 11744 7958
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11716 7410 11744 7482
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11612 6928 11664 6934
rect 11610 6896 11612 6905
rect 11664 6896 11666 6905
rect 11610 6831 11666 6840
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11428 6792 11480 6798
rect 11612 6792 11664 6798
rect 11428 6734 11480 6740
rect 11610 6760 11612 6769
rect 11664 6760 11666 6769
rect 11610 6695 11666 6704
rect 11610 6624 11666 6633
rect 11610 6559 11666 6568
rect 11348 6038 11560 6066
rect 11334 5944 11390 5953
rect 11334 5879 11336 5888
rect 11388 5879 11390 5888
rect 11336 5850 11388 5856
rect 11334 5536 11390 5545
rect 11334 5471 11390 5480
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11242 4992 11298 5001
rect 11242 4927 11298 4936
rect 11256 4826 11284 4927
rect 11348 4826 11376 5471
rect 11532 5370 11560 6038
rect 11624 5778 11652 6559
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11428 5296 11480 5302
rect 11716 5250 11744 6802
rect 11428 5238 11480 5244
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11256 4282 11284 4626
rect 11334 4312 11390 4321
rect 11244 4276 11296 4282
rect 11440 4282 11468 5238
rect 11532 5222 11744 5250
rect 11532 5137 11560 5222
rect 11612 5160 11664 5166
rect 11518 5128 11574 5137
rect 11612 5102 11664 5108
rect 11518 5063 11574 5072
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11334 4247 11390 4256
rect 11428 4276 11480 4282
rect 11244 4218 11296 4224
rect 11348 4146 11376 4247
rect 11428 4218 11480 4224
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11440 4026 11468 4218
rect 11348 3998 11468 4026
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11256 3738 11284 3878
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10704 2582 10732 3402
rect 10796 3369 10824 3470
rect 10782 3360 10838 3369
rect 10782 3295 10838 3304
rect 10782 3224 10838 3233
rect 10888 3210 10916 3470
rect 10838 3182 10916 3210
rect 10782 3159 10838 3168
rect 10796 3126 10824 3159
rect 10784 3120 10836 3126
rect 11256 3097 11284 3538
rect 10784 3062 10836 3068
rect 11242 3088 11298 3097
rect 10968 3052 11020 3058
rect 11242 3023 11298 3032
rect 10968 2994 11020 3000
rect 10980 2922 11008 2994
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10817 2672 11113 2692
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 11348 2446 11376 3998
rect 11426 3904 11482 3913
rect 11426 3839 11482 3848
rect 11440 3398 11468 3839
rect 11428 3392 11480 3398
rect 11428 3334 11480 3340
rect 11426 3088 11482 3097
rect 11426 3023 11482 3032
rect 11440 2854 11468 3023
rect 11532 2990 11560 4626
rect 11624 4622 11652 5102
rect 11808 5098 11836 9318
rect 11900 5914 11928 12242
rect 11992 8129 12020 12407
rect 12084 10266 12112 15914
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12070 10160 12126 10169
rect 12070 10095 12126 10104
rect 12084 10062 12112 10095
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12070 9888 12126 9897
rect 12070 9823 12126 9832
rect 11978 8120 12034 8129
rect 11978 8055 12034 8064
rect 12084 7954 12112 9823
rect 12176 9722 12204 16662
rect 12268 16561 12296 16730
rect 12254 16552 12310 16561
rect 12254 16487 12310 16496
rect 12360 16250 12388 19520
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12348 16040 12400 16046
rect 12254 16008 12310 16017
rect 12348 15982 12400 15988
rect 12254 15943 12310 15952
rect 12268 15706 12296 15943
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12268 13410 12296 15506
rect 12360 13870 12388 15982
rect 12452 15337 12480 16594
rect 12438 15328 12494 15337
rect 12438 15263 12494 15272
rect 12440 14952 12492 14958
rect 12438 14920 12440 14929
rect 12492 14920 12494 14929
rect 12438 14855 12494 14864
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12348 13864 12400 13870
rect 12452 13841 12480 14758
rect 12348 13806 12400 13812
rect 12438 13832 12494 13841
rect 12438 13767 12494 13776
rect 12544 13716 12572 17070
rect 12452 13688 12572 13716
rect 12268 13382 12388 13410
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12268 12850 12296 13262
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12360 12594 12388 13382
rect 12268 12566 12388 12594
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12268 9518 12296 12566
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12360 10538 12388 12378
rect 12452 12209 12480 13688
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 12544 12442 12572 13330
rect 12636 12753 12664 19520
rect 12808 17944 12860 17950
rect 12808 17886 12860 17892
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12728 16266 12756 17614
rect 12820 16522 12848 17886
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12728 16238 12848 16266
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12728 14113 12756 14418
rect 12714 14104 12770 14113
rect 12714 14039 12770 14048
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12622 12744 12678 12753
rect 12728 12714 12756 13806
rect 12622 12679 12678 12688
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12714 12608 12770 12617
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12530 12336 12586 12345
rect 12530 12271 12586 12280
rect 12438 12200 12494 12209
rect 12438 12135 12494 12144
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12452 11014 12480 12038
rect 12544 11694 12572 12271
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12636 11286 12664 12582
rect 12714 12543 12770 12552
rect 12728 11665 12756 12543
rect 12820 12458 12848 16238
rect 12912 16182 12940 16934
rect 12900 16176 12952 16182
rect 12900 16118 12952 16124
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12912 13977 12940 15438
rect 12898 13968 12954 13977
rect 12898 13903 12954 13912
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12912 12617 12940 13670
rect 12898 12608 12954 12617
rect 12898 12543 12954 12552
rect 12820 12430 12940 12458
rect 12808 12096 12860 12102
rect 12806 12064 12808 12073
rect 12860 12064 12862 12073
rect 12806 11999 12862 12008
rect 12912 11898 12940 12430
rect 12900 11892 12952 11898
rect 13004 11880 13032 19520
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 13096 13530 13124 17070
rect 13188 15144 13216 17750
rect 13372 17649 13400 19520
rect 13358 17640 13414 17649
rect 13358 17575 13414 17584
rect 13282 17436 13578 17456
rect 13338 17434 13362 17436
rect 13418 17434 13442 17436
rect 13498 17434 13522 17436
rect 13360 17382 13362 17434
rect 13424 17382 13436 17434
rect 13498 17382 13500 17434
rect 13338 17380 13362 17382
rect 13418 17380 13442 17382
rect 13498 17380 13522 17382
rect 13282 17360 13578 17380
rect 13740 16833 13768 19520
rect 13912 18012 13964 18018
rect 13912 17954 13964 17960
rect 13726 16824 13782 16833
rect 13726 16759 13782 16768
rect 13924 16697 13952 17954
rect 13726 16688 13782 16697
rect 13726 16623 13782 16632
rect 13910 16688 13966 16697
rect 13910 16623 13966 16632
rect 13282 16348 13578 16368
rect 13338 16346 13362 16348
rect 13418 16346 13442 16348
rect 13498 16346 13522 16348
rect 13360 16294 13362 16346
rect 13424 16294 13436 16346
rect 13498 16294 13500 16346
rect 13338 16292 13362 16294
rect 13418 16292 13442 16294
rect 13498 16292 13522 16294
rect 13282 16272 13578 16292
rect 13282 15260 13578 15280
rect 13338 15258 13362 15260
rect 13418 15258 13442 15260
rect 13498 15258 13522 15260
rect 13360 15206 13362 15258
rect 13424 15206 13436 15258
rect 13498 15206 13500 15258
rect 13338 15204 13362 15206
rect 13418 15204 13442 15206
rect 13498 15204 13522 15206
rect 13282 15184 13578 15204
rect 13188 15116 13308 15144
rect 13174 15056 13230 15065
rect 13174 14991 13230 15000
rect 13188 13530 13216 14991
rect 13280 14618 13308 15116
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13282 14172 13578 14192
rect 13338 14170 13362 14172
rect 13418 14170 13442 14172
rect 13498 14170 13522 14172
rect 13360 14118 13362 14170
rect 13424 14118 13436 14170
rect 13498 14118 13500 14170
rect 13338 14116 13362 14118
rect 13418 14116 13442 14118
rect 13498 14116 13522 14118
rect 13282 14096 13578 14116
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13096 12170 13124 13466
rect 13280 13326 13308 13874
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13282 13084 13578 13104
rect 13338 13082 13362 13084
rect 13418 13082 13442 13084
rect 13498 13082 13522 13084
rect 13360 13030 13362 13082
rect 13424 13030 13436 13082
rect 13498 13030 13500 13082
rect 13338 13028 13362 13030
rect 13418 13028 13442 13030
rect 13498 13028 13522 13030
rect 13282 13008 13578 13028
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13280 12753 13308 12854
rect 13648 12850 13676 14418
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13266 12744 13322 12753
rect 13176 12708 13228 12714
rect 13740 12730 13768 16623
rect 14016 15586 14044 19520
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14292 16794 14320 17682
rect 14384 17542 14412 19520
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 14108 16561 14136 16594
rect 14094 16552 14150 16561
rect 14094 16487 14150 16496
rect 14016 15558 14320 15586
rect 14004 15496 14056 15502
rect 13818 15464 13874 15473
rect 14004 15438 14056 15444
rect 13818 15399 13874 15408
rect 13832 13870 13860 15399
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13266 12679 13322 12688
rect 13648 12702 13768 12730
rect 13176 12650 13228 12656
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 13004 11852 13124 11880
rect 12900 11834 12952 11840
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12714 11656 12770 11665
rect 12714 11591 12770 11600
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12728 11370 12756 11494
rect 12728 11342 12848 11370
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12360 9897 12388 10474
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12346 9888 12402 9897
rect 12346 9823 12402 9832
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12164 8968 12216 8974
rect 12268 8945 12296 9318
rect 12164 8910 12216 8916
rect 12254 8936 12310 8945
rect 12176 8673 12204 8910
rect 12254 8871 12310 8880
rect 12162 8664 12218 8673
rect 12162 8599 12218 8608
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12072 7948 12124 7954
rect 11992 7908 12072 7936
rect 11992 7177 12020 7908
rect 12072 7890 12124 7896
rect 12176 7818 12204 8502
rect 12360 8265 12388 9590
rect 12452 9489 12480 10406
rect 12636 10146 12664 10950
rect 12544 10118 12664 10146
rect 12438 9480 12494 9489
rect 12438 9415 12494 9424
rect 12438 9208 12494 9217
rect 12438 9143 12494 9152
rect 12452 9042 12480 9143
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12440 8832 12492 8838
rect 12544 8809 12572 10118
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 9761 12664 9998
rect 12622 9752 12678 9761
rect 12622 9687 12678 9696
rect 12728 9654 12756 11222
rect 12820 9654 12848 11342
rect 13004 11121 13032 11698
rect 13096 11393 13124 11852
rect 13082 11384 13138 11393
rect 13082 11319 13138 11328
rect 13188 11286 13216 12650
rect 13282 11996 13578 12016
rect 13338 11994 13362 11996
rect 13418 11994 13442 11996
rect 13498 11994 13522 11996
rect 13360 11942 13362 11994
rect 13424 11942 13436 11994
rect 13498 11942 13500 11994
rect 13338 11940 13362 11942
rect 13418 11940 13442 11942
rect 13498 11940 13522 11942
rect 13282 11920 13578 11940
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12990 11112 13046 11121
rect 12900 11076 12952 11082
rect 12990 11047 13046 11056
rect 12900 11018 12952 11024
rect 12912 10962 12940 11018
rect 12912 10934 13032 10962
rect 12900 10192 12952 10198
rect 12898 10160 12900 10169
rect 12952 10160 12954 10169
rect 12898 10095 12954 10104
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12440 8774 12492 8780
rect 12530 8800 12586 8809
rect 12452 8548 12480 8774
rect 12530 8735 12586 8744
rect 12452 8520 12572 8548
rect 12438 8392 12494 8401
rect 12438 8327 12494 8336
rect 12346 8256 12402 8265
rect 12346 8191 12402 8200
rect 12346 7984 12402 7993
rect 12256 7948 12308 7954
rect 12452 7954 12480 8327
rect 12346 7919 12402 7928
rect 12440 7948 12492 7954
rect 12256 7890 12308 7896
rect 12268 7857 12296 7890
rect 12254 7848 12310 7857
rect 12164 7812 12216 7818
rect 12360 7834 12388 7919
rect 12440 7890 12492 7896
rect 12544 7886 12572 8520
rect 12636 8498 12664 9522
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12532 7880 12584 7886
rect 12360 7806 12480 7834
rect 12532 7822 12584 7828
rect 12254 7783 12310 7792
rect 12164 7754 12216 7760
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11978 7168 12034 7177
rect 11978 7103 12034 7112
rect 11978 6760 12034 6769
rect 11978 6695 12034 6704
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11796 5092 11848 5098
rect 11796 5034 11848 5040
rect 11794 4992 11850 5001
rect 11794 4927 11850 4936
rect 11808 4690 11836 4927
rect 11900 4758 11928 5306
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11612 4004 11664 4010
rect 11612 3946 11664 3952
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11426 2680 11482 2689
rect 11426 2615 11428 2624
rect 11480 2615 11482 2624
rect 11428 2586 11480 2592
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11336 2304 11388 2310
rect 10966 2272 11022 2281
rect 11336 2246 11388 2252
rect 10966 2207 11022 2216
rect 10980 480 11008 2207
rect 11348 480 11376 2246
rect 11440 1562 11468 2586
rect 11428 1556 11480 1562
rect 11428 1498 11480 1504
rect 11624 480 11652 3946
rect 11716 3534 11744 4558
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11900 4146 11928 4422
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11808 3126 11836 3878
rect 11900 3534 11928 4082
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11808 2145 11836 2926
rect 11794 2136 11850 2145
rect 11794 2071 11850 2080
rect 11992 480 12020 6695
rect 12084 3738 12112 7346
rect 12176 5846 12204 7754
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12268 7002 12296 7686
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12360 7002 12388 7142
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12254 6896 12310 6905
rect 12254 6831 12310 6840
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12176 5234 12204 5646
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12176 4185 12204 4218
rect 12162 4176 12218 4185
rect 12162 4111 12218 4120
rect 12162 3904 12218 3913
rect 12162 3839 12218 3848
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12176 2582 12204 3839
rect 12268 3618 12296 6831
rect 12452 6458 12480 7806
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12544 7410 12572 7686
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12636 6882 12664 8298
rect 12728 8022 12756 9454
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12820 9353 12848 9386
rect 12806 9344 12862 9353
rect 12806 9279 12862 9288
rect 12912 9194 12940 9998
rect 12820 9166 12940 9194
rect 12820 8974 12848 9166
rect 13004 9058 13032 10934
rect 13096 10674 13124 11154
rect 13280 11098 13308 11630
rect 13648 11354 13676 12702
rect 13726 11792 13782 11801
rect 13726 11727 13782 11736
rect 13740 11694 13768 11727
rect 13832 11694 13860 13806
rect 13910 13424 13966 13433
rect 13910 13359 13912 13368
rect 13964 13359 13966 13368
rect 13912 13330 13964 13336
rect 13910 13016 13966 13025
rect 13910 12951 13966 12960
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13740 11286 13768 11630
rect 13924 11626 13952 12951
rect 13912 11620 13964 11626
rect 13912 11562 13964 11568
rect 13728 11280 13780 11286
rect 13634 11248 13690 11257
rect 13728 11222 13780 11228
rect 13634 11183 13690 11192
rect 13188 11070 13308 11098
rect 13542 11112 13598 11121
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13096 9586 13124 10474
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 13096 9353 13124 9386
rect 13082 9344 13138 9353
rect 13082 9279 13138 9288
rect 13188 9178 13216 11070
rect 13542 11047 13544 11056
rect 13596 11047 13598 11056
rect 13544 11018 13596 11024
rect 13282 10908 13578 10928
rect 13338 10906 13362 10908
rect 13418 10906 13442 10908
rect 13498 10906 13522 10908
rect 13360 10854 13362 10906
rect 13424 10854 13436 10906
rect 13498 10854 13500 10906
rect 13338 10852 13362 10854
rect 13418 10852 13442 10854
rect 13498 10852 13522 10854
rect 13282 10832 13578 10852
rect 13282 9820 13578 9840
rect 13338 9818 13362 9820
rect 13418 9818 13442 9820
rect 13498 9818 13522 9820
rect 13360 9766 13362 9818
rect 13424 9766 13436 9818
rect 13498 9766 13500 9818
rect 13338 9764 13362 9766
rect 13418 9764 13442 9766
rect 13498 9764 13522 9766
rect 13282 9744 13578 9764
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 12912 9030 13032 9058
rect 13176 9036 13228 9042
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12820 7886 12848 8434
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12716 7472 12768 7478
rect 12820 7449 12848 7686
rect 12716 7414 12768 7420
rect 12806 7440 12862 7449
rect 12728 7324 12756 7414
rect 12912 7410 12940 9030
rect 13176 8978 13228 8984
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 13004 7546 13032 8910
rect 13188 8537 13216 8978
rect 13282 8732 13578 8752
rect 13338 8730 13362 8732
rect 13418 8730 13442 8732
rect 13498 8730 13522 8732
rect 13360 8678 13362 8730
rect 13424 8678 13436 8730
rect 13498 8678 13500 8730
rect 13338 8676 13362 8678
rect 13418 8676 13442 8678
rect 13498 8676 13522 8678
rect 13282 8656 13578 8676
rect 13648 8634 13676 11183
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13740 10266 13768 11086
rect 13820 10736 13872 10742
rect 13818 10704 13820 10713
rect 13872 10704 13874 10713
rect 13818 10639 13874 10648
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13832 10062 13860 10542
rect 13924 10130 13952 11562
rect 14016 10606 14044 15438
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13820 10056 13872 10062
rect 13740 10016 13820 10044
rect 13740 9654 13768 10016
rect 13820 9998 13872 10004
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13740 8974 13768 9590
rect 13832 9110 13860 9658
rect 13910 9616 13966 9625
rect 13910 9551 13966 9560
rect 13924 9518 13952 9551
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13360 8560 13412 8566
rect 13174 8528 13230 8537
rect 13360 8502 13412 8508
rect 13174 8463 13230 8472
rect 13372 8090 13400 8502
rect 13740 8498 13768 8910
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13452 8424 13504 8430
rect 13504 8401 13584 8412
rect 13504 8392 13598 8401
rect 13504 8384 13542 8392
rect 13452 8366 13504 8372
rect 13542 8327 13598 8336
rect 13728 8356 13780 8362
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 13004 7410 13032 7482
rect 12806 7375 12862 7384
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12728 7296 12848 7324
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12544 6854 12664 6882
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12544 6322 12572 6854
rect 12728 6390 12756 7142
rect 12820 7002 12848 7296
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12452 6066 12480 6190
rect 12360 6038 12480 6066
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12360 5370 12388 6038
rect 12728 5914 12756 6054
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12452 5030 12480 5714
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12346 4856 12402 4865
rect 12346 4791 12402 4800
rect 12360 3924 12388 4791
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12452 4078 12480 4694
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12440 3936 12492 3942
rect 12360 3896 12440 3924
rect 12440 3878 12492 3884
rect 12268 3590 12480 3618
rect 12256 3460 12308 3466
rect 12256 3402 12308 3408
rect 12268 2650 12296 3402
rect 12452 3380 12480 3590
rect 12360 3352 12480 3380
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 12360 2496 12388 3352
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 2650 12480 2790
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12440 2508 12492 2514
rect 12360 2468 12440 2496
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12176 1630 12204 2246
rect 12268 2038 12296 2246
rect 12256 2032 12308 2038
rect 12256 1974 12308 1980
rect 12164 1624 12216 1630
rect 12164 1566 12216 1572
rect 12360 480 12388 2468
rect 12440 2450 12492 2456
rect 12438 2408 12494 2417
rect 12438 2343 12440 2352
rect 12492 2343 12494 2352
rect 12440 2314 12492 2320
rect 12544 2038 12572 5850
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12636 3505 12664 5238
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 12622 3496 12678 3505
rect 12622 3431 12678 3440
rect 12622 3360 12678 3369
rect 12622 3295 12678 3304
rect 12532 2032 12584 2038
rect 12532 1974 12584 1980
rect 12636 480 12664 3295
rect 12728 2582 12756 4694
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 12820 2378 12848 6734
rect 12912 6089 12940 7142
rect 12898 6080 12954 6089
rect 12898 6015 12954 6024
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12912 3097 12940 5850
rect 13004 5710 13032 7346
rect 13096 6361 13124 8026
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13082 6352 13138 6361
rect 13082 6287 13138 6296
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 13004 5234 13032 5646
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 12992 4548 13044 4554
rect 12992 4490 13044 4496
rect 13004 4146 13032 4490
rect 13096 4146 13124 6190
rect 13188 4826 13216 7890
rect 13464 7818 13492 8026
rect 13556 7818 13584 8327
rect 13728 8298 13780 8304
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13282 7644 13578 7664
rect 13338 7642 13362 7644
rect 13418 7642 13442 7644
rect 13498 7642 13522 7644
rect 13360 7590 13362 7642
rect 13424 7590 13436 7642
rect 13498 7590 13500 7642
rect 13338 7588 13362 7590
rect 13418 7588 13442 7590
rect 13498 7588 13522 7590
rect 13282 7568 13578 7588
rect 13648 7449 13676 7686
rect 13634 7440 13690 7449
rect 13634 7375 13690 7384
rect 13634 7304 13690 7313
rect 13634 7239 13690 7248
rect 13648 7206 13676 7239
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13740 7018 13768 8298
rect 13648 6990 13768 7018
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13648 6338 13676 6990
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13556 6310 13676 6338
rect 13360 6180 13412 6186
rect 13360 6122 13412 6128
rect 13372 5710 13400 6122
rect 13556 5930 13584 6310
rect 13634 6216 13690 6225
rect 13634 6151 13690 6160
rect 13648 6118 13676 6151
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13556 5902 13676 5930
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13648 5370 13676 5902
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13450 5264 13506 5273
rect 13450 5199 13452 5208
rect 13504 5199 13506 5208
rect 13452 5170 13504 5176
rect 13634 5128 13690 5137
rect 13268 5092 13320 5098
rect 13634 5063 13636 5072
rect 13268 5034 13320 5040
rect 13688 5063 13690 5072
rect 13636 5034 13688 5040
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13280 4706 13308 5034
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13188 4678 13308 4706
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13096 3194 13124 4082
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 12898 3088 12954 3097
rect 12898 3023 12954 3032
rect 12992 2916 13044 2922
rect 12992 2858 13044 2864
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 12912 2553 12940 2790
rect 13004 2582 13032 2858
rect 12992 2576 13044 2582
rect 12898 2544 12954 2553
rect 12992 2518 13044 2524
rect 12898 2479 12954 2488
rect 13188 2428 13216 4678
rect 13282 4380 13578 4400
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 13648 4282 13676 4762
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13266 4176 13322 4185
rect 13266 4111 13322 4120
rect 13280 4078 13308 4111
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13634 3904 13690 3913
rect 13280 3738 13308 3878
rect 13634 3839 13690 3848
rect 13648 3738 13676 3839
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13266 3496 13322 3505
rect 13266 3431 13268 3440
rect 13320 3431 13322 3440
rect 13268 3402 13320 3408
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 13740 3194 13768 6870
rect 13832 6769 13860 8774
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13818 6760 13874 6769
rect 13818 6695 13874 6704
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5166 13860 6054
rect 13924 5778 13952 8366
rect 14016 7478 14044 9658
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 14108 6882 14136 12038
rect 14200 10470 14228 13806
rect 14292 12646 14320 15558
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 9722 14228 10406
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14200 9081 14228 9318
rect 14186 9072 14242 9081
rect 14186 9007 14242 9016
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14200 7886 14228 8434
rect 14292 8401 14320 12582
rect 14384 11257 14412 14758
rect 14476 13870 14504 18022
rect 14554 16144 14610 16153
rect 14554 16079 14610 16088
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14370 11248 14426 11257
rect 14370 11183 14426 11192
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 14278 8392 14334 8401
rect 14278 8327 14334 8336
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14016 6854 14136 6882
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13832 3670 13860 4966
rect 13924 3738 13952 5510
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13832 3058 13860 3402
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13636 2848 13688 2854
rect 13634 2816 13636 2825
rect 13688 2816 13690 2825
rect 13634 2751 13690 2760
rect 13004 2400 13216 2428
rect 12808 2372 12860 2378
rect 12808 2314 12860 2320
rect 13004 480 13032 2400
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 13360 2032 13412 2038
rect 13360 1974 13412 1980
rect 13372 480 13400 1974
rect 13648 1902 13676 2751
rect 13924 2446 13952 2926
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 13728 2372 13780 2378
rect 13728 2314 13780 2320
rect 13636 1896 13688 1902
rect 13636 1838 13688 1844
rect 13740 480 13768 2314
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 13912 2304 13964 2310
rect 13912 2246 13964 2252
rect 13832 1766 13860 2246
rect 13924 2106 13952 2246
rect 13912 2100 13964 2106
rect 13912 2042 13964 2048
rect 13820 1760 13872 1766
rect 13820 1702 13872 1708
rect 14016 480 14044 6854
rect 14292 6440 14320 8230
rect 14108 6412 14320 6440
rect 14108 4865 14136 6412
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14200 5642 14228 6054
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14094 4856 14150 4865
rect 14094 4791 14150 4800
rect 14200 4622 14228 5170
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14094 3904 14150 3913
rect 14094 3839 14150 3848
rect 14108 3602 14136 3839
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14094 3496 14150 3505
rect 14094 3431 14150 3440
rect 14108 3058 14136 3431
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14094 2952 14150 2961
rect 14094 2887 14150 2896
rect 14108 2854 14136 2887
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 14200 2650 14228 3606
rect 14292 3058 14320 6258
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14384 2938 14412 11018
rect 14476 9042 14504 13262
rect 14568 10130 14596 16079
rect 14752 12866 14780 19520
rect 15028 18170 15056 19520
rect 15028 18142 15332 18170
rect 15304 17898 15332 18142
rect 15212 17870 15332 17898
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 14660 12838 14780 12866
rect 14830 12880 14886 12889
rect 14660 10130 14688 12838
rect 14830 12815 14886 12824
rect 14844 12782 14872 12815
rect 14832 12776 14884 12782
rect 14738 12744 14794 12753
rect 14832 12718 14884 12724
rect 14738 12679 14794 12688
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14462 8936 14518 8945
rect 14462 8871 14518 8880
rect 14476 6866 14504 8871
rect 14568 8430 14596 10066
rect 14646 10024 14702 10033
rect 14646 9959 14648 9968
rect 14700 9959 14702 9968
rect 14648 9930 14700 9936
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14752 7698 14780 12679
rect 14936 11676 14964 13942
rect 15028 12753 15056 14214
rect 15014 12744 15070 12753
rect 15014 12679 15070 12688
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 14568 7670 14780 7698
rect 14844 11648 14964 11676
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14476 4214 14504 5646
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14476 3097 14504 3878
rect 14462 3088 14518 3097
rect 14462 3023 14518 3032
rect 14292 2910 14412 2938
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14292 2378 14320 2910
rect 14568 2836 14596 7670
rect 14844 7290 14872 11648
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14936 9178 14964 10066
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14936 8430 14964 9114
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14924 7812 14976 7818
rect 14924 7754 14976 7760
rect 14936 7342 14964 7754
rect 14752 7262 14872 7290
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14660 5030 14688 6802
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14646 4584 14702 4593
rect 14646 4519 14648 4528
rect 14700 4519 14702 4528
rect 14648 4490 14700 4496
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14660 3777 14688 3878
rect 14646 3768 14702 3777
rect 14646 3703 14702 3712
rect 14384 2808 14596 2836
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 14384 480 14412 2808
rect 14752 480 14780 7262
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 14844 1834 14872 7142
rect 14936 5953 14964 7142
rect 14922 5944 14978 5953
rect 14922 5879 14978 5888
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 14936 4185 14964 5102
rect 14922 4176 14978 4185
rect 14922 4111 14978 4120
rect 14832 1828 14884 1834
rect 14832 1770 14884 1776
rect 15028 480 15056 12582
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15120 10033 15148 11698
rect 15212 10810 15240 17870
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15212 10713 15240 10746
rect 15198 10704 15254 10713
rect 15198 10639 15254 10648
rect 15304 10588 15332 13670
rect 15396 13326 15424 19520
rect 15764 13734 15792 19520
rect 16040 18086 16068 19520
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16408 16153 16436 19520
rect 16394 16144 16450 16153
rect 16394 16079 16450 16088
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15212 10560 15332 10588
rect 15106 10024 15162 10033
rect 15106 9959 15162 9968
rect 15212 7188 15240 10560
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15120 7160 15240 7188
rect 15120 6186 15148 7160
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15120 2922 15148 5714
rect 15198 4992 15254 5001
rect 15198 4927 15254 4936
rect 15212 4078 15240 4927
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 15304 2514 15332 9862
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15396 480 15424 12174
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15488 6254 15516 9998
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15580 3369 15608 10134
rect 15566 3360 15622 3369
rect 15566 3295 15622 3304
rect 15764 480 15792 12650
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16028 1964 16080 1970
rect 16028 1906 16080 1912
rect 16040 480 16068 1906
rect 16408 480 16436 11562
rect 16776 10606 16804 19520
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16762 4040 16818 4049
rect 16762 3975 16818 3984
rect 16776 480 16804 3975
rect 2870 439 2926 448
rect 3146 0 3202 480
rect 3514 0 3570 480
rect 3790 0 3846 480
rect 4158 0 4214 480
rect 4526 0 4582 480
rect 4802 0 4858 480
rect 5170 0 5226 480
rect 5538 0 5594 480
rect 5814 0 5870 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7194 0 7250 480
rect 7562 0 7618 480
rect 7930 0 7986 480
rect 8206 0 8262 480
rect 8574 0 8630 480
rect 8942 0 8998 480
rect 9218 0 9274 480
rect 9586 0 9642 480
rect 9954 0 10010 480
rect 10322 0 10378 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11610 0 11666 480
rect 11978 0 12034 480
rect 12346 0 12402 480
rect 12622 0 12678 480
rect 12990 0 13046 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14002 0 14058 480
rect 14370 0 14426 480
rect 14738 0 14794 480
rect 15014 0 15070 480
rect 15382 0 15438 480
rect 15750 0 15806 480
rect 16026 0 16082 480
rect 16394 0 16450 480
rect 16762 0 16818 480
<< via2 >>
rect 1490 19352 1546 19408
rect 1674 18400 1730 18456
rect 1306 15000 1362 15056
rect 1398 12824 1454 12880
rect 1214 8356 1270 8392
rect 1214 8336 1216 8356
rect 1216 8336 1268 8356
rect 1268 8336 1270 8356
rect 1214 8200 1270 8256
rect 1582 8064 1638 8120
rect 1950 11212 2006 11248
rect 1950 11192 1952 11212
rect 1952 11192 2004 11212
rect 2004 11192 2006 11212
rect 1858 10376 1914 10432
rect 1766 8064 1822 8120
rect 1582 7928 1638 7984
rect 1766 7928 1822 7984
rect 1122 2896 1178 2952
rect 1858 7248 1914 7304
rect 1858 4684 1914 4720
rect 1858 4664 1860 4684
rect 1860 4664 1912 4684
rect 1912 4664 1914 4684
rect 1766 3576 1822 3632
rect 1490 3168 1546 3224
rect 2226 13268 2228 13288
rect 2228 13268 2280 13288
rect 2280 13268 2282 13288
rect 2226 13232 2282 13268
rect 2226 12144 2282 12200
rect 2410 14456 2466 14512
rect 3054 17312 3110 17368
rect 2778 16360 2834 16416
rect 2686 15544 2742 15600
rect 2594 12688 2650 12744
rect 3421 17434 3477 17436
rect 3501 17434 3557 17436
rect 3581 17434 3637 17436
rect 3661 17434 3717 17436
rect 3421 17382 3447 17434
rect 3447 17382 3477 17434
rect 3501 17382 3511 17434
rect 3511 17382 3557 17434
rect 3581 17382 3627 17434
rect 3627 17382 3637 17434
rect 3661 17382 3691 17434
rect 3691 17382 3717 17434
rect 3421 17380 3477 17382
rect 3501 17380 3557 17382
rect 3581 17380 3637 17382
rect 3661 17380 3717 17382
rect 3330 16768 3386 16824
rect 2962 12416 3018 12472
rect 2502 9444 2558 9480
rect 2502 9424 2504 9444
rect 2504 9424 2556 9444
rect 2556 9424 2558 9444
rect 2870 9968 2926 10024
rect 3146 13776 3202 13832
rect 3421 16346 3477 16348
rect 3501 16346 3557 16348
rect 3581 16346 3637 16348
rect 3661 16346 3717 16348
rect 3421 16294 3447 16346
rect 3447 16294 3477 16346
rect 3501 16294 3511 16346
rect 3511 16294 3557 16346
rect 3581 16294 3627 16346
rect 3627 16294 3637 16346
rect 3661 16294 3691 16346
rect 3691 16294 3717 16346
rect 3421 16292 3477 16294
rect 3501 16292 3557 16294
rect 3581 16292 3637 16294
rect 3661 16292 3717 16294
rect 3606 15408 3662 15464
rect 3421 15258 3477 15260
rect 3501 15258 3557 15260
rect 3581 15258 3637 15260
rect 3661 15258 3717 15260
rect 3421 15206 3447 15258
rect 3447 15206 3477 15258
rect 3501 15206 3511 15258
rect 3511 15206 3557 15258
rect 3581 15206 3627 15258
rect 3627 15206 3637 15258
rect 3661 15206 3691 15258
rect 3691 15206 3717 15258
rect 3421 15204 3477 15206
rect 3501 15204 3557 15206
rect 3581 15204 3637 15206
rect 3661 15204 3717 15206
rect 3421 14170 3477 14172
rect 3501 14170 3557 14172
rect 3581 14170 3637 14172
rect 3661 14170 3717 14172
rect 3421 14118 3447 14170
rect 3447 14118 3477 14170
rect 3501 14118 3511 14170
rect 3511 14118 3557 14170
rect 3581 14118 3627 14170
rect 3627 14118 3637 14170
rect 3661 14118 3691 14170
rect 3691 14118 3717 14170
rect 3421 14116 3477 14118
rect 3501 14116 3557 14118
rect 3581 14116 3637 14118
rect 3661 14116 3717 14118
rect 3054 11328 3110 11384
rect 2134 7792 2190 7848
rect 2502 7520 2558 7576
rect 2686 8064 2742 8120
rect 2594 6160 2650 6216
rect 2134 4528 2190 4584
rect 2042 1400 2098 1456
rect 2778 7656 2834 7712
rect 2502 3984 2558 4040
rect 2594 3440 2650 3496
rect 2962 9152 3018 9208
rect 2962 7656 3018 7712
rect 2870 6840 2926 6896
rect 3054 7384 3110 7440
rect 3421 13082 3477 13084
rect 3501 13082 3557 13084
rect 3581 13082 3637 13084
rect 3661 13082 3717 13084
rect 3421 13030 3447 13082
rect 3447 13030 3477 13082
rect 3501 13030 3511 13082
rect 3511 13030 3557 13082
rect 3581 13030 3627 13082
rect 3627 13030 3637 13082
rect 3661 13030 3691 13082
rect 3691 13030 3717 13082
rect 3421 13028 3477 13030
rect 3501 13028 3557 13030
rect 3581 13028 3637 13030
rect 3661 13028 3717 13030
rect 3421 11994 3477 11996
rect 3501 11994 3557 11996
rect 3581 11994 3637 11996
rect 3661 11994 3717 11996
rect 3421 11942 3447 11994
rect 3447 11942 3477 11994
rect 3501 11942 3511 11994
rect 3511 11942 3557 11994
rect 3581 11942 3627 11994
rect 3627 11942 3637 11994
rect 3661 11942 3691 11994
rect 3691 11942 3717 11994
rect 3421 11940 3477 11942
rect 3501 11940 3557 11942
rect 3581 11940 3637 11942
rect 3661 11940 3717 11942
rect 3421 10906 3477 10908
rect 3501 10906 3557 10908
rect 3581 10906 3637 10908
rect 3661 10906 3717 10908
rect 3421 10854 3447 10906
rect 3447 10854 3477 10906
rect 3501 10854 3511 10906
rect 3511 10854 3557 10906
rect 3581 10854 3627 10906
rect 3627 10854 3637 10906
rect 3661 10854 3691 10906
rect 3691 10854 3717 10906
rect 3421 10852 3477 10854
rect 3501 10852 3557 10854
rect 3581 10852 3637 10854
rect 3661 10852 3717 10854
rect 4158 16360 4214 16416
rect 3421 9818 3477 9820
rect 3501 9818 3557 9820
rect 3581 9818 3637 9820
rect 3661 9818 3717 9820
rect 3421 9766 3447 9818
rect 3447 9766 3477 9818
rect 3501 9766 3511 9818
rect 3511 9766 3557 9818
rect 3581 9766 3627 9818
rect 3627 9766 3637 9818
rect 3661 9766 3691 9818
rect 3691 9766 3717 9818
rect 3421 9764 3477 9766
rect 3501 9764 3557 9766
rect 3581 9764 3637 9766
rect 3661 9764 3717 9766
rect 3421 8730 3477 8732
rect 3501 8730 3557 8732
rect 3581 8730 3637 8732
rect 3661 8730 3717 8732
rect 3421 8678 3447 8730
rect 3447 8678 3477 8730
rect 3501 8678 3511 8730
rect 3511 8678 3557 8730
rect 3581 8678 3627 8730
rect 3627 8678 3637 8730
rect 3661 8678 3691 8730
rect 3691 8678 3717 8730
rect 3421 8676 3477 8678
rect 3501 8676 3557 8678
rect 3581 8676 3637 8678
rect 3661 8676 3717 8678
rect 3606 8336 3662 8392
rect 2962 5344 3018 5400
rect 2962 4392 3018 4448
rect 3514 7928 3570 7984
rect 3422 7792 3478 7848
rect 3698 7792 3754 7848
rect 3421 7642 3477 7644
rect 3501 7642 3557 7644
rect 3581 7642 3637 7644
rect 3661 7642 3717 7644
rect 3421 7590 3447 7642
rect 3447 7590 3477 7642
rect 3501 7590 3511 7642
rect 3511 7590 3557 7642
rect 3581 7590 3627 7642
rect 3627 7590 3637 7642
rect 3661 7590 3691 7642
rect 3691 7590 3717 7642
rect 3421 7588 3477 7590
rect 3501 7588 3557 7590
rect 3581 7588 3637 7590
rect 3661 7588 3717 7590
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 3422 5092 3478 5128
rect 3422 5072 3424 5092
rect 3424 5072 3476 5092
rect 3476 5072 3478 5092
rect 4250 14320 4306 14376
rect 4250 13776 4306 13832
rect 4710 16244 4766 16280
rect 4986 17196 5042 17232
rect 4986 17176 4988 17196
rect 4988 17176 5040 17196
rect 5040 17176 5042 17196
rect 5354 16652 5410 16688
rect 5354 16632 5356 16652
rect 5356 16632 5408 16652
rect 5408 16632 5410 16652
rect 4710 16224 4712 16244
rect 4712 16224 4764 16244
rect 4764 16224 4766 16244
rect 4894 16088 4950 16144
rect 4894 14320 4950 14376
rect 4526 12960 4582 13016
rect 4710 12300 4766 12336
rect 4710 12280 4712 12300
rect 4712 12280 4764 12300
rect 4764 12280 4766 12300
rect 4342 11872 4398 11928
rect 4342 11600 4398 11656
rect 3882 8472 3938 8528
rect 4618 12144 4674 12200
rect 4526 8916 4528 8936
rect 4528 8916 4580 8936
rect 4580 8916 4582 8936
rect 4526 8880 4582 8916
rect 4158 8336 4214 8392
rect 3882 5480 3938 5536
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 2778 3032 2834 3088
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 3054 2488 3110 2544
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 2870 448 2926 504
rect 4342 8608 4398 8664
rect 4434 8084 4490 8120
rect 4434 8064 4436 8084
rect 4436 8064 4488 8084
rect 4488 8064 4490 8084
rect 4250 7792 4306 7848
rect 4618 7656 4674 7712
rect 4618 7520 4674 7576
rect 4434 6840 4490 6896
rect 4250 5072 4306 5128
rect 4342 4256 4398 4312
rect 4526 5752 4582 5808
rect 4894 11636 4896 11656
rect 4896 11636 4948 11656
rect 4948 11636 4950 11656
rect 4894 11600 4950 11636
rect 4802 9968 4858 10024
rect 5886 16890 5942 16892
rect 5966 16890 6022 16892
rect 6046 16890 6102 16892
rect 6126 16890 6182 16892
rect 5886 16838 5912 16890
rect 5912 16838 5942 16890
rect 5966 16838 5976 16890
rect 5976 16838 6022 16890
rect 6046 16838 6092 16890
rect 6092 16838 6102 16890
rect 6126 16838 6156 16890
rect 6156 16838 6182 16890
rect 5886 16836 5942 16838
rect 5966 16836 6022 16838
rect 6046 16836 6102 16838
rect 6126 16836 6182 16838
rect 5814 16496 5870 16552
rect 5170 12960 5226 13016
rect 5722 15444 5724 15464
rect 5724 15444 5776 15464
rect 5776 15444 5778 15464
rect 5722 15408 5778 15444
rect 5630 13776 5686 13832
rect 5886 15802 5942 15804
rect 5966 15802 6022 15804
rect 6046 15802 6102 15804
rect 6126 15802 6182 15804
rect 5886 15750 5912 15802
rect 5912 15750 5942 15802
rect 5966 15750 5976 15802
rect 5976 15750 6022 15802
rect 6046 15750 6092 15802
rect 6092 15750 6102 15802
rect 6126 15750 6156 15802
rect 6156 15750 6182 15802
rect 5886 15748 5942 15750
rect 5966 15748 6022 15750
rect 6046 15748 6102 15750
rect 6126 15748 6182 15750
rect 7010 16224 7066 16280
rect 6826 16124 6828 16144
rect 6828 16124 6880 16144
rect 6880 16124 6882 16144
rect 6550 15952 6606 16008
rect 6366 14864 6422 14920
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 6126 14714 6182 14716
rect 5886 14662 5912 14714
rect 5912 14662 5942 14714
rect 5966 14662 5976 14714
rect 5976 14662 6022 14714
rect 6046 14662 6092 14714
rect 6092 14662 6102 14714
rect 6126 14662 6156 14714
rect 6156 14662 6182 14714
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 6126 14660 6182 14662
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 6126 13626 6182 13628
rect 5886 13574 5912 13626
rect 5912 13574 5942 13626
rect 5966 13574 5976 13626
rect 5976 13574 6022 13626
rect 6046 13574 6092 13626
rect 6092 13574 6102 13626
rect 6126 13574 6156 13626
rect 6156 13574 6182 13626
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 6126 13572 6182 13574
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 6126 12538 6182 12540
rect 5886 12486 5912 12538
rect 5912 12486 5942 12538
rect 5966 12486 5976 12538
rect 5976 12486 6022 12538
rect 6046 12486 6092 12538
rect 6092 12486 6102 12538
rect 6126 12486 6156 12538
rect 6156 12486 6182 12538
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 6126 12484 6182 12486
rect 6826 16088 6882 16124
rect 6642 14728 6698 14784
rect 6918 15408 6974 15464
rect 7194 16088 7250 16144
rect 7194 15000 7250 15056
rect 7102 13504 7158 13560
rect 6550 12688 6606 12744
rect 5538 11872 5594 11928
rect 6918 13232 6974 13288
rect 7102 12416 7158 12472
rect 5078 9868 5080 9888
rect 5080 9868 5132 9888
rect 5132 9868 5134 9888
rect 5078 9832 5134 9868
rect 6366 11736 6422 11792
rect 5814 11600 5870 11656
rect 6274 11464 6330 11520
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 6126 11450 6182 11452
rect 5886 11398 5912 11450
rect 5912 11398 5942 11450
rect 5966 11398 5976 11450
rect 5976 11398 6022 11450
rect 6046 11398 6092 11450
rect 6092 11398 6102 11450
rect 6126 11398 6156 11450
rect 6156 11398 6182 11450
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 6126 11396 6182 11398
rect 5814 11076 5870 11112
rect 5814 11056 5816 11076
rect 5816 11056 5868 11076
rect 5868 11056 5870 11076
rect 4986 8916 4988 8936
rect 4988 8916 5040 8936
rect 5040 8916 5042 8936
rect 4986 8880 5042 8916
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 6126 10362 6182 10364
rect 5886 10310 5912 10362
rect 5912 10310 5942 10362
rect 5966 10310 5976 10362
rect 5976 10310 6022 10362
rect 6046 10310 6092 10362
rect 6092 10310 6102 10362
rect 6126 10310 6156 10362
rect 6156 10310 6182 10362
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 6126 10308 6182 10310
rect 5538 9832 5594 9888
rect 5630 9152 5686 9208
rect 5722 9016 5778 9072
rect 4434 3168 4490 3224
rect 4158 1944 4214 2000
rect 4618 4392 4674 4448
rect 5262 6296 5318 6352
rect 5078 5480 5134 5536
rect 4986 4256 5042 4312
rect 5078 4120 5134 4176
rect 4618 2760 4674 2816
rect 4986 2760 5042 2816
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 6126 9274 6182 9276
rect 5886 9222 5912 9274
rect 5912 9222 5942 9274
rect 5966 9222 5976 9274
rect 5976 9222 6022 9274
rect 6046 9222 6092 9274
rect 6092 9222 6102 9274
rect 6126 9222 6156 9274
rect 6156 9222 6182 9274
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 6126 9220 6182 9222
rect 5814 8608 5870 8664
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 6126 8186 6182 8188
rect 5886 8134 5912 8186
rect 5912 8134 5942 8186
rect 5966 8134 5976 8186
rect 5976 8134 6022 8186
rect 6046 8134 6092 8186
rect 6092 8134 6102 8186
rect 6126 8134 6156 8186
rect 6156 8134 6182 8186
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 6126 8132 6182 8134
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 6126 7098 6182 7100
rect 5886 7046 5912 7098
rect 5912 7046 5942 7098
rect 5966 7046 5976 7098
rect 5976 7046 6022 7098
rect 6046 7046 6092 7098
rect 6092 7046 6102 7098
rect 6126 7046 6156 7098
rect 6156 7046 6182 7098
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 6126 7044 6182 7046
rect 6274 6704 6330 6760
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 5354 4256 5410 4312
rect 5630 3168 5686 3224
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 7010 11328 7066 11384
rect 6642 10648 6698 10704
rect 6550 9968 6606 10024
rect 7286 13232 7342 13288
rect 7746 16940 7748 16960
rect 7748 16940 7800 16960
rect 7800 16940 7802 16960
rect 7746 16904 7802 16940
rect 7746 16768 7802 16824
rect 7562 16224 7618 16280
rect 7746 16088 7802 16144
rect 7654 15408 7710 15464
rect 8114 16788 8170 16824
rect 8114 16768 8116 16788
rect 8116 16768 8168 16788
rect 8168 16768 8170 16788
rect 8850 17892 8852 17912
rect 8852 17892 8904 17912
rect 8904 17892 8906 17912
rect 8850 17856 8906 17892
rect 8352 17434 8408 17436
rect 8432 17434 8488 17436
rect 8512 17434 8568 17436
rect 8592 17434 8648 17436
rect 8352 17382 8378 17434
rect 8378 17382 8408 17434
rect 8432 17382 8442 17434
rect 8442 17382 8488 17434
rect 8512 17382 8558 17434
rect 8558 17382 8568 17434
rect 8592 17382 8622 17434
rect 8622 17382 8648 17434
rect 8352 17380 8408 17382
rect 8432 17380 8488 17382
rect 8512 17380 8568 17382
rect 8592 17380 8648 17382
rect 8482 17060 8538 17096
rect 8482 17040 8484 17060
rect 8484 17040 8536 17060
rect 8536 17040 8538 17060
rect 8298 16788 8354 16824
rect 8298 16768 8300 16788
rect 8300 16768 8352 16788
rect 8352 16768 8354 16788
rect 8758 17584 8814 17640
rect 8206 16360 8262 16416
rect 8352 16346 8408 16348
rect 8432 16346 8488 16348
rect 8512 16346 8568 16348
rect 8592 16346 8648 16348
rect 8352 16294 8378 16346
rect 8378 16294 8408 16346
rect 8432 16294 8442 16346
rect 8442 16294 8488 16346
rect 8512 16294 8558 16346
rect 8558 16294 8568 16346
rect 8592 16294 8622 16346
rect 8622 16294 8648 16346
rect 8352 16292 8408 16294
rect 8432 16292 8488 16294
rect 8512 16292 8568 16294
rect 8592 16292 8648 16294
rect 8114 15700 8170 15736
rect 8114 15680 8116 15700
rect 8116 15680 8168 15700
rect 8168 15680 8170 15700
rect 7562 14728 7618 14784
rect 7930 15000 7986 15056
rect 8352 15258 8408 15260
rect 8432 15258 8488 15260
rect 8512 15258 8568 15260
rect 8592 15258 8648 15260
rect 8352 15206 8378 15258
rect 8378 15206 8408 15258
rect 8432 15206 8442 15258
rect 8442 15206 8488 15258
rect 8512 15206 8558 15258
rect 8558 15206 8568 15258
rect 8592 15206 8622 15258
rect 8622 15206 8648 15258
rect 8352 15204 8408 15206
rect 8432 15204 8488 15206
rect 8512 15204 8568 15206
rect 8592 15204 8648 15206
rect 8390 14884 8446 14920
rect 8390 14864 8392 14884
rect 8392 14864 8444 14884
rect 8444 14864 8446 14884
rect 8666 14456 8722 14512
rect 8352 14170 8408 14172
rect 8432 14170 8488 14172
rect 8512 14170 8568 14172
rect 8592 14170 8648 14172
rect 8352 14118 8378 14170
rect 8378 14118 8408 14170
rect 8432 14118 8442 14170
rect 8442 14118 8488 14170
rect 8512 14118 8558 14170
rect 8558 14118 8568 14170
rect 8592 14118 8622 14170
rect 8622 14118 8648 14170
rect 8352 14116 8408 14118
rect 8432 14116 8488 14118
rect 8512 14116 8568 14118
rect 8592 14116 8648 14118
rect 8206 13640 8262 13696
rect 7470 10376 7526 10432
rect 7102 9288 7158 9344
rect 7654 9868 7656 9888
rect 7656 9868 7708 9888
rect 7708 9868 7710 9888
rect 7654 9832 7710 9868
rect 7654 9560 7710 9616
rect 7562 9152 7618 9208
rect 7194 8880 7250 8936
rect 7470 8900 7526 8936
rect 7930 12300 7986 12336
rect 7930 12280 7932 12300
rect 7932 12280 7984 12300
rect 7984 12280 7986 12300
rect 7930 12144 7986 12200
rect 8352 13082 8408 13084
rect 8432 13082 8488 13084
rect 8512 13082 8568 13084
rect 8592 13082 8648 13084
rect 8352 13030 8378 13082
rect 8378 13030 8408 13082
rect 8432 13030 8442 13082
rect 8442 13030 8488 13082
rect 8512 13030 8558 13082
rect 8558 13030 8568 13082
rect 8592 13030 8622 13082
rect 8622 13030 8648 13082
rect 8352 13028 8408 13030
rect 8432 13028 8488 13030
rect 8512 13028 8568 13030
rect 8592 13028 8648 13030
rect 8942 14184 8998 14240
rect 8206 12008 8262 12064
rect 8352 11994 8408 11996
rect 8432 11994 8488 11996
rect 8512 11994 8568 11996
rect 8592 11994 8648 11996
rect 8352 11942 8378 11994
rect 8378 11942 8408 11994
rect 8432 11942 8442 11994
rect 8442 11942 8488 11994
rect 8512 11942 8558 11994
rect 8558 11942 8568 11994
rect 8592 11942 8622 11994
rect 8622 11942 8648 11994
rect 8352 11940 8408 11942
rect 8432 11940 8488 11942
rect 8512 11940 8568 11942
rect 8592 11940 8648 11942
rect 8206 11872 8262 11928
rect 8482 11600 8538 11656
rect 8666 11600 8722 11656
rect 8666 11056 8722 11112
rect 8352 10906 8408 10908
rect 8432 10906 8488 10908
rect 8512 10906 8568 10908
rect 8592 10906 8648 10908
rect 8352 10854 8378 10906
rect 8378 10854 8408 10906
rect 8432 10854 8442 10906
rect 8442 10854 8488 10906
rect 8512 10854 8558 10906
rect 8558 10854 8568 10906
rect 8592 10854 8622 10906
rect 8622 10854 8648 10906
rect 8352 10852 8408 10854
rect 8432 10852 8488 10854
rect 8512 10852 8568 10854
rect 8592 10852 8648 10854
rect 8206 10376 8262 10432
rect 8206 10240 8262 10296
rect 7470 8880 7472 8900
rect 7472 8880 7524 8900
rect 7524 8880 7526 8900
rect 7470 8064 7526 8120
rect 7838 7656 7894 7712
rect 7010 6996 7066 7032
rect 7010 6976 7012 6996
rect 7012 6976 7064 6996
rect 7064 6976 7066 6996
rect 7838 7112 7894 7168
rect 7838 6704 7894 6760
rect 6642 4800 6698 4856
rect 6826 4800 6882 4856
rect 6918 4664 6974 4720
rect 7010 2760 7066 2816
rect 7470 4428 7472 4448
rect 7472 4428 7524 4448
rect 7524 4428 7526 4448
rect 7470 4392 7526 4428
rect 7838 5480 7894 5536
rect 7746 5344 7802 5400
rect 7746 4256 7802 4312
rect 7562 4120 7618 4176
rect 7562 3712 7618 3768
rect 7562 2488 7618 2544
rect 8022 9560 8078 9616
rect 8352 9818 8408 9820
rect 8432 9818 8488 9820
rect 8512 9818 8568 9820
rect 8592 9818 8648 9820
rect 8352 9766 8378 9818
rect 8378 9766 8408 9818
rect 8432 9766 8442 9818
rect 8442 9766 8488 9818
rect 8512 9766 8558 9818
rect 8558 9766 8568 9818
rect 8592 9766 8622 9818
rect 8622 9766 8648 9818
rect 8352 9764 8408 9766
rect 8432 9764 8488 9766
rect 8512 9764 8568 9766
rect 8592 9764 8648 9766
rect 8114 9288 8170 9344
rect 8390 9288 8446 9344
rect 8666 9152 8722 9208
rect 8352 8730 8408 8732
rect 8432 8730 8488 8732
rect 8512 8730 8568 8732
rect 8592 8730 8648 8732
rect 8352 8678 8378 8730
rect 8378 8678 8408 8730
rect 8432 8678 8442 8730
rect 8442 8678 8488 8730
rect 8512 8678 8558 8730
rect 8558 8678 8568 8730
rect 8592 8678 8622 8730
rect 8622 8678 8648 8730
rect 8352 8676 8408 8678
rect 8432 8676 8488 8678
rect 8512 8676 8568 8678
rect 8592 8676 8648 8678
rect 8206 7792 8262 7848
rect 8352 7642 8408 7644
rect 8432 7642 8488 7644
rect 8512 7642 8568 7644
rect 8592 7642 8648 7644
rect 8352 7590 8378 7642
rect 8378 7590 8408 7642
rect 8432 7590 8442 7642
rect 8442 7590 8488 7642
rect 8512 7590 8558 7642
rect 8558 7590 8568 7642
rect 8592 7590 8622 7642
rect 8622 7590 8648 7642
rect 8352 7588 8408 7590
rect 8432 7588 8488 7590
rect 8512 7588 8568 7590
rect 8592 7588 8648 7590
rect 8206 7520 8262 7576
rect 8482 6976 8538 7032
rect 8666 6840 8722 6896
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 8206 6060 8208 6080
rect 8208 6060 8260 6080
rect 8260 6060 8262 6080
rect 8206 6024 8262 6060
rect 8022 4664 8078 4720
rect 7930 3848 7986 3904
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 8482 4800 8538 4856
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 8206 3168 8262 3224
rect 8574 2488 8630 2544
rect 8666 2352 8722 2408
rect 8850 12436 8906 12472
rect 8850 12416 8852 12436
rect 8852 12416 8904 12436
rect 8904 12416 8906 12436
rect 8850 12008 8906 12064
rect 9402 16360 9458 16416
rect 9310 15680 9366 15736
rect 9586 16768 9642 16824
rect 9494 16224 9550 16280
rect 9494 15272 9550 15328
rect 9402 13776 9458 13832
rect 9310 13640 9366 13696
rect 9218 13096 9274 13152
rect 9586 14728 9642 14784
rect 9586 14048 9642 14104
rect 9862 16244 9918 16280
rect 9862 16224 9864 16244
rect 9864 16224 9916 16244
rect 9916 16224 9918 16244
rect 9770 15408 9826 15464
rect 9954 14884 10010 14920
rect 9954 14864 9956 14884
rect 9956 14864 10008 14884
rect 10008 14864 10010 14884
rect 9770 14592 9826 14648
rect 10138 16768 10194 16824
rect 10138 15680 10194 15736
rect 10138 14764 10140 14784
rect 10140 14764 10192 14784
rect 10192 14764 10194 14784
rect 10138 14728 10194 14764
rect 9770 14048 9826 14104
rect 9678 13232 9734 13288
rect 9862 13232 9918 13288
rect 9862 12688 9918 12744
rect 9310 12552 9366 12608
rect 9310 12436 9366 12472
rect 9310 12416 9312 12436
rect 9312 12416 9364 12436
rect 9364 12416 9366 12436
rect 8942 11056 8998 11112
rect 9034 10920 9090 10976
rect 8942 8084 8998 8120
rect 8942 8064 8944 8084
rect 8944 8064 8996 8084
rect 8996 8064 8998 8084
rect 9586 11464 9642 11520
rect 9402 10512 9458 10568
rect 9218 8200 9274 8256
rect 9126 7112 9182 7168
rect 9034 5344 9090 5400
rect 9218 6024 9274 6080
rect 9586 10512 9642 10568
rect 10138 13404 10140 13424
rect 10140 13404 10192 13424
rect 10192 13404 10194 13424
rect 10138 13368 10194 13404
rect 10138 12416 10194 12472
rect 9770 11600 9826 11656
rect 9586 9288 9642 9344
rect 9954 11872 10010 11928
rect 10046 11464 10102 11520
rect 10690 17856 10746 17912
rect 10322 12552 10378 12608
rect 10598 17040 10654 17096
rect 10506 16904 10562 16960
rect 10966 17040 11022 17096
rect 10817 16890 10873 16892
rect 10897 16890 10953 16892
rect 10977 16890 11033 16892
rect 11057 16890 11113 16892
rect 10817 16838 10843 16890
rect 10843 16838 10873 16890
rect 10897 16838 10907 16890
rect 10907 16838 10953 16890
rect 10977 16838 11023 16890
rect 11023 16838 11033 16890
rect 11057 16838 11087 16890
rect 11087 16838 11113 16890
rect 10817 16836 10873 16838
rect 10897 16836 10953 16838
rect 10977 16836 11033 16838
rect 11057 16836 11113 16838
rect 10817 15802 10873 15804
rect 10897 15802 10953 15804
rect 10977 15802 11033 15804
rect 11057 15802 11113 15804
rect 10817 15750 10843 15802
rect 10843 15750 10873 15802
rect 10897 15750 10907 15802
rect 10907 15750 10953 15802
rect 10977 15750 11023 15802
rect 11023 15750 11033 15802
rect 11057 15750 11087 15802
rect 11087 15750 11113 15802
rect 10817 15748 10873 15750
rect 10897 15748 10953 15750
rect 10977 15748 11033 15750
rect 11057 15748 11113 15750
rect 10782 15136 10838 15192
rect 10966 15136 11022 15192
rect 11058 14864 11114 14920
rect 10817 14714 10873 14716
rect 10897 14714 10953 14716
rect 10977 14714 11033 14716
rect 11057 14714 11113 14716
rect 10817 14662 10843 14714
rect 10843 14662 10873 14714
rect 10897 14662 10907 14714
rect 10907 14662 10953 14714
rect 10977 14662 11023 14714
rect 11023 14662 11033 14714
rect 11057 14662 11087 14714
rect 11087 14662 11113 14714
rect 10817 14660 10873 14662
rect 10897 14660 10953 14662
rect 10977 14660 11033 14662
rect 11057 14660 11113 14662
rect 10690 14340 10746 14376
rect 10690 14320 10692 14340
rect 10692 14320 10744 14340
rect 10744 14320 10746 14340
rect 10874 14320 10930 14376
rect 10598 14184 10654 14240
rect 11150 14476 11206 14512
rect 11150 14456 11152 14476
rect 11152 14456 11204 14476
rect 11204 14456 11206 14476
rect 11242 14184 11298 14240
rect 10817 13626 10873 13628
rect 10897 13626 10953 13628
rect 10977 13626 11033 13628
rect 11057 13626 11113 13628
rect 10817 13574 10843 13626
rect 10843 13574 10873 13626
rect 10897 13574 10907 13626
rect 10907 13574 10953 13626
rect 10977 13574 11023 13626
rect 11023 13574 11033 13626
rect 11057 13574 11087 13626
rect 11087 13574 11113 13626
rect 10817 13572 10873 13574
rect 10897 13572 10953 13574
rect 10977 13572 11033 13574
rect 11057 13572 11113 13574
rect 10506 12960 10562 13016
rect 10506 12416 10562 12472
rect 10230 12144 10286 12200
rect 10230 11328 10286 11384
rect 9954 10240 10010 10296
rect 10817 12538 10873 12540
rect 10897 12538 10953 12540
rect 10977 12538 11033 12540
rect 11057 12538 11113 12540
rect 10817 12486 10843 12538
rect 10843 12486 10873 12538
rect 10897 12486 10907 12538
rect 10907 12486 10953 12538
rect 10977 12486 11023 12538
rect 11023 12486 11033 12538
rect 11057 12486 11087 12538
rect 11087 12486 11113 12538
rect 10817 12484 10873 12486
rect 10897 12484 10953 12486
rect 10977 12484 11033 12486
rect 11057 12484 11113 12486
rect 11058 12144 11114 12200
rect 10966 11872 11022 11928
rect 10782 11600 10838 11656
rect 9954 9832 10010 9888
rect 9402 8744 9458 8800
rect 9494 8064 9550 8120
rect 9310 5480 9366 5536
rect 9218 5344 9274 5400
rect 9034 4936 9090 4992
rect 9862 8744 9918 8800
rect 9678 6840 9734 6896
rect 9586 6296 9642 6352
rect 9678 5888 9734 5944
rect 9586 5752 9642 5808
rect 9402 4800 9458 4856
rect 9678 4800 9734 4856
rect 9126 4392 9182 4448
rect 9586 4120 9642 4176
rect 8850 3304 8906 3360
rect 9034 3304 9090 3360
rect 8850 2352 8906 2408
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 9034 2080 9090 2136
rect 9494 3304 9550 3360
rect 9218 2624 9274 2680
rect 9862 5752 9918 5808
rect 10046 6996 10102 7032
rect 10046 6976 10048 6996
rect 10048 6976 10100 6996
rect 10100 6976 10102 6996
rect 10138 6876 10140 6896
rect 10140 6876 10192 6896
rect 10192 6876 10194 6896
rect 10138 6840 10194 6876
rect 10046 5616 10102 5672
rect 10230 6704 10286 6760
rect 10414 8064 10470 8120
rect 10817 11450 10873 11452
rect 10897 11450 10953 11452
rect 10977 11450 11033 11452
rect 11057 11450 11113 11452
rect 10817 11398 10843 11450
rect 10843 11398 10873 11450
rect 10897 11398 10907 11450
rect 10907 11398 10953 11450
rect 10977 11398 11023 11450
rect 11023 11398 11033 11450
rect 11057 11398 11087 11450
rect 11087 11398 11113 11450
rect 10817 11396 10873 11398
rect 10897 11396 10953 11398
rect 10977 11396 11033 11398
rect 11057 11396 11113 11398
rect 10782 10784 10838 10840
rect 10817 10362 10873 10364
rect 10897 10362 10953 10364
rect 10977 10362 11033 10364
rect 11057 10362 11113 10364
rect 10817 10310 10843 10362
rect 10843 10310 10873 10362
rect 10897 10310 10907 10362
rect 10907 10310 10953 10362
rect 10977 10310 11023 10362
rect 11023 10310 11033 10362
rect 11057 10310 11087 10362
rect 11087 10310 11113 10362
rect 10817 10308 10873 10310
rect 10897 10308 10953 10310
rect 10977 10308 11033 10310
rect 11057 10308 11113 10310
rect 11058 9696 11114 9752
rect 11334 12552 11390 12608
rect 11242 11500 11244 11520
rect 11244 11500 11296 11520
rect 11296 11500 11298 11520
rect 11242 11464 11298 11500
rect 11242 11328 11298 11384
rect 11242 10920 11298 10976
rect 11702 16360 11758 16416
rect 11794 15428 11850 15464
rect 11794 15408 11796 15428
rect 11796 15408 11848 15428
rect 11848 15408 11850 15428
rect 11794 15020 11850 15056
rect 11794 15000 11796 15020
rect 11796 15000 11848 15020
rect 11848 15000 11850 15020
rect 11702 14764 11704 14784
rect 11704 14764 11756 14784
rect 11756 14764 11758 14784
rect 11702 14728 11758 14764
rect 11794 13912 11850 13968
rect 11794 13268 11796 13288
rect 11796 13268 11848 13288
rect 11848 13268 11850 13288
rect 11794 13232 11850 13268
rect 11794 13096 11850 13152
rect 11610 12552 11666 12608
rect 11518 12280 11574 12336
rect 11794 12280 11850 12336
rect 11978 12552 12034 12608
rect 11978 12416 12034 12472
rect 11702 12144 11758 12200
rect 10598 8064 10654 8120
rect 10598 7792 10654 7848
rect 10817 9274 10873 9276
rect 10897 9274 10953 9276
rect 10977 9274 11033 9276
rect 11057 9274 11113 9276
rect 10817 9222 10843 9274
rect 10843 9222 10873 9274
rect 10897 9222 10907 9274
rect 10907 9222 10953 9274
rect 10977 9222 11023 9274
rect 11023 9222 11033 9274
rect 11057 9222 11087 9274
rect 11087 9222 11113 9274
rect 10817 9220 10873 9222
rect 10897 9220 10953 9222
rect 10977 9220 11033 9222
rect 11057 9220 11113 9222
rect 11334 9716 11390 9752
rect 11334 9696 11336 9716
rect 11336 9696 11388 9716
rect 11388 9696 11390 9716
rect 11702 10548 11704 10568
rect 11704 10548 11756 10568
rect 11756 10548 11758 10568
rect 11702 10512 11758 10548
rect 11702 10376 11758 10432
rect 11702 9868 11704 9888
rect 11704 9868 11756 9888
rect 11756 9868 11758 9888
rect 11702 9832 11758 9868
rect 10817 8186 10873 8188
rect 10897 8186 10953 8188
rect 10977 8186 11033 8188
rect 11057 8186 11113 8188
rect 10817 8134 10843 8186
rect 10843 8134 10873 8186
rect 10897 8134 10907 8186
rect 10907 8134 10953 8186
rect 10977 8134 11023 8186
rect 11023 8134 11033 8186
rect 11057 8134 11087 8186
rect 11087 8134 11113 8186
rect 10817 8132 10873 8134
rect 10897 8132 10953 8134
rect 10977 8132 11033 8134
rect 11057 8132 11113 8134
rect 11242 8492 11298 8528
rect 11242 8472 11244 8492
rect 11244 8472 11296 8492
rect 11296 8472 11298 8492
rect 11426 8336 11482 8392
rect 10598 7692 10600 7712
rect 10600 7692 10652 7712
rect 10652 7692 10654 7712
rect 10598 7656 10654 7692
rect 10782 7656 10838 7712
rect 10322 6568 10378 6624
rect 11150 7792 11206 7848
rect 10817 7098 10873 7100
rect 10897 7098 10953 7100
rect 10977 7098 11033 7100
rect 11057 7098 11113 7100
rect 10817 7046 10843 7098
rect 10843 7046 10873 7098
rect 10897 7046 10907 7098
rect 10907 7046 10953 7098
rect 10977 7046 11023 7098
rect 11023 7046 11033 7098
rect 11057 7046 11087 7098
rect 11087 7046 11113 7098
rect 10817 7044 10873 7046
rect 10897 7044 10953 7046
rect 10977 7044 11033 7046
rect 11057 7044 11113 7046
rect 10506 6024 10562 6080
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 10506 5616 10562 5672
rect 9862 4800 9918 4856
rect 10046 3884 10048 3904
rect 10048 3884 10100 3904
rect 10100 3884 10102 3904
rect 10046 3848 10102 3884
rect 9678 3304 9734 3360
rect 9770 3068 9772 3088
rect 9772 3068 9824 3088
rect 9824 3068 9826 3088
rect 9770 3032 9826 3068
rect 10046 2796 10048 2816
rect 10048 2796 10100 2816
rect 10100 2796 10102 2816
rect 10046 2760 10102 2796
rect 9954 2624 10010 2680
rect 10230 3848 10286 3904
rect 10230 3712 10286 3768
rect 10506 5344 10562 5400
rect 10414 3712 10470 3768
rect 10966 5752 11022 5808
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 11610 6876 11612 6896
rect 11612 6876 11664 6896
rect 11664 6876 11666 6896
rect 11610 6840 11666 6876
rect 11610 6740 11612 6760
rect 11612 6740 11664 6760
rect 11664 6740 11666 6760
rect 11610 6704 11666 6740
rect 11610 6568 11666 6624
rect 11334 5908 11390 5944
rect 11334 5888 11336 5908
rect 11336 5888 11388 5908
rect 11388 5888 11390 5908
rect 11334 5480 11390 5536
rect 11242 4936 11298 4992
rect 11334 4256 11390 4312
rect 11518 5072 11574 5128
rect 10782 3304 10838 3360
rect 10782 3168 10838 3224
rect 11242 3032 11298 3088
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 11426 3848 11482 3904
rect 11426 3032 11482 3088
rect 12070 10104 12126 10160
rect 12070 9832 12126 9888
rect 11978 8064 12034 8120
rect 12254 16496 12310 16552
rect 12254 15952 12310 16008
rect 12438 15272 12494 15328
rect 12438 14900 12440 14920
rect 12440 14900 12492 14920
rect 12492 14900 12494 14920
rect 12438 14864 12494 14900
rect 12438 13776 12494 13832
rect 12714 14048 12770 14104
rect 12622 12688 12678 12744
rect 12530 12280 12586 12336
rect 12438 12144 12494 12200
rect 12714 12552 12770 12608
rect 12898 13912 12954 13968
rect 12898 12552 12954 12608
rect 12806 12044 12808 12064
rect 12808 12044 12860 12064
rect 12860 12044 12862 12064
rect 12806 12008 12862 12044
rect 13358 17584 13414 17640
rect 13282 17434 13338 17436
rect 13362 17434 13418 17436
rect 13442 17434 13498 17436
rect 13522 17434 13578 17436
rect 13282 17382 13308 17434
rect 13308 17382 13338 17434
rect 13362 17382 13372 17434
rect 13372 17382 13418 17434
rect 13442 17382 13488 17434
rect 13488 17382 13498 17434
rect 13522 17382 13552 17434
rect 13552 17382 13578 17434
rect 13282 17380 13338 17382
rect 13362 17380 13418 17382
rect 13442 17380 13498 17382
rect 13522 17380 13578 17382
rect 13726 16768 13782 16824
rect 13726 16632 13782 16688
rect 13910 16632 13966 16688
rect 13282 16346 13338 16348
rect 13362 16346 13418 16348
rect 13442 16346 13498 16348
rect 13522 16346 13578 16348
rect 13282 16294 13308 16346
rect 13308 16294 13338 16346
rect 13362 16294 13372 16346
rect 13372 16294 13418 16346
rect 13442 16294 13488 16346
rect 13488 16294 13498 16346
rect 13522 16294 13552 16346
rect 13552 16294 13578 16346
rect 13282 16292 13338 16294
rect 13362 16292 13418 16294
rect 13442 16292 13498 16294
rect 13522 16292 13578 16294
rect 13282 15258 13338 15260
rect 13362 15258 13418 15260
rect 13442 15258 13498 15260
rect 13522 15258 13578 15260
rect 13282 15206 13308 15258
rect 13308 15206 13338 15258
rect 13362 15206 13372 15258
rect 13372 15206 13418 15258
rect 13442 15206 13488 15258
rect 13488 15206 13498 15258
rect 13522 15206 13552 15258
rect 13552 15206 13578 15258
rect 13282 15204 13338 15206
rect 13362 15204 13418 15206
rect 13442 15204 13498 15206
rect 13522 15204 13578 15206
rect 13174 15000 13230 15056
rect 13282 14170 13338 14172
rect 13362 14170 13418 14172
rect 13442 14170 13498 14172
rect 13522 14170 13578 14172
rect 13282 14118 13308 14170
rect 13308 14118 13338 14170
rect 13362 14118 13372 14170
rect 13372 14118 13418 14170
rect 13442 14118 13488 14170
rect 13488 14118 13498 14170
rect 13522 14118 13552 14170
rect 13552 14118 13578 14170
rect 13282 14116 13338 14118
rect 13362 14116 13418 14118
rect 13442 14116 13498 14118
rect 13522 14116 13578 14118
rect 13282 13082 13338 13084
rect 13362 13082 13418 13084
rect 13442 13082 13498 13084
rect 13522 13082 13578 13084
rect 13282 13030 13308 13082
rect 13308 13030 13338 13082
rect 13362 13030 13372 13082
rect 13372 13030 13418 13082
rect 13442 13030 13488 13082
rect 13488 13030 13498 13082
rect 13522 13030 13552 13082
rect 13552 13030 13578 13082
rect 13282 13028 13338 13030
rect 13362 13028 13418 13030
rect 13442 13028 13498 13030
rect 13522 13028 13578 13030
rect 13266 12688 13322 12744
rect 14094 16496 14150 16552
rect 13818 15408 13874 15464
rect 12714 11600 12770 11656
rect 12346 9832 12402 9888
rect 12254 8880 12310 8936
rect 12162 8608 12218 8664
rect 12438 9424 12494 9480
rect 12438 9152 12494 9208
rect 12622 9696 12678 9752
rect 13082 11328 13138 11384
rect 13282 11994 13338 11996
rect 13362 11994 13418 11996
rect 13442 11994 13498 11996
rect 13522 11994 13578 11996
rect 13282 11942 13308 11994
rect 13308 11942 13338 11994
rect 13362 11942 13372 11994
rect 13372 11942 13418 11994
rect 13442 11942 13488 11994
rect 13488 11942 13498 11994
rect 13522 11942 13552 11994
rect 13552 11942 13578 11994
rect 13282 11940 13338 11942
rect 13362 11940 13418 11942
rect 13442 11940 13498 11942
rect 13522 11940 13578 11942
rect 12990 11056 13046 11112
rect 12898 10140 12900 10160
rect 12900 10140 12952 10160
rect 12952 10140 12954 10160
rect 12898 10104 12954 10140
rect 12530 8744 12586 8800
rect 12438 8336 12494 8392
rect 12346 8200 12402 8256
rect 12346 7928 12402 7984
rect 12254 7792 12310 7848
rect 11978 7112 12034 7168
rect 11978 6704 12034 6760
rect 11794 4936 11850 4992
rect 11426 2644 11482 2680
rect 11426 2624 11428 2644
rect 11428 2624 11480 2644
rect 11480 2624 11482 2644
rect 10966 2216 11022 2272
rect 11794 2080 11850 2136
rect 12254 6840 12310 6896
rect 12162 4120 12218 4176
rect 12162 3848 12218 3904
rect 12806 9288 12862 9344
rect 13726 11736 13782 11792
rect 13910 13388 13966 13424
rect 13910 13368 13912 13388
rect 13912 13368 13964 13388
rect 13964 13368 13966 13388
rect 13910 12960 13966 13016
rect 13634 11192 13690 11248
rect 13542 11076 13598 11112
rect 13082 9288 13138 9344
rect 13542 11056 13544 11076
rect 13544 11056 13596 11076
rect 13596 11056 13598 11076
rect 13282 10906 13338 10908
rect 13362 10906 13418 10908
rect 13442 10906 13498 10908
rect 13522 10906 13578 10908
rect 13282 10854 13308 10906
rect 13308 10854 13338 10906
rect 13362 10854 13372 10906
rect 13372 10854 13418 10906
rect 13442 10854 13488 10906
rect 13488 10854 13498 10906
rect 13522 10854 13552 10906
rect 13552 10854 13578 10906
rect 13282 10852 13338 10854
rect 13362 10852 13418 10854
rect 13442 10852 13498 10854
rect 13522 10852 13578 10854
rect 13282 9818 13338 9820
rect 13362 9818 13418 9820
rect 13442 9818 13498 9820
rect 13522 9818 13578 9820
rect 13282 9766 13308 9818
rect 13308 9766 13338 9818
rect 13362 9766 13372 9818
rect 13372 9766 13418 9818
rect 13442 9766 13488 9818
rect 13488 9766 13498 9818
rect 13522 9766 13552 9818
rect 13552 9766 13578 9818
rect 13282 9764 13338 9766
rect 13362 9764 13418 9766
rect 13442 9764 13498 9766
rect 13522 9764 13578 9766
rect 12806 7384 12862 7440
rect 13282 8730 13338 8732
rect 13362 8730 13418 8732
rect 13442 8730 13498 8732
rect 13522 8730 13578 8732
rect 13282 8678 13308 8730
rect 13308 8678 13338 8730
rect 13362 8678 13372 8730
rect 13372 8678 13418 8730
rect 13442 8678 13488 8730
rect 13488 8678 13498 8730
rect 13522 8678 13552 8730
rect 13552 8678 13578 8730
rect 13282 8676 13338 8678
rect 13362 8676 13418 8678
rect 13442 8676 13498 8678
rect 13522 8676 13578 8678
rect 13818 10684 13820 10704
rect 13820 10684 13872 10704
rect 13872 10684 13874 10704
rect 13818 10648 13874 10684
rect 13910 9560 13966 9616
rect 13174 8472 13230 8528
rect 13542 8336 13598 8392
rect 12346 4800 12402 4856
rect 12438 2372 12494 2408
rect 12438 2352 12440 2372
rect 12440 2352 12492 2372
rect 12492 2352 12494 2372
rect 12622 3440 12678 3496
rect 12622 3304 12678 3360
rect 12898 6024 12954 6080
rect 13082 6296 13138 6352
rect 13282 7642 13338 7644
rect 13362 7642 13418 7644
rect 13442 7642 13498 7644
rect 13522 7642 13578 7644
rect 13282 7590 13308 7642
rect 13308 7590 13338 7642
rect 13362 7590 13372 7642
rect 13372 7590 13418 7642
rect 13442 7590 13488 7642
rect 13488 7590 13498 7642
rect 13522 7590 13552 7642
rect 13552 7590 13578 7642
rect 13282 7588 13338 7590
rect 13362 7588 13418 7590
rect 13442 7588 13498 7590
rect 13522 7588 13578 7590
rect 13634 7384 13690 7440
rect 13634 7248 13690 7304
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 13634 6160 13690 6216
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 13450 5228 13506 5264
rect 13450 5208 13452 5228
rect 13452 5208 13504 5228
rect 13504 5208 13506 5228
rect 13634 5092 13690 5128
rect 13634 5072 13636 5092
rect 13636 5072 13688 5092
rect 13688 5072 13690 5092
rect 12898 3032 12954 3088
rect 12898 2488 12954 2544
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 13266 4120 13322 4176
rect 13634 3848 13690 3904
rect 13266 3460 13322 3496
rect 13266 3440 13268 3460
rect 13268 3440 13320 3460
rect 13320 3440 13322 3460
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 13818 6704 13874 6760
rect 14186 9016 14242 9072
rect 14554 16088 14610 16144
rect 14370 11192 14426 11248
rect 14278 8336 14334 8392
rect 13634 2796 13636 2816
rect 13636 2796 13688 2816
rect 13688 2796 13690 2816
rect 13634 2760 13690 2796
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
rect 14094 4800 14150 4856
rect 14094 3848 14150 3904
rect 14094 3440 14150 3496
rect 14094 2896 14150 2952
rect 14830 12824 14886 12880
rect 14738 12688 14794 12744
rect 14462 8880 14518 8936
rect 14646 9988 14702 10024
rect 14646 9968 14648 9988
rect 14648 9968 14700 9988
rect 14700 9968 14702 9988
rect 15014 12688 15070 12744
rect 14462 3032 14518 3088
rect 14646 4548 14702 4584
rect 14646 4528 14648 4548
rect 14648 4528 14700 4548
rect 14700 4528 14702 4548
rect 14646 3712 14702 3768
rect 14922 5888 14978 5944
rect 14922 4120 14978 4176
rect 15198 10648 15254 10704
rect 16394 16088 16450 16144
rect 15106 9968 15162 10024
rect 15198 4936 15254 4992
rect 15566 3304 15622 3360
rect 16762 3984 16818 4040
<< metal3 >>
rect 0 19410 480 19440
rect 1485 19410 1551 19413
rect 0 19408 1551 19410
rect 0 19352 1490 19408
rect 1546 19352 1551 19408
rect 0 19350 1551 19352
rect 0 19320 480 19350
rect 1485 19347 1551 19350
rect 0 18458 480 18488
rect 1669 18458 1735 18461
rect 0 18456 1735 18458
rect 0 18400 1674 18456
rect 1730 18400 1735 18456
rect 0 18398 1735 18400
rect 0 18368 480 18398
rect 1669 18395 1735 18398
rect 8845 17914 8911 17917
rect 10685 17914 10751 17917
rect 8845 17912 10751 17914
rect 8845 17856 8850 17912
rect 8906 17856 10690 17912
rect 10746 17856 10751 17912
rect 8845 17854 10751 17856
rect 8845 17851 8911 17854
rect 10685 17851 10751 17854
rect 8753 17642 8819 17645
rect 13118 17642 13124 17644
rect 8753 17640 13124 17642
rect 8753 17584 8758 17640
rect 8814 17584 13124 17640
rect 8753 17582 13124 17584
rect 8753 17579 8819 17582
rect 13118 17580 13124 17582
rect 13188 17642 13194 17644
rect 13353 17642 13419 17645
rect 13188 17640 13419 17642
rect 13188 17584 13358 17640
rect 13414 17584 13419 17640
rect 13188 17582 13419 17584
rect 13188 17580 13194 17582
rect 13353 17579 13419 17582
rect 3409 17440 3729 17441
rect 0 17370 480 17400
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 17375 3729 17376
rect 8340 17440 8660 17441
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 17375 8660 17376
rect 13270 17440 13590 17441
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 13270 17375 13590 17376
rect 3049 17370 3115 17373
rect 0 17368 3115 17370
rect 0 17312 3054 17368
rect 3110 17312 3115 17368
rect 0 17310 3115 17312
rect 0 17280 480 17310
rect 3049 17307 3115 17310
rect 4981 17234 5047 17237
rect 9806 17234 9812 17236
rect 4981 17232 9812 17234
rect 4981 17176 4986 17232
rect 5042 17176 9812 17232
rect 4981 17174 9812 17176
rect 4981 17171 5047 17174
rect 9806 17172 9812 17174
rect 9876 17172 9882 17236
rect 8477 17098 8543 17101
rect 10593 17098 10659 17101
rect 8477 17096 10659 17098
rect 8477 17040 8482 17096
rect 8538 17040 10598 17096
rect 10654 17040 10659 17096
rect 8477 17038 10659 17040
rect 8477 17035 8543 17038
rect 10593 17035 10659 17038
rect 10961 17098 11027 17101
rect 11278 17098 11284 17100
rect 10961 17096 11284 17098
rect 10961 17040 10966 17096
rect 11022 17040 11284 17096
rect 10961 17038 11284 17040
rect 10961 17035 11027 17038
rect 11278 17036 11284 17038
rect 11348 17036 11354 17100
rect 7741 16962 7807 16965
rect 10501 16962 10567 16965
rect 7741 16960 10567 16962
rect 7741 16904 7746 16960
rect 7802 16904 10506 16960
rect 10562 16904 10567 16960
rect 7741 16902 10567 16904
rect 7741 16899 7807 16902
rect 10501 16899 10567 16902
rect 5874 16896 6194 16897
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6194 16896
rect 5874 16831 6194 16832
rect 10805 16896 11125 16897
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 16831 11125 16832
rect 3325 16826 3391 16829
rect 4286 16826 4292 16828
rect 3325 16824 4292 16826
rect 3325 16768 3330 16824
rect 3386 16768 4292 16824
rect 3325 16766 4292 16768
rect 3325 16763 3391 16766
rect 4286 16764 4292 16766
rect 4356 16764 4362 16828
rect 7741 16826 7807 16829
rect 8109 16826 8175 16829
rect 7741 16824 8175 16826
rect 7741 16768 7746 16824
rect 7802 16768 8114 16824
rect 8170 16768 8175 16824
rect 7741 16766 8175 16768
rect 7741 16763 7807 16766
rect 8109 16763 8175 16766
rect 8293 16826 8359 16829
rect 9581 16826 9647 16829
rect 8293 16824 9647 16826
rect 8293 16768 8298 16824
rect 8354 16768 9586 16824
rect 9642 16768 9647 16824
rect 8293 16766 9647 16768
rect 8293 16763 8359 16766
rect 9581 16763 9647 16766
rect 9990 16764 9996 16828
rect 10060 16826 10066 16828
rect 10133 16826 10199 16829
rect 10060 16824 10199 16826
rect 10060 16768 10138 16824
rect 10194 16768 10199 16824
rect 10060 16766 10199 16768
rect 10060 16764 10066 16766
rect 10133 16763 10199 16766
rect 13721 16826 13787 16829
rect 14038 16826 14044 16828
rect 13721 16824 14044 16826
rect 13721 16768 13726 16824
rect 13782 16768 14044 16824
rect 13721 16766 14044 16768
rect 13721 16763 13787 16766
rect 14038 16764 14044 16766
rect 14108 16764 14114 16828
rect 5349 16690 5415 16693
rect 13721 16690 13787 16693
rect 13905 16692 13971 16693
rect 5349 16688 13787 16690
rect 5349 16632 5354 16688
rect 5410 16632 13726 16688
rect 13782 16632 13787 16688
rect 5349 16630 13787 16632
rect 5349 16627 5415 16630
rect 13721 16627 13787 16630
rect 13854 16628 13860 16692
rect 13924 16690 13971 16692
rect 16520 16690 17000 16720
rect 13924 16688 17000 16690
rect 13966 16632 17000 16688
rect 13924 16630 17000 16632
rect 13924 16628 13971 16630
rect 13905 16627 13971 16628
rect 16520 16600 17000 16630
rect 5809 16554 5875 16557
rect 12249 16554 12315 16557
rect 5809 16552 12315 16554
rect 5809 16496 5814 16552
rect 5870 16496 12254 16552
rect 12310 16496 12315 16552
rect 5809 16494 12315 16496
rect 5809 16491 5875 16494
rect 12249 16491 12315 16494
rect 13670 16492 13676 16556
rect 13740 16554 13746 16556
rect 14089 16554 14155 16557
rect 13740 16552 14155 16554
rect 13740 16496 14094 16552
rect 14150 16496 14155 16552
rect 13740 16494 14155 16496
rect 13740 16492 13746 16494
rect 14089 16491 14155 16494
rect 0 16418 480 16448
rect 2773 16418 2839 16421
rect 0 16416 2839 16418
rect 0 16360 2778 16416
rect 2834 16360 2839 16416
rect 0 16358 2839 16360
rect 0 16328 480 16358
rect 2773 16355 2839 16358
rect 4153 16418 4219 16421
rect 8201 16418 8267 16421
rect 4153 16416 8267 16418
rect 4153 16360 4158 16416
rect 4214 16360 8206 16416
rect 8262 16360 8267 16416
rect 4153 16358 8267 16360
rect 4153 16355 4219 16358
rect 8201 16355 8267 16358
rect 9397 16418 9463 16421
rect 11697 16418 11763 16421
rect 9397 16416 11763 16418
rect 9397 16360 9402 16416
rect 9458 16360 11702 16416
rect 11758 16360 11763 16416
rect 9397 16358 11763 16360
rect 9397 16355 9463 16358
rect 11697 16355 11763 16358
rect 3409 16352 3729 16353
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 16287 3729 16288
rect 8340 16352 8660 16353
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 16287 8660 16288
rect 13270 16352 13590 16353
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 16287 13590 16288
rect 4705 16282 4771 16285
rect 7005 16282 7071 16285
rect 4705 16280 7071 16282
rect 4705 16224 4710 16280
rect 4766 16224 7010 16280
rect 7066 16224 7071 16280
rect 4705 16222 7071 16224
rect 4705 16219 4771 16222
rect 7005 16219 7071 16222
rect 7557 16282 7623 16285
rect 7966 16282 7972 16284
rect 7557 16280 7972 16282
rect 7557 16224 7562 16280
rect 7618 16224 7972 16280
rect 7557 16222 7972 16224
rect 7557 16219 7623 16222
rect 7966 16220 7972 16222
rect 8036 16220 8042 16284
rect 9254 16220 9260 16284
rect 9324 16282 9330 16284
rect 9489 16282 9555 16285
rect 9324 16280 9555 16282
rect 9324 16224 9494 16280
rect 9550 16224 9555 16280
rect 9324 16222 9555 16224
rect 9324 16220 9330 16222
rect 9489 16219 9555 16222
rect 9857 16282 9923 16285
rect 9990 16282 9996 16284
rect 9857 16280 9996 16282
rect 9857 16224 9862 16280
rect 9918 16224 9996 16280
rect 9857 16222 9996 16224
rect 9857 16219 9923 16222
rect 9990 16220 9996 16222
rect 10060 16220 10066 16284
rect 4889 16146 4955 16149
rect 6821 16146 6887 16149
rect 4889 16144 6887 16146
rect 4889 16088 4894 16144
rect 4950 16088 6826 16144
rect 6882 16088 6887 16144
rect 4889 16086 6887 16088
rect 4889 16083 4955 16086
rect 6821 16083 6887 16086
rect 7189 16146 7255 16149
rect 7741 16146 7807 16149
rect 7189 16144 7807 16146
rect 7189 16088 7194 16144
rect 7250 16088 7746 16144
rect 7802 16088 7807 16144
rect 7189 16086 7807 16088
rect 7189 16083 7255 16086
rect 7741 16083 7807 16086
rect 8150 16084 8156 16148
rect 8220 16146 8226 16148
rect 14549 16146 14615 16149
rect 16389 16146 16455 16149
rect 8220 16144 16455 16146
rect 8220 16088 14554 16144
rect 14610 16088 16394 16144
rect 16450 16088 16455 16144
rect 8220 16086 16455 16088
rect 8220 16084 8226 16086
rect 14549 16083 14615 16086
rect 16389 16083 16455 16086
rect 6545 16010 6611 16013
rect 12249 16010 12315 16013
rect 6545 16008 12315 16010
rect 6545 15952 6550 16008
rect 6606 15952 12254 16008
rect 12310 15952 12315 16008
rect 6545 15950 12315 15952
rect 6545 15947 6611 15950
rect 12249 15947 12315 15950
rect 5874 15808 6194 15809
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6194 15808
rect 5874 15743 6194 15744
rect 10805 15808 11125 15809
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 15743 11125 15744
rect 8109 15740 8175 15741
rect 8109 15738 8156 15740
rect 8064 15736 8156 15738
rect 8064 15680 8114 15736
rect 8064 15678 8156 15680
rect 8109 15676 8156 15678
rect 8220 15676 8226 15740
rect 9305 15738 9371 15741
rect 9622 15738 9628 15740
rect 9305 15736 9628 15738
rect 9305 15680 9310 15736
rect 9366 15680 9628 15736
rect 9305 15678 9628 15680
rect 8109 15675 8175 15676
rect 9305 15675 9371 15678
rect 9622 15676 9628 15678
rect 9692 15676 9698 15740
rect 9990 15676 9996 15740
rect 10060 15738 10066 15740
rect 10133 15738 10199 15741
rect 10060 15736 10199 15738
rect 10060 15680 10138 15736
rect 10194 15680 10199 15736
rect 10060 15678 10199 15680
rect 10060 15676 10066 15678
rect 10133 15675 10199 15678
rect 2681 15602 2747 15605
rect 2681 15600 13876 15602
rect 2681 15544 2686 15600
rect 2742 15544 13876 15600
rect 2681 15542 13876 15544
rect 2681 15539 2747 15542
rect 0 15466 480 15496
rect 13816 15469 13876 15542
rect 3601 15466 3667 15469
rect 0 15464 3667 15466
rect 0 15408 3606 15464
rect 3662 15408 3667 15464
rect 0 15406 3667 15408
rect 0 15376 480 15406
rect 3601 15403 3667 15406
rect 5717 15466 5783 15469
rect 6913 15466 6979 15469
rect 5717 15464 6979 15466
rect 5717 15408 5722 15464
rect 5778 15408 6918 15464
rect 6974 15408 6979 15464
rect 5717 15406 6979 15408
rect 5717 15403 5783 15406
rect 6913 15403 6979 15406
rect 7649 15466 7715 15469
rect 9765 15466 9831 15469
rect 11789 15466 11855 15469
rect 7649 15464 8954 15466
rect 7649 15408 7654 15464
rect 7710 15408 8954 15464
rect 7649 15406 8954 15408
rect 7649 15403 7715 15406
rect 3409 15264 3729 15265
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 15199 3729 15200
rect 8340 15264 8660 15265
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 15199 8660 15200
rect 8894 15194 8954 15406
rect 9765 15464 11855 15466
rect 9765 15408 9770 15464
rect 9826 15408 11794 15464
rect 11850 15408 11855 15464
rect 9765 15406 11855 15408
rect 9765 15403 9831 15406
rect 11789 15403 11855 15406
rect 13813 15464 13879 15469
rect 13813 15408 13818 15464
rect 13874 15408 13879 15464
rect 13813 15403 13879 15408
rect 9489 15330 9555 15333
rect 11830 15330 11836 15332
rect 9489 15328 11836 15330
rect 9489 15272 9494 15328
rect 9550 15272 11836 15328
rect 9489 15270 11836 15272
rect 9489 15267 9555 15270
rect 11830 15268 11836 15270
rect 11900 15330 11906 15332
rect 12433 15330 12499 15333
rect 11900 15328 12499 15330
rect 11900 15272 12438 15328
rect 12494 15272 12499 15328
rect 11900 15270 12499 15272
rect 11900 15268 11906 15270
rect 12433 15267 12499 15270
rect 13270 15264 13590 15265
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 15199 13590 15200
rect 10777 15194 10843 15197
rect 8894 15192 10843 15194
rect 8894 15136 10782 15192
rect 10838 15136 10843 15192
rect 8894 15134 10843 15136
rect 10777 15131 10843 15134
rect 10961 15194 11027 15197
rect 10961 15192 13186 15194
rect 10961 15136 10966 15192
rect 11022 15136 13186 15192
rect 10961 15134 13186 15136
rect 10961 15131 11027 15134
rect 13126 15061 13186 15134
rect 1301 15058 1367 15061
rect 7189 15058 7255 15061
rect 1301 15056 7255 15058
rect 1301 15000 1306 15056
rect 1362 15000 7194 15056
rect 7250 15000 7255 15056
rect 1301 14998 7255 15000
rect 1301 14995 1367 14998
rect 7189 14995 7255 14998
rect 7925 15058 7991 15061
rect 11789 15058 11855 15061
rect 7925 15056 11855 15058
rect 7925 15000 7930 15056
rect 7986 15000 11794 15056
rect 11850 15000 11855 15056
rect 7925 14998 11855 15000
rect 13126 15056 13235 15061
rect 13126 15000 13174 15056
rect 13230 15000 13235 15056
rect 13126 14998 13235 15000
rect 7925 14995 7991 14998
rect 11789 14995 11855 14998
rect 13169 14995 13235 14998
rect 6361 14922 6427 14925
rect 8385 14922 8451 14925
rect 6361 14920 8451 14922
rect 6361 14864 6366 14920
rect 6422 14864 8390 14920
rect 8446 14864 8451 14920
rect 6361 14862 8451 14864
rect 6361 14859 6427 14862
rect 8385 14859 8451 14862
rect 9949 14922 10015 14925
rect 11053 14922 11119 14925
rect 9949 14920 11119 14922
rect 9949 14864 9954 14920
rect 10010 14864 11058 14920
rect 11114 14864 11119 14920
rect 9949 14862 11119 14864
rect 9949 14859 10015 14862
rect 11053 14859 11119 14862
rect 12433 14922 12499 14925
rect 13670 14922 13676 14924
rect 12433 14920 13676 14922
rect 12433 14864 12438 14920
rect 12494 14864 13676 14920
rect 12433 14862 13676 14864
rect 12433 14859 12499 14862
rect 13670 14860 13676 14862
rect 13740 14860 13746 14924
rect 6637 14786 6703 14789
rect 7557 14786 7623 14789
rect 6637 14784 7623 14786
rect 6637 14728 6642 14784
rect 6698 14728 7562 14784
rect 7618 14728 7623 14784
rect 6637 14726 7623 14728
rect 6637 14723 6703 14726
rect 7557 14723 7623 14726
rect 7966 14724 7972 14788
rect 8036 14786 8042 14788
rect 9581 14786 9647 14789
rect 8036 14784 9647 14786
rect 8036 14728 9586 14784
rect 9642 14728 9647 14784
rect 8036 14726 9647 14728
rect 8036 14724 8042 14726
rect 9581 14723 9647 14726
rect 10133 14786 10199 14789
rect 10542 14786 10548 14788
rect 10133 14784 10548 14786
rect 10133 14728 10138 14784
rect 10194 14728 10548 14784
rect 10133 14726 10548 14728
rect 10133 14723 10199 14726
rect 10542 14724 10548 14726
rect 10612 14724 10618 14788
rect 11697 14786 11763 14789
rect 12934 14786 12940 14788
rect 11697 14784 12940 14786
rect 11697 14728 11702 14784
rect 11758 14728 12940 14784
rect 11697 14726 12940 14728
rect 11697 14723 11763 14726
rect 12934 14724 12940 14726
rect 13004 14724 13010 14788
rect 5874 14720 6194 14721
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6194 14720
rect 5874 14655 6194 14656
rect 10805 14720 11125 14721
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 14655 11125 14656
rect 9765 14650 9831 14653
rect 6272 14648 9831 14650
rect 6272 14592 9770 14648
rect 9826 14592 9831 14648
rect 6272 14590 9831 14592
rect 2405 14514 2471 14517
rect 6272 14514 6332 14590
rect 9765 14587 9831 14590
rect 2405 14512 6332 14514
rect 2405 14456 2410 14512
rect 2466 14456 6332 14512
rect 2405 14454 6332 14456
rect 8661 14514 8727 14517
rect 11145 14514 11211 14517
rect 11278 14514 11284 14516
rect 8661 14512 11284 14514
rect 8661 14456 8666 14512
rect 8722 14456 11150 14512
rect 11206 14456 11284 14512
rect 8661 14454 11284 14456
rect 2405 14451 2471 14454
rect 8661 14451 8727 14454
rect 11145 14451 11211 14454
rect 11278 14452 11284 14454
rect 11348 14514 11354 14516
rect 12198 14514 12204 14516
rect 11348 14454 12204 14514
rect 11348 14452 11354 14454
rect 12198 14452 12204 14454
rect 12268 14452 12274 14516
rect 0 14378 480 14408
rect 4245 14378 4311 14381
rect 0 14376 4311 14378
rect 0 14320 4250 14376
rect 4306 14320 4311 14376
rect 0 14318 4311 14320
rect 0 14288 480 14318
rect 4245 14315 4311 14318
rect 4889 14378 4955 14381
rect 10685 14378 10751 14381
rect 4889 14376 10751 14378
rect 4889 14320 4894 14376
rect 4950 14320 10690 14376
rect 10746 14320 10751 14376
rect 4889 14318 10751 14320
rect 4889 14315 4955 14318
rect 10685 14315 10751 14318
rect 10869 14378 10935 14381
rect 11646 14378 11652 14380
rect 10869 14376 11652 14378
rect 10869 14320 10874 14376
rect 10930 14320 11652 14376
rect 10869 14318 11652 14320
rect 10869 14315 10935 14318
rect 11646 14316 11652 14318
rect 11716 14316 11722 14380
rect 8937 14242 9003 14245
rect 10593 14242 10659 14245
rect 8937 14240 10659 14242
rect 8937 14184 8942 14240
rect 8998 14184 10598 14240
rect 10654 14184 10659 14240
rect 8937 14182 10659 14184
rect 8937 14179 9003 14182
rect 10593 14179 10659 14182
rect 11237 14242 11303 14245
rect 11462 14242 11468 14244
rect 11237 14240 11468 14242
rect 11237 14184 11242 14240
rect 11298 14184 11468 14240
rect 11237 14182 11468 14184
rect 11237 14179 11303 14182
rect 11462 14180 11468 14182
rect 11532 14180 11538 14244
rect 3409 14176 3729 14177
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 14111 3729 14112
rect 8340 14176 8660 14177
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 14111 8660 14112
rect 13270 14176 13590 14177
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 14111 13590 14112
rect 9438 14044 9444 14108
rect 9508 14106 9514 14108
rect 9581 14106 9647 14109
rect 9508 14104 9647 14106
rect 9508 14048 9586 14104
rect 9642 14048 9647 14104
rect 9508 14046 9647 14048
rect 9508 14044 9514 14046
rect 9581 14043 9647 14046
rect 9765 14106 9831 14109
rect 12709 14106 12775 14109
rect 9765 14104 12775 14106
rect 9765 14048 9770 14104
rect 9826 14048 12714 14104
rect 12770 14048 12775 14104
rect 9765 14046 12775 14048
rect 9765 14043 9831 14046
rect 12709 14043 12775 14046
rect 11789 13970 11855 13973
rect 3190 13968 11855 13970
rect 3190 13912 11794 13968
rect 11850 13912 11855 13968
rect 3190 13910 11855 13912
rect 3190 13837 3250 13910
rect 11789 13907 11855 13910
rect 12382 13908 12388 13972
rect 12452 13970 12458 13972
rect 12893 13970 12959 13973
rect 12452 13968 12959 13970
rect 12452 13912 12898 13968
rect 12954 13912 12959 13968
rect 12452 13910 12959 13912
rect 12452 13908 12458 13910
rect 12893 13907 12959 13910
rect 3141 13832 3250 13837
rect 3141 13776 3146 13832
rect 3202 13776 3250 13832
rect 3141 13774 3250 13776
rect 4245 13834 4311 13837
rect 5625 13834 5691 13837
rect 4245 13832 5691 13834
rect 4245 13776 4250 13832
rect 4306 13776 5630 13832
rect 5686 13776 5691 13832
rect 4245 13774 5691 13776
rect 3141 13771 3207 13774
rect 4245 13771 4311 13774
rect 5625 13771 5691 13774
rect 9070 13772 9076 13836
rect 9140 13834 9146 13836
rect 9397 13834 9463 13837
rect 9140 13832 9463 13834
rect 9140 13776 9402 13832
rect 9458 13776 9463 13832
rect 9140 13774 9463 13776
rect 9140 13772 9146 13774
rect 9397 13771 9463 13774
rect 10358 13772 10364 13836
rect 10428 13834 10434 13836
rect 12433 13834 12499 13837
rect 10428 13832 12499 13834
rect 10428 13776 12438 13832
rect 12494 13776 12499 13832
rect 10428 13774 12499 13776
rect 10428 13772 10434 13774
rect 12433 13771 12499 13774
rect 8201 13698 8267 13701
rect 9305 13698 9371 13701
rect 8201 13696 9371 13698
rect 8201 13640 8206 13696
rect 8262 13640 9310 13696
rect 9366 13640 9371 13696
rect 8201 13638 9371 13640
rect 8201 13635 8267 13638
rect 9305 13635 9371 13638
rect 5874 13632 6194 13633
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6194 13632
rect 5874 13567 6194 13568
rect 10805 13632 11125 13633
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 13567 11125 13568
rect 7097 13562 7163 13565
rect 7097 13560 10656 13562
rect 7097 13504 7102 13560
rect 7158 13504 10656 13560
rect 7097 13502 10656 13504
rect 7097 13499 7163 13502
rect 0 13426 480 13456
rect 10133 13426 10199 13429
rect 0 13424 10199 13426
rect 0 13368 10138 13424
rect 10194 13368 10199 13424
rect 0 13366 10199 13368
rect 10596 13426 10656 13502
rect 13905 13426 13971 13429
rect 10596 13424 13971 13426
rect 10596 13368 13910 13424
rect 13966 13368 13971 13424
rect 10596 13366 13971 13368
rect 0 13336 480 13366
rect 10133 13363 10199 13366
rect 13905 13363 13971 13366
rect 2221 13290 2287 13293
rect 6913 13290 6979 13293
rect 2221 13288 6979 13290
rect 2221 13232 2226 13288
rect 2282 13232 6918 13288
rect 6974 13232 6979 13288
rect 2221 13230 6979 13232
rect 2221 13227 2287 13230
rect 6913 13227 6979 13230
rect 7281 13290 7347 13293
rect 9673 13290 9739 13293
rect 7281 13288 9739 13290
rect 7281 13232 7286 13288
rect 7342 13232 9678 13288
rect 9734 13232 9739 13288
rect 7281 13230 9739 13232
rect 7281 13227 7347 13230
rect 9673 13227 9739 13230
rect 9857 13290 9923 13293
rect 11789 13290 11855 13293
rect 9857 13288 11855 13290
rect 9857 13232 9862 13288
rect 9918 13232 11794 13288
rect 11850 13232 11855 13288
rect 9857 13230 11855 13232
rect 9857 13227 9923 13230
rect 11789 13227 11855 13230
rect 13118 13228 13124 13292
rect 13188 13290 13194 13292
rect 13188 13230 13738 13290
rect 13188 13228 13194 13230
rect 8886 13092 8892 13156
rect 8956 13154 8962 13156
rect 9213 13154 9279 13157
rect 11789 13154 11855 13157
rect 8956 13152 9279 13154
rect 8956 13096 9218 13152
rect 9274 13096 9279 13152
rect 8956 13094 9279 13096
rect 8956 13092 8962 13094
rect 9213 13091 9279 13094
rect 10366 13152 11855 13154
rect 10366 13096 11794 13152
rect 11850 13096 11855 13152
rect 10366 13094 11855 13096
rect 3409 13088 3729 13089
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 13023 3729 13024
rect 8340 13088 8660 13089
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 13023 8660 13024
rect 4521 13018 4587 13021
rect 5165 13018 5231 13021
rect 4521 13016 5231 13018
rect 4521 12960 4526 13016
rect 4582 12960 5170 13016
rect 5226 12960 5231 13016
rect 4521 12958 5231 12960
rect 4521 12955 4587 12958
rect 5165 12955 5231 12958
rect 9254 12956 9260 13020
rect 9324 13018 9330 13020
rect 10366 13018 10426 13094
rect 11789 13091 11855 13094
rect 13270 13088 13590 13089
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 13023 13590 13024
rect 9324 12958 10426 13018
rect 10501 13018 10567 13021
rect 11278 13018 11284 13020
rect 10501 13016 11284 13018
rect 10501 12960 10506 13016
rect 10562 12960 11284 13016
rect 10501 12958 11284 12960
rect 9324 12956 9330 12958
rect 10501 12955 10567 12958
rect 11278 12956 11284 12958
rect 11348 12956 11354 13020
rect 13678 13018 13738 13230
rect 13905 13018 13971 13021
rect 13678 13016 13971 13018
rect 13678 12960 13910 13016
rect 13966 12960 13971 13016
rect 13678 12958 13971 12960
rect 13905 12955 13971 12958
rect 1393 12882 1459 12885
rect 14825 12882 14891 12885
rect 1393 12880 14891 12882
rect 1393 12824 1398 12880
rect 1454 12824 14830 12880
rect 14886 12824 14891 12880
rect 1393 12822 14891 12824
rect 1393 12819 1459 12822
rect 14825 12819 14891 12822
rect 2589 12746 2655 12749
rect 6545 12746 6611 12749
rect 9857 12746 9923 12749
rect 2589 12744 6424 12746
rect 2589 12688 2594 12744
rect 2650 12688 6424 12744
rect 2589 12686 6424 12688
rect 2589 12683 2655 12686
rect 6364 12610 6424 12686
rect 6545 12744 9923 12746
rect 6545 12688 6550 12744
rect 6606 12688 9862 12744
rect 9918 12688 9923 12744
rect 6545 12686 9923 12688
rect 6545 12683 6611 12686
rect 9857 12683 9923 12686
rect 10174 12684 10180 12748
rect 10244 12746 10250 12748
rect 11462 12746 11468 12748
rect 10244 12686 11468 12746
rect 10244 12684 10250 12686
rect 11462 12684 11468 12686
rect 11532 12684 11538 12748
rect 12617 12746 12683 12749
rect 13261 12746 13327 12749
rect 14038 12746 14044 12748
rect 12617 12744 12818 12746
rect 12617 12688 12622 12744
rect 12678 12688 12818 12744
rect 12617 12686 12818 12688
rect 12617 12683 12683 12686
rect 12758 12613 12818 12686
rect 13261 12744 14044 12746
rect 13261 12688 13266 12744
rect 13322 12688 14044 12744
rect 13261 12686 14044 12688
rect 13261 12683 13327 12686
rect 14038 12684 14044 12686
rect 14108 12684 14114 12748
rect 14733 12746 14799 12749
rect 15009 12746 15075 12749
rect 14733 12744 15075 12746
rect 14733 12688 14738 12744
rect 14794 12688 15014 12744
rect 15070 12688 15075 12744
rect 14733 12686 15075 12688
rect 14733 12683 14799 12686
rect 15009 12683 15075 12686
rect 8886 12610 8892 12612
rect 6364 12550 8892 12610
rect 8886 12548 8892 12550
rect 8956 12610 8962 12612
rect 9305 12610 9371 12613
rect 10317 12610 10383 12613
rect 8956 12550 9184 12610
rect 8956 12548 8962 12550
rect 5874 12544 6194 12545
rect 0 12474 480 12504
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6194 12544
rect 5874 12479 6194 12480
rect 2957 12474 3023 12477
rect 0 12472 3023 12474
rect 0 12416 2962 12472
rect 3018 12416 3023 12472
rect 0 12414 3023 12416
rect 0 12384 480 12414
rect 2957 12411 3023 12414
rect 7097 12474 7163 12477
rect 8845 12474 8911 12477
rect 7097 12472 8911 12474
rect 7097 12416 7102 12472
rect 7158 12416 8850 12472
rect 8906 12416 8911 12472
rect 7097 12414 8911 12416
rect 7097 12411 7163 12414
rect 8845 12411 8911 12414
rect 4705 12338 4771 12341
rect 7925 12338 7991 12341
rect 4705 12336 7991 12338
rect 4705 12280 4710 12336
rect 4766 12280 7930 12336
rect 7986 12280 7991 12336
rect 4705 12278 7991 12280
rect 9124 12338 9184 12550
rect 9305 12608 10383 12610
rect 9305 12552 9310 12608
rect 9366 12552 10322 12608
rect 10378 12552 10383 12608
rect 9305 12550 10383 12552
rect 9305 12547 9371 12550
rect 10317 12547 10383 12550
rect 11329 12610 11395 12613
rect 11462 12610 11468 12612
rect 11329 12608 11468 12610
rect 11329 12552 11334 12608
rect 11390 12552 11468 12608
rect 11329 12550 11468 12552
rect 11329 12547 11395 12550
rect 11462 12548 11468 12550
rect 11532 12548 11538 12612
rect 11605 12610 11671 12613
rect 11973 12612 12039 12613
rect 11605 12608 11898 12610
rect 11605 12552 11610 12608
rect 11666 12552 11898 12608
rect 11605 12550 11898 12552
rect 11605 12547 11671 12550
rect 10805 12544 11125 12545
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 12479 11125 12480
rect 9305 12476 9371 12477
rect 9254 12412 9260 12476
rect 9324 12474 9371 12476
rect 10133 12474 10199 12477
rect 10501 12474 10567 12477
rect 9324 12472 9416 12474
rect 9366 12416 9416 12472
rect 9324 12414 9416 12416
rect 10133 12472 10567 12474
rect 10133 12416 10138 12472
rect 10194 12416 10506 12472
rect 10562 12416 10567 12472
rect 10133 12414 10567 12416
rect 11838 12474 11898 12550
rect 11973 12608 12020 12612
rect 12084 12610 12090 12612
rect 11973 12552 11978 12608
rect 11973 12548 12020 12552
rect 12084 12550 12130 12610
rect 12709 12608 12818 12613
rect 12709 12552 12714 12608
rect 12770 12552 12818 12608
rect 12709 12550 12818 12552
rect 12893 12608 12959 12613
rect 12893 12552 12898 12608
rect 12954 12552 12959 12608
rect 12084 12548 12090 12550
rect 11973 12547 12039 12548
rect 12709 12547 12775 12550
rect 12893 12547 12959 12552
rect 11973 12474 12039 12477
rect 11838 12472 12039 12474
rect 11838 12416 11978 12472
rect 12034 12416 12039 12472
rect 11838 12414 12039 12416
rect 9324 12412 9371 12414
rect 9305 12411 9371 12412
rect 10133 12411 10199 12414
rect 10501 12411 10567 12414
rect 11973 12411 12039 12414
rect 11513 12338 11579 12341
rect 9124 12336 11579 12338
rect 9124 12280 11518 12336
rect 11574 12280 11579 12336
rect 9124 12278 11579 12280
rect 4705 12275 4771 12278
rect 7925 12275 7991 12278
rect 11513 12275 11579 12278
rect 11646 12276 11652 12340
rect 11716 12338 11722 12340
rect 11789 12338 11855 12341
rect 11716 12336 11855 12338
rect 11716 12280 11794 12336
rect 11850 12280 11855 12336
rect 11716 12278 11855 12280
rect 11716 12276 11722 12278
rect 11789 12275 11855 12278
rect 12525 12338 12591 12341
rect 12896 12338 12956 12547
rect 12525 12336 12956 12338
rect 12525 12280 12530 12336
rect 12586 12280 12956 12336
rect 12525 12278 12956 12280
rect 12525 12275 12591 12278
rect 2221 12202 2287 12205
rect 4613 12202 4679 12205
rect 7925 12202 7991 12205
rect 9990 12202 9996 12204
rect 2221 12200 4538 12202
rect 2221 12144 2226 12200
rect 2282 12144 4538 12200
rect 2221 12142 4538 12144
rect 2221 12139 2287 12142
rect 4478 12066 4538 12142
rect 4613 12200 9996 12202
rect 4613 12144 4618 12200
rect 4674 12144 7930 12200
rect 7986 12144 9996 12200
rect 4613 12142 9996 12144
rect 4613 12139 4679 12142
rect 7925 12139 7991 12142
rect 9990 12140 9996 12142
rect 10060 12140 10066 12204
rect 10225 12202 10291 12205
rect 11053 12202 11119 12205
rect 10225 12200 11119 12202
rect 10225 12144 10230 12200
rect 10286 12144 11058 12200
rect 11114 12144 11119 12200
rect 10225 12142 11119 12144
rect 10225 12139 10291 12142
rect 11053 12139 11119 12142
rect 11278 12140 11284 12204
rect 11348 12202 11354 12204
rect 11697 12202 11763 12205
rect 11348 12200 11763 12202
rect 11348 12144 11702 12200
rect 11758 12144 11763 12200
rect 11348 12142 11763 12144
rect 11348 12140 11354 12142
rect 11697 12139 11763 12142
rect 12433 12202 12499 12205
rect 12750 12202 12756 12204
rect 12433 12200 12756 12202
rect 12433 12144 12438 12200
rect 12494 12144 12756 12200
rect 12433 12142 12756 12144
rect 12433 12139 12499 12142
rect 12750 12140 12756 12142
rect 12820 12140 12826 12204
rect 8201 12066 8267 12069
rect 4478 12064 8267 12066
rect 4478 12008 8206 12064
rect 8262 12008 8267 12064
rect 4478 12006 8267 12008
rect 8201 12003 8267 12006
rect 8845 12066 8911 12069
rect 12801 12066 12867 12069
rect 8845 12064 12867 12066
rect 8845 12008 8850 12064
rect 8906 12008 12806 12064
rect 12862 12008 12867 12064
rect 8845 12006 12867 12008
rect 8845 12003 8911 12006
rect 12801 12003 12867 12006
rect 3409 12000 3729 12001
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 11935 3729 11936
rect 8340 12000 8660 12001
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 11935 8660 11936
rect 13270 12000 13590 12001
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 11935 13590 11936
rect 4337 11930 4403 11933
rect 4294 11928 4403 11930
rect 4294 11872 4342 11928
rect 4398 11872 4403 11928
rect 4294 11867 4403 11872
rect 5533 11930 5599 11933
rect 8201 11930 8267 11933
rect 9949 11932 10015 11933
rect 9949 11930 9996 11932
rect 5533 11928 8267 11930
rect 5533 11872 5538 11928
rect 5594 11872 8206 11928
rect 8262 11872 8267 11928
rect 5533 11870 8267 11872
rect 9904 11928 9996 11930
rect 9904 11872 9954 11928
rect 9904 11870 9996 11872
rect 5533 11867 5599 11870
rect 8201 11867 8267 11870
rect 9949 11868 9996 11870
rect 10060 11868 10066 11932
rect 10542 11868 10548 11932
rect 10612 11930 10618 11932
rect 10961 11930 11027 11933
rect 12566 11930 12572 11932
rect 10612 11928 12572 11930
rect 10612 11872 10966 11928
rect 11022 11872 12572 11928
rect 10612 11870 12572 11872
rect 10612 11868 10618 11870
rect 9949 11867 10015 11868
rect 10961 11867 11027 11870
rect 12566 11868 12572 11870
rect 12636 11868 12642 11932
rect 4294 11661 4354 11867
rect 6361 11794 6427 11797
rect 13721 11794 13787 11797
rect 13854 11794 13860 11796
rect 6361 11792 11668 11794
rect 6361 11736 6366 11792
rect 6422 11736 11668 11792
rect 6361 11734 11668 11736
rect 6361 11731 6427 11734
rect 4294 11656 4403 11661
rect 4294 11600 4342 11656
rect 4398 11600 4403 11656
rect 4294 11598 4403 11600
rect 4337 11595 4403 11598
rect 4889 11658 4955 11661
rect 5809 11658 5875 11661
rect 8477 11658 8543 11661
rect 4889 11656 8543 11658
rect 4889 11600 4894 11656
rect 4950 11600 5814 11656
rect 5870 11600 8482 11656
rect 8538 11600 8543 11656
rect 4889 11598 8543 11600
rect 4889 11595 4955 11598
rect 5809 11595 5875 11598
rect 8477 11595 8543 11598
rect 8661 11658 8727 11661
rect 9622 11658 9628 11660
rect 8661 11656 9628 11658
rect 8661 11600 8666 11656
rect 8722 11600 9628 11656
rect 8661 11598 9628 11600
rect 8661 11595 8727 11598
rect 9622 11596 9628 11598
rect 9692 11658 9698 11660
rect 9765 11658 9831 11661
rect 9692 11656 9831 11658
rect 9692 11600 9770 11656
rect 9826 11600 9831 11656
rect 9692 11598 9831 11600
rect 9692 11596 9698 11598
rect 9765 11595 9831 11598
rect 10777 11658 10843 11661
rect 11462 11658 11468 11660
rect 10777 11656 11468 11658
rect 10777 11600 10782 11656
rect 10838 11600 11468 11656
rect 10777 11598 11468 11600
rect 10777 11595 10843 11598
rect 11462 11596 11468 11598
rect 11532 11596 11538 11660
rect 6269 11522 6335 11525
rect 9581 11522 9647 11525
rect 6269 11520 9647 11522
rect 6269 11464 6274 11520
rect 6330 11464 9586 11520
rect 9642 11464 9647 11520
rect 6269 11462 9647 11464
rect 6269 11459 6335 11462
rect 9581 11459 9647 11462
rect 10041 11520 10107 11525
rect 10041 11464 10046 11520
rect 10102 11464 10107 11520
rect 10041 11459 10107 11464
rect 11237 11522 11303 11525
rect 11608 11522 11668 11734
rect 13721 11792 13860 11794
rect 13721 11736 13726 11792
rect 13782 11736 13860 11792
rect 13721 11734 13860 11736
rect 13721 11731 13787 11734
rect 13854 11732 13860 11734
rect 13924 11732 13930 11796
rect 12709 11658 12775 11661
rect 11237 11520 11668 11522
rect 11237 11464 11242 11520
rect 11298 11464 11668 11520
rect 11237 11462 11668 11464
rect 11792 11656 12775 11658
rect 11792 11600 12714 11656
rect 12770 11600 12775 11656
rect 11792 11598 12775 11600
rect 11237 11459 11303 11462
rect 5874 11456 6194 11457
rect 0 11386 480 11416
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6194 11456
rect 5874 11391 6194 11392
rect 3049 11386 3115 11389
rect 0 11384 3115 11386
rect 0 11328 3054 11384
rect 3110 11328 3115 11384
rect 0 11326 3115 11328
rect 0 11296 480 11326
rect 3049 11323 3115 11326
rect 7005 11386 7071 11389
rect 10044 11386 10104 11459
rect 10805 11456 11125 11457
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 11391 11125 11392
rect 10225 11388 10291 11389
rect 7005 11384 10104 11386
rect 7005 11328 7010 11384
rect 7066 11328 10104 11384
rect 7005 11326 10104 11328
rect 7005 11323 7071 11326
rect 10174 11324 10180 11388
rect 10244 11386 10291 11388
rect 11237 11386 11303 11389
rect 11792 11386 11852 11598
rect 12709 11595 12775 11598
rect 10244 11384 10336 11386
rect 10286 11328 10336 11384
rect 10244 11326 10336 11328
rect 11237 11384 11852 11386
rect 11237 11328 11242 11384
rect 11298 11328 11852 11384
rect 11237 11326 11852 11328
rect 10244 11324 10291 11326
rect 10225 11323 10291 11324
rect 11237 11323 11303 11326
rect 12934 11324 12940 11388
rect 13004 11386 13010 11388
rect 13077 11386 13143 11389
rect 13004 11384 13143 11386
rect 13004 11328 13082 11384
rect 13138 11328 13143 11384
rect 13004 11326 13143 11328
rect 13004 11324 13010 11326
rect 13077 11323 13143 11326
rect 1945 11250 2011 11253
rect 13629 11250 13695 11253
rect 1945 11248 13695 11250
rect 1945 11192 1950 11248
rect 2006 11192 13634 11248
rect 13690 11192 13695 11248
rect 1945 11190 13695 11192
rect 1945 11187 2011 11190
rect 13629 11187 13695 11190
rect 13854 11188 13860 11252
rect 13924 11250 13930 11252
rect 14365 11250 14431 11253
rect 13924 11248 14431 11250
rect 13924 11192 14370 11248
rect 14426 11192 14431 11248
rect 13924 11190 14431 11192
rect 13924 11188 13930 11190
rect 14365 11187 14431 11190
rect 5809 11114 5875 11117
rect 8661 11114 8727 11117
rect 5809 11112 8727 11114
rect 5809 11056 5814 11112
rect 5870 11056 8666 11112
rect 8722 11056 8727 11112
rect 5809 11054 8727 11056
rect 5809 11051 5875 11054
rect 8661 11051 8727 11054
rect 8937 11114 9003 11117
rect 12985 11114 13051 11117
rect 13537 11114 13603 11117
rect 8937 11112 11530 11114
rect 8937 11056 8942 11112
rect 8998 11056 11530 11112
rect 8937 11054 11530 11056
rect 8937 11051 9003 11054
rect 9029 10980 9095 10981
rect 9029 10978 9076 10980
rect 8984 10976 9076 10978
rect 8984 10920 9034 10976
rect 8984 10918 9076 10920
rect 9029 10916 9076 10918
rect 9140 10916 9146 10980
rect 10174 10916 10180 10980
rect 10244 10978 10250 10980
rect 11237 10978 11303 10981
rect 10244 10976 11303 10978
rect 10244 10920 11242 10976
rect 11298 10920 11303 10976
rect 10244 10918 11303 10920
rect 11470 10978 11530 11054
rect 11976 11112 13603 11114
rect 11976 11056 12990 11112
rect 13046 11056 13542 11112
rect 13598 11056 13603 11112
rect 11976 11054 13603 11056
rect 11976 10978 12036 11054
rect 12985 11051 13051 11054
rect 13537 11051 13603 11054
rect 11470 10918 12036 10978
rect 10244 10916 10250 10918
rect 9029 10915 9095 10916
rect 11237 10915 11303 10918
rect 3409 10912 3729 10913
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 10847 3729 10848
rect 8340 10912 8660 10913
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 10847 8660 10848
rect 13270 10912 13590 10913
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 10847 13590 10848
rect 10777 10842 10843 10845
rect 12382 10842 12388 10844
rect 10777 10840 12388 10842
rect 10777 10784 10782 10840
rect 10838 10784 12388 10840
rect 10777 10782 12388 10784
rect 10777 10779 10843 10782
rect 12382 10780 12388 10782
rect 12452 10780 12458 10844
rect 6637 10706 6703 10709
rect 13813 10706 13879 10709
rect 6637 10704 13879 10706
rect 6637 10648 6642 10704
rect 6698 10648 13818 10704
rect 13874 10648 13879 10704
rect 6637 10646 13879 10648
rect 6637 10643 6703 10646
rect 13813 10643 13879 10646
rect 14406 10644 14412 10708
rect 14476 10706 14482 10708
rect 15193 10706 15259 10709
rect 14476 10704 15259 10706
rect 14476 10648 15198 10704
rect 15254 10648 15259 10704
rect 14476 10646 15259 10648
rect 14476 10644 14482 10646
rect 15193 10643 15259 10646
rect 9397 10572 9463 10573
rect 9397 10570 9444 10572
rect 9352 10568 9444 10570
rect 9352 10512 9402 10568
rect 9352 10510 9444 10512
rect 9397 10508 9444 10510
rect 9508 10508 9514 10572
rect 9581 10570 9647 10573
rect 11697 10572 11763 10573
rect 11646 10570 11652 10572
rect 9581 10568 11652 10570
rect 11716 10570 11763 10572
rect 11716 10568 11808 10570
rect 9581 10512 9586 10568
rect 9642 10512 11652 10568
rect 11758 10512 11808 10568
rect 9581 10510 11652 10512
rect 9397 10507 9463 10508
rect 9581 10507 9647 10510
rect 11646 10508 11652 10510
rect 11716 10510 11808 10512
rect 11716 10508 11763 10510
rect 11697 10507 11763 10508
rect 0 10434 480 10464
rect 1853 10434 1919 10437
rect 0 10432 1919 10434
rect 0 10376 1858 10432
rect 1914 10376 1919 10432
rect 0 10374 1919 10376
rect 0 10344 480 10374
rect 1853 10371 1919 10374
rect 7465 10434 7531 10437
rect 8201 10434 8267 10437
rect 7465 10432 8267 10434
rect 7465 10376 7470 10432
rect 7526 10376 8206 10432
rect 8262 10376 8267 10432
rect 7465 10374 8267 10376
rect 7465 10371 7531 10374
rect 8201 10371 8267 10374
rect 11697 10434 11763 10437
rect 12014 10434 12020 10436
rect 11697 10432 12020 10434
rect 11697 10376 11702 10432
rect 11758 10376 12020 10432
rect 11697 10374 12020 10376
rect 11697 10371 11763 10374
rect 12014 10372 12020 10374
rect 12084 10372 12090 10436
rect 5874 10368 6194 10369
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6194 10368
rect 5874 10303 6194 10304
rect 10805 10368 11125 10369
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 10303 11125 10304
rect 8201 10298 8267 10301
rect 9949 10298 10015 10301
rect 8201 10296 10015 10298
rect 8201 10240 8206 10296
rect 8262 10240 9954 10296
rect 10010 10240 10015 10296
rect 8201 10238 10015 10240
rect 8201 10235 8267 10238
rect 9949 10235 10015 10238
rect 12065 10162 12131 10165
rect 12198 10162 12204 10164
rect 5214 10160 12204 10162
rect 5214 10104 12070 10160
rect 12126 10104 12204 10160
rect 5214 10102 12204 10104
rect 2865 10026 2931 10029
rect 4797 10026 4863 10029
rect 5214 10026 5274 10102
rect 12065 10099 12131 10102
rect 12198 10100 12204 10102
rect 12268 10100 12274 10164
rect 12893 10162 12959 10165
rect 13670 10162 13676 10164
rect 12893 10160 13676 10162
rect 12893 10104 12898 10160
rect 12954 10104 13676 10160
rect 12893 10102 13676 10104
rect 12893 10099 12959 10102
rect 13670 10100 13676 10102
rect 13740 10100 13746 10164
rect 2865 10024 5274 10026
rect 2865 9968 2870 10024
rect 2926 9968 4802 10024
rect 4858 9968 5274 10024
rect 2865 9966 5274 9968
rect 6545 10026 6611 10029
rect 14641 10026 14707 10029
rect 6545 10024 14707 10026
rect 6545 9968 6550 10024
rect 6606 9968 14646 10024
rect 14702 9968 14707 10024
rect 6545 9966 14707 9968
rect 2865 9963 2931 9966
rect 4797 9963 4863 9966
rect 6545 9963 6611 9966
rect 14641 9963 14707 9966
rect 15101 10026 15167 10029
rect 16520 10026 17000 10056
rect 15101 10024 17000 10026
rect 15101 9968 15106 10024
rect 15162 9968 17000 10024
rect 15101 9966 17000 9968
rect 15101 9963 15167 9966
rect 16520 9936 17000 9966
rect 5073 9890 5139 9893
rect 5533 9890 5599 9893
rect 7649 9890 7715 9893
rect 5073 9888 7715 9890
rect 5073 9832 5078 9888
rect 5134 9832 5538 9888
rect 5594 9832 7654 9888
rect 7710 9832 7715 9888
rect 5073 9830 7715 9832
rect 5073 9827 5139 9830
rect 5533 9827 5599 9830
rect 7649 9827 7715 9830
rect 9949 9890 10015 9893
rect 11697 9890 11763 9893
rect 9949 9888 11763 9890
rect 9949 9832 9954 9888
rect 10010 9832 11702 9888
rect 11758 9832 11763 9888
rect 9949 9830 11763 9832
rect 9949 9827 10015 9830
rect 11697 9827 11763 9830
rect 12065 9890 12131 9893
rect 12341 9890 12407 9893
rect 12065 9888 12407 9890
rect 12065 9832 12070 9888
rect 12126 9832 12346 9888
rect 12402 9832 12407 9888
rect 12065 9830 12407 9832
rect 12065 9827 12131 9830
rect 12341 9827 12407 9830
rect 3409 9824 3729 9825
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 9759 3729 9760
rect 8340 9824 8660 9825
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 9759 8660 9760
rect 13270 9824 13590 9825
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 9759 13590 9760
rect 11053 9754 11119 9757
rect 9630 9752 11119 9754
rect 9630 9696 11058 9752
rect 11114 9696 11119 9752
rect 9630 9694 11119 9696
rect 7649 9618 7715 9621
rect 2270 9616 7715 9618
rect 2270 9560 7654 9616
rect 7710 9560 7715 9616
rect 2270 9558 7715 9560
rect 0 9482 480 9512
rect 2270 9482 2330 9558
rect 7649 9555 7715 9558
rect 8017 9618 8083 9621
rect 9630 9618 9690 9694
rect 11053 9691 11119 9694
rect 11329 9754 11395 9757
rect 12617 9756 12683 9757
rect 12566 9754 12572 9756
rect 11329 9752 12572 9754
rect 12636 9754 12683 9756
rect 12636 9752 12764 9754
rect 11329 9696 11334 9752
rect 11390 9696 12572 9752
rect 12678 9696 12764 9752
rect 11329 9694 12572 9696
rect 11329 9691 11395 9694
rect 12566 9692 12572 9694
rect 12636 9694 12764 9696
rect 12636 9692 12683 9694
rect 12617 9691 12683 9692
rect 8017 9616 9690 9618
rect 8017 9560 8022 9616
rect 8078 9560 9690 9616
rect 8017 9558 9690 9560
rect 8017 9555 8083 9558
rect 9990 9556 9996 9620
rect 10060 9618 10066 9620
rect 13118 9618 13124 9620
rect 10060 9558 13124 9618
rect 10060 9556 10066 9558
rect 13118 9556 13124 9558
rect 13188 9618 13194 9620
rect 13905 9618 13971 9621
rect 13188 9616 13971 9618
rect 13188 9560 13910 9616
rect 13966 9560 13971 9616
rect 13188 9558 13971 9560
rect 13188 9556 13194 9558
rect 13905 9555 13971 9558
rect 0 9422 2330 9482
rect 2497 9482 2563 9485
rect 12433 9482 12499 9485
rect 2497 9480 12499 9482
rect 2497 9424 2502 9480
rect 2558 9424 12438 9480
rect 12494 9424 12499 9480
rect 2497 9422 12499 9424
rect 0 9392 480 9422
rect 2497 9419 2563 9422
rect 12433 9419 12499 9422
rect 7097 9346 7163 9349
rect 8109 9346 8175 9349
rect 7097 9344 8175 9346
rect 7097 9288 7102 9344
rect 7158 9288 8114 9344
rect 8170 9288 8175 9344
rect 7097 9286 8175 9288
rect 7097 9283 7163 9286
rect 8109 9283 8175 9286
rect 8385 9346 8451 9349
rect 8886 9346 8892 9348
rect 8385 9344 8892 9346
rect 8385 9288 8390 9344
rect 8446 9288 8892 9344
rect 8385 9286 8892 9288
rect 8385 9283 8451 9286
rect 8886 9284 8892 9286
rect 8956 9346 8962 9348
rect 9581 9346 9647 9349
rect 8956 9344 9647 9346
rect 8956 9288 9586 9344
rect 9642 9288 9647 9344
rect 8956 9286 9647 9288
rect 8956 9284 8962 9286
rect 9581 9283 9647 9286
rect 9768 9286 10426 9346
rect 5874 9280 6194 9281
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6194 9280
rect 5874 9215 6194 9216
rect 2957 9210 3023 9213
rect 5625 9210 5691 9213
rect 2957 9208 5691 9210
rect 2957 9152 2962 9208
rect 3018 9152 5630 9208
rect 5686 9152 5691 9208
rect 2957 9150 5691 9152
rect 2957 9147 3023 9150
rect 5625 9147 5691 9150
rect 7557 9210 7623 9213
rect 8661 9210 8727 9213
rect 7557 9208 8727 9210
rect 7557 9152 7562 9208
rect 7618 9152 8666 9208
rect 8722 9152 8727 9208
rect 7557 9150 8727 9152
rect 7557 9147 7623 9150
rect 8661 9147 8727 9150
rect 5717 9074 5783 9077
rect 9768 9074 9828 9286
rect 5717 9072 9828 9074
rect 5717 9016 5722 9072
rect 5778 9016 9828 9072
rect 5717 9014 9828 9016
rect 10366 9074 10426 9286
rect 11278 9284 11284 9348
rect 11348 9346 11354 9348
rect 12801 9346 12867 9349
rect 11348 9344 12867 9346
rect 11348 9288 12806 9344
rect 12862 9288 12867 9344
rect 11348 9286 12867 9288
rect 11348 9284 11354 9286
rect 12801 9283 12867 9286
rect 13077 9348 13143 9349
rect 13077 9344 13124 9348
rect 13188 9346 13194 9348
rect 13077 9288 13082 9344
rect 13077 9284 13124 9288
rect 13188 9286 13234 9346
rect 13188 9284 13194 9286
rect 13077 9283 13143 9284
rect 10805 9280 11125 9281
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 9215 11125 9216
rect 12433 9210 12499 9213
rect 12934 9210 12940 9212
rect 12433 9208 12940 9210
rect 12433 9152 12438 9208
rect 12494 9152 12940 9208
rect 12433 9150 12940 9152
rect 12433 9147 12499 9150
rect 12934 9148 12940 9150
rect 13004 9148 13010 9212
rect 14181 9074 14247 9077
rect 10366 9072 14247 9074
rect 10366 9016 14186 9072
rect 14242 9016 14247 9072
rect 10366 9014 14247 9016
rect 5717 9011 5783 9014
rect 14181 9011 14247 9014
rect 4521 8940 4587 8941
rect 4470 8876 4476 8940
rect 4540 8938 4587 8940
rect 4981 8938 5047 8941
rect 7189 8938 7255 8941
rect 4540 8936 4632 8938
rect 4582 8880 4632 8936
rect 4540 8878 4632 8880
rect 4981 8936 7255 8938
rect 4981 8880 4986 8936
rect 5042 8880 7194 8936
rect 7250 8880 7255 8936
rect 4981 8878 7255 8880
rect 4540 8876 4587 8878
rect 4521 8875 4587 8876
rect 4981 8875 5047 8878
rect 7189 8875 7255 8878
rect 7465 8938 7531 8941
rect 10542 8938 10548 8940
rect 7465 8936 10548 8938
rect 7465 8880 7470 8936
rect 7526 8880 10548 8936
rect 7465 8878 10548 8880
rect 7465 8875 7531 8878
rect 10542 8876 10548 8878
rect 10612 8938 10618 8940
rect 11278 8938 11284 8940
rect 10612 8878 11284 8938
rect 10612 8876 10618 8878
rect 11278 8876 11284 8878
rect 11348 8876 11354 8940
rect 11646 8876 11652 8940
rect 11716 8938 11722 8940
rect 12249 8938 12315 8941
rect 12382 8938 12388 8940
rect 11716 8936 12388 8938
rect 11716 8880 12254 8936
rect 12310 8880 12388 8936
rect 11716 8878 12388 8880
rect 11716 8876 11722 8878
rect 12249 8875 12315 8878
rect 12382 8876 12388 8878
rect 12452 8876 12458 8940
rect 14038 8876 14044 8940
rect 14108 8938 14114 8940
rect 14457 8938 14523 8941
rect 14108 8936 14523 8938
rect 14108 8880 14462 8936
rect 14518 8880 14523 8936
rect 14108 8878 14523 8880
rect 14108 8876 14114 8878
rect 14457 8875 14523 8878
rect 9397 8802 9463 8805
rect 9857 8802 9923 8805
rect 9397 8800 9923 8802
rect 9397 8744 9402 8800
rect 9458 8744 9862 8800
rect 9918 8744 9923 8800
rect 9397 8742 9923 8744
rect 9397 8739 9463 8742
rect 9857 8739 9923 8742
rect 12382 8740 12388 8804
rect 12452 8802 12458 8804
rect 12525 8802 12591 8805
rect 12452 8800 12591 8802
rect 12452 8744 12530 8800
rect 12586 8744 12591 8800
rect 12452 8742 12591 8744
rect 12452 8740 12458 8742
rect 12525 8739 12591 8742
rect 3409 8736 3729 8737
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 8671 3729 8672
rect 8340 8736 8660 8737
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 8671 8660 8672
rect 13270 8736 13590 8737
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 8671 13590 8672
rect 4337 8666 4403 8669
rect 5809 8666 5875 8669
rect 4337 8664 5875 8666
rect 4337 8608 4342 8664
rect 4398 8608 5814 8664
rect 5870 8608 5875 8664
rect 4337 8606 5875 8608
rect 4337 8603 4403 8606
rect 5809 8603 5875 8606
rect 9622 8604 9628 8668
rect 9692 8666 9698 8668
rect 12157 8666 12223 8669
rect 12750 8666 12756 8668
rect 9692 8606 11484 8666
rect 9692 8604 9698 8606
rect 3877 8530 3943 8533
rect 9438 8530 9444 8532
rect 3877 8528 9444 8530
rect 3877 8472 3882 8528
rect 3938 8472 9444 8528
rect 3877 8470 9444 8472
rect 3877 8467 3943 8470
rect 9438 8468 9444 8470
rect 9508 8468 9514 8532
rect 11237 8530 11303 8533
rect 10734 8528 11303 8530
rect 10734 8472 11242 8528
rect 11298 8472 11303 8528
rect 10734 8470 11303 8472
rect 0 8394 480 8424
rect 1209 8394 1275 8397
rect 0 8392 1275 8394
rect 0 8336 1214 8392
rect 1270 8336 1275 8392
rect 0 8334 1275 8336
rect 0 8304 480 8334
rect 1209 8331 1275 8334
rect 3601 8394 3667 8397
rect 4153 8394 4219 8397
rect 10734 8394 10794 8470
rect 11237 8467 11303 8470
rect 11424 8530 11484 8606
rect 12157 8664 12756 8666
rect 12157 8608 12162 8664
rect 12218 8608 12756 8664
rect 12157 8606 12756 8608
rect 12157 8603 12223 8606
rect 12750 8604 12756 8606
rect 12820 8604 12826 8668
rect 13169 8530 13235 8533
rect 11424 8528 13235 8530
rect 11424 8472 13174 8528
rect 13230 8472 13235 8528
rect 11424 8470 13235 8472
rect 11424 8397 11484 8470
rect 13169 8467 13235 8470
rect 3601 8392 4219 8394
rect 3601 8336 3606 8392
rect 3662 8336 4158 8392
rect 4214 8336 4219 8392
rect 3601 8334 4219 8336
rect 3601 8331 3667 8334
rect 4153 8331 4219 8334
rect 4294 8334 10794 8394
rect 11421 8392 11487 8397
rect 12433 8396 12499 8397
rect 12382 8394 12388 8396
rect 11421 8336 11426 8392
rect 11482 8336 11487 8392
rect 1209 8258 1275 8261
rect 4294 8258 4354 8334
rect 11421 8331 11487 8336
rect 12342 8334 12388 8394
rect 12452 8392 12499 8396
rect 12494 8336 12499 8392
rect 12382 8332 12388 8334
rect 12452 8332 12499 8336
rect 12433 8331 12499 8332
rect 13537 8394 13603 8397
rect 14273 8394 14339 8397
rect 13537 8392 14339 8394
rect 13537 8336 13542 8392
rect 13598 8336 14278 8392
rect 14334 8336 14339 8392
rect 13537 8334 14339 8336
rect 13537 8331 13603 8334
rect 14273 8331 14339 8334
rect 1209 8256 4354 8258
rect 1209 8200 1214 8256
rect 1270 8200 4354 8256
rect 1209 8198 4354 8200
rect 9213 8260 9279 8261
rect 12341 8260 12407 8261
rect 9213 8256 9260 8260
rect 9324 8258 9330 8260
rect 9213 8200 9218 8256
rect 1209 8195 1275 8198
rect 9213 8196 9260 8200
rect 9324 8198 9370 8258
rect 9324 8196 9330 8198
rect 9438 8196 9444 8260
rect 9508 8258 9514 8260
rect 12341 8258 12388 8260
rect 9508 8198 10656 8258
rect 12296 8256 12388 8258
rect 12296 8200 12346 8256
rect 12296 8198 12388 8200
rect 9508 8196 9514 8198
rect 9213 8195 9279 8196
rect 5874 8192 6194 8193
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6194 8192
rect 5874 8127 6194 8128
rect 10596 8125 10656 8198
rect 12341 8196 12388 8198
rect 12452 8196 12458 8260
rect 12341 8195 12407 8196
rect 10805 8192 11125 8193
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 8127 11125 8128
rect 1577 8122 1643 8125
rect 1534 8120 1643 8122
rect 1534 8064 1582 8120
rect 1638 8064 1643 8120
rect 1534 8059 1643 8064
rect 1761 8120 1827 8125
rect 1761 8064 1766 8120
rect 1822 8064 1827 8120
rect 1761 8059 1827 8064
rect 2681 8122 2747 8125
rect 4429 8122 4495 8125
rect 2681 8120 4495 8122
rect 2681 8064 2686 8120
rect 2742 8064 4434 8120
rect 4490 8064 4495 8120
rect 2681 8062 4495 8064
rect 2681 8059 2747 8062
rect 4429 8059 4495 8062
rect 7465 8122 7531 8125
rect 8937 8122 9003 8125
rect 7465 8120 9003 8122
rect 7465 8064 7470 8120
rect 7526 8064 8942 8120
rect 8998 8064 9003 8120
rect 7465 8062 9003 8064
rect 7465 8059 7531 8062
rect 8937 8059 9003 8062
rect 9489 8122 9555 8125
rect 10409 8122 10475 8125
rect 9489 8120 10475 8122
rect 9489 8064 9494 8120
rect 9550 8064 10414 8120
rect 10470 8064 10475 8120
rect 9489 8062 10475 8064
rect 9489 8059 9555 8062
rect 10409 8059 10475 8062
rect 10593 8120 10659 8125
rect 10593 8064 10598 8120
rect 10654 8064 10659 8120
rect 10593 8059 10659 8064
rect 11973 8122 12039 8125
rect 14038 8122 14044 8124
rect 11973 8120 14044 8122
rect 11973 8064 11978 8120
rect 12034 8064 14044 8120
rect 11973 8062 14044 8064
rect 11973 8059 12039 8062
rect 14038 8060 14044 8062
rect 14108 8060 14114 8124
rect 1534 7989 1594 8059
rect 1764 7989 1824 8059
rect 1534 7984 1643 7989
rect 1534 7928 1582 7984
rect 1638 7928 1643 7984
rect 1534 7926 1643 7928
rect 1577 7923 1643 7926
rect 1761 7984 1827 7989
rect 1761 7928 1766 7984
rect 1822 7928 1827 7984
rect 1761 7923 1827 7928
rect 3509 7986 3575 7989
rect 7966 7986 7972 7988
rect 3509 7984 7972 7986
rect 3509 7928 3514 7984
rect 3570 7928 7972 7984
rect 3509 7926 7972 7928
rect 3509 7923 3575 7926
rect 7966 7924 7972 7926
rect 8036 7924 8042 7988
rect 8150 7924 8156 7988
rect 8220 7986 8226 7988
rect 12341 7986 12407 7989
rect 8220 7984 12407 7986
rect 8220 7928 12346 7984
rect 12402 7928 12407 7984
rect 8220 7926 12407 7928
rect 8220 7924 8226 7926
rect 12341 7923 12407 7926
rect 2129 7850 2195 7853
rect 3417 7850 3483 7853
rect 2129 7848 3483 7850
rect 2129 7792 2134 7848
rect 2190 7792 3422 7848
rect 3478 7792 3483 7848
rect 2129 7790 3483 7792
rect 2129 7787 2195 7790
rect 3417 7787 3483 7790
rect 3693 7850 3759 7853
rect 4245 7850 4311 7853
rect 3693 7848 4311 7850
rect 3693 7792 3698 7848
rect 3754 7792 4250 7848
rect 4306 7792 4311 7848
rect 3693 7790 4311 7792
rect 3693 7787 3759 7790
rect 4245 7787 4311 7790
rect 8201 7850 8267 7853
rect 10593 7850 10659 7853
rect 11145 7850 11211 7853
rect 8201 7848 10472 7850
rect 8201 7792 8206 7848
rect 8262 7792 10472 7848
rect 8201 7790 10472 7792
rect 8201 7787 8267 7790
rect 2773 7714 2839 7717
rect 2957 7714 3023 7717
rect 2773 7712 3023 7714
rect 2773 7656 2778 7712
rect 2834 7656 2962 7712
rect 3018 7656 3023 7712
rect 2773 7654 3023 7656
rect 2773 7651 2839 7654
rect 2957 7651 3023 7654
rect 4613 7714 4679 7717
rect 7833 7714 7899 7717
rect 4613 7712 7899 7714
rect 4613 7656 4618 7712
rect 4674 7656 7838 7712
rect 7894 7656 7899 7712
rect 4613 7654 7899 7656
rect 10412 7714 10472 7790
rect 10593 7848 11211 7850
rect 10593 7792 10598 7848
rect 10654 7792 11150 7848
rect 11206 7792 11211 7848
rect 10593 7790 11211 7792
rect 10593 7787 10659 7790
rect 11145 7787 11211 7790
rect 12014 7788 12020 7852
rect 12084 7850 12090 7852
rect 12249 7850 12315 7853
rect 13854 7850 13860 7852
rect 12084 7848 12315 7850
rect 12084 7792 12254 7848
rect 12310 7792 12315 7848
rect 12084 7790 12315 7792
rect 12084 7788 12090 7790
rect 12249 7787 12315 7790
rect 12390 7790 13860 7850
rect 10593 7714 10659 7717
rect 10412 7712 10659 7714
rect 10412 7656 10598 7712
rect 10654 7656 10659 7712
rect 10412 7654 10659 7656
rect 4613 7651 4679 7654
rect 7833 7651 7899 7654
rect 10593 7651 10659 7654
rect 10777 7714 10843 7717
rect 12390 7714 12450 7790
rect 13854 7788 13860 7790
rect 13924 7788 13930 7852
rect 10777 7712 12450 7714
rect 10777 7656 10782 7712
rect 10838 7656 12450 7712
rect 10777 7654 12450 7656
rect 10777 7651 10843 7654
rect 3409 7648 3729 7649
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 7583 3729 7584
rect 8340 7648 8660 7649
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 7583 8660 7584
rect 13270 7648 13590 7649
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 7583 13590 7584
rect 2497 7578 2563 7581
rect 4613 7578 4679 7581
rect 8201 7578 8267 7581
rect 2497 7576 3250 7578
rect 2497 7520 2502 7576
rect 2558 7520 3250 7576
rect 2497 7518 3250 7520
rect 2497 7515 2563 7518
rect 0 7442 480 7472
rect 3049 7442 3115 7445
rect 0 7440 3115 7442
rect 0 7384 3054 7440
rect 3110 7384 3115 7440
rect 0 7382 3115 7384
rect 3190 7442 3250 7518
rect 4613 7576 8267 7578
rect 4613 7520 4618 7576
rect 4674 7520 8206 7576
rect 8262 7520 8267 7576
rect 4613 7518 8267 7520
rect 4613 7515 4679 7518
rect 8201 7515 8267 7518
rect 9070 7516 9076 7580
rect 9140 7578 9146 7580
rect 9140 7518 13002 7578
rect 9140 7516 9146 7518
rect 12801 7442 12867 7445
rect 3190 7440 12867 7442
rect 3190 7384 12806 7440
rect 12862 7384 12867 7440
rect 3190 7382 12867 7384
rect 12942 7442 13002 7518
rect 13629 7442 13695 7445
rect 12942 7440 13695 7442
rect 12942 7384 13634 7440
rect 13690 7384 13695 7440
rect 12942 7382 13695 7384
rect 0 7352 480 7382
rect 3049 7379 3115 7382
rect 12801 7379 12867 7382
rect 13629 7379 13695 7382
rect 1853 7306 1919 7309
rect 13629 7306 13695 7309
rect 1853 7304 13695 7306
rect 1853 7248 1858 7304
rect 1914 7248 13634 7304
rect 13690 7248 13695 7304
rect 1853 7246 13695 7248
rect 1853 7243 1919 7246
rect 13629 7243 13695 7246
rect 7833 7170 7899 7173
rect 9121 7170 9187 7173
rect 7833 7168 9187 7170
rect 7833 7112 7838 7168
rect 7894 7112 9126 7168
rect 9182 7112 9187 7168
rect 7833 7110 9187 7112
rect 7833 7107 7899 7110
rect 9121 7107 9187 7110
rect 11278 7108 11284 7172
rect 11348 7170 11354 7172
rect 11973 7170 12039 7173
rect 11348 7168 12039 7170
rect 11348 7112 11978 7168
rect 12034 7112 12039 7168
rect 11348 7110 12039 7112
rect 11348 7108 11354 7110
rect 11973 7107 12039 7110
rect 5874 7104 6194 7105
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6194 7104
rect 5874 7039 6194 7040
rect 10805 7104 11125 7105
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 7039 11125 7040
rect 7005 7034 7071 7037
rect 8477 7034 8543 7037
rect 7005 7032 8543 7034
rect 7005 6976 7010 7032
rect 7066 6976 8482 7032
rect 8538 6976 8543 7032
rect 7005 6974 8543 6976
rect 7005 6971 7071 6974
rect 8477 6971 8543 6974
rect 10041 7034 10107 7037
rect 10174 7034 10180 7036
rect 10041 7032 10180 7034
rect 10041 6976 10046 7032
rect 10102 6976 10180 7032
rect 10041 6974 10180 6976
rect 10041 6971 10107 6974
rect 10174 6972 10180 6974
rect 10244 6972 10250 7036
rect 2865 6898 2931 6901
rect 1350 6896 2931 6898
rect 1350 6840 2870 6896
rect 2926 6840 2931 6896
rect 1350 6838 2931 6840
rect 0 6490 480 6520
rect 1350 6490 1410 6838
rect 2865 6835 2931 6838
rect 4429 6898 4495 6901
rect 8661 6898 8727 6901
rect 4429 6896 8727 6898
rect 4429 6840 4434 6896
rect 4490 6840 8666 6896
rect 8722 6840 8727 6896
rect 4429 6838 8727 6840
rect 4429 6835 4495 6838
rect 8661 6835 8727 6838
rect 9673 6898 9739 6901
rect 10133 6898 10199 6901
rect 11605 6898 11671 6901
rect 9673 6896 11671 6898
rect 9673 6840 9678 6896
rect 9734 6840 10138 6896
rect 10194 6840 11610 6896
rect 11666 6840 11671 6896
rect 9673 6838 11671 6840
rect 9673 6835 9739 6838
rect 10133 6835 10199 6838
rect 11605 6835 11671 6838
rect 11830 6836 11836 6900
rect 11900 6898 11906 6900
rect 12249 6898 12315 6901
rect 11900 6896 12315 6898
rect 11900 6840 12254 6896
rect 12310 6840 12315 6896
rect 11900 6838 12315 6840
rect 11900 6836 11906 6838
rect 12249 6835 12315 6838
rect 6269 6762 6335 6765
rect 7833 6762 7899 6765
rect 10225 6762 10291 6765
rect 11605 6762 11671 6765
rect 6269 6760 11671 6762
rect 6269 6704 6274 6760
rect 6330 6704 7838 6760
rect 7894 6704 10230 6760
rect 10286 6704 11610 6760
rect 11666 6704 11671 6760
rect 6269 6702 11671 6704
rect 6269 6699 6335 6702
rect 7833 6699 7899 6702
rect 10225 6699 10291 6702
rect 11605 6699 11671 6702
rect 11973 6762 12039 6765
rect 12382 6762 12388 6764
rect 11973 6760 12388 6762
rect 11973 6704 11978 6760
rect 12034 6704 12388 6760
rect 11973 6702 12388 6704
rect 11973 6699 12039 6702
rect 12382 6700 12388 6702
rect 12452 6700 12458 6764
rect 13813 6762 13879 6765
rect 13126 6760 13879 6762
rect 13126 6704 13818 6760
rect 13874 6704 13879 6760
rect 13126 6702 13879 6704
rect 10317 6626 10383 6629
rect 11605 6626 11671 6629
rect 10317 6624 11671 6626
rect 10317 6568 10322 6624
rect 10378 6568 11610 6624
rect 11666 6568 11671 6624
rect 10317 6566 11671 6568
rect 10317 6563 10383 6566
rect 11605 6563 11671 6566
rect 3409 6560 3729 6561
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 13126 6490 13186 6702
rect 13813 6699 13879 6702
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 0 6430 1410 6490
rect 8848 6430 13186 6490
rect 0 6400 480 6430
rect 5257 6354 5323 6357
rect 8848 6354 8908 6430
rect 5257 6352 8908 6354
rect 5257 6296 5262 6352
rect 5318 6296 8908 6352
rect 5257 6294 8908 6296
rect 9581 6354 9647 6357
rect 13077 6354 13143 6357
rect 9581 6352 13143 6354
rect 9581 6296 9586 6352
rect 9642 6296 13082 6352
rect 13138 6296 13143 6352
rect 9581 6294 13143 6296
rect 5257 6291 5323 6294
rect 9581 6291 9647 6294
rect 13077 6291 13143 6294
rect 2589 6218 2655 6221
rect 13629 6218 13695 6221
rect 2589 6216 13695 6218
rect 2589 6160 2594 6216
rect 2650 6160 13634 6216
rect 13690 6160 13695 6216
rect 2589 6158 13695 6160
rect 2589 6155 2655 6158
rect 13629 6155 13695 6158
rect 8201 6084 8267 6085
rect 8150 6082 8156 6084
rect 8110 6022 8156 6082
rect 8220 6080 8267 6084
rect 8262 6024 8267 6080
rect 8150 6020 8156 6022
rect 8220 6020 8267 6024
rect 8201 6019 8267 6020
rect 9213 6082 9279 6085
rect 10501 6082 10567 6085
rect 9213 6080 10567 6082
rect 9213 6024 9218 6080
rect 9274 6024 10506 6080
rect 10562 6024 10567 6080
rect 9213 6022 10567 6024
rect 9213 6019 9279 6022
rect 10501 6019 10567 6022
rect 11830 6020 11836 6084
rect 11900 6082 11906 6084
rect 12893 6082 12959 6085
rect 11900 6080 12959 6082
rect 11900 6024 12898 6080
rect 12954 6024 12959 6080
rect 11900 6022 12959 6024
rect 11900 6020 11906 6022
rect 12893 6019 12959 6022
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 9673 5946 9739 5949
rect 11329 5946 11395 5949
rect 14917 5946 14983 5949
rect 9673 5944 10656 5946
rect 9673 5888 9678 5944
rect 9734 5888 10656 5944
rect 9673 5886 10656 5888
rect 9673 5883 9739 5886
rect 4521 5810 4587 5813
rect 9581 5810 9647 5813
rect 4521 5808 9647 5810
rect 4521 5752 4526 5808
rect 4582 5752 9586 5808
rect 9642 5752 9647 5808
rect 4521 5750 9647 5752
rect 4521 5747 4587 5750
rect 9581 5747 9647 5750
rect 9857 5810 9923 5813
rect 10596 5810 10656 5886
rect 11329 5944 14983 5946
rect 11329 5888 11334 5944
rect 11390 5888 14922 5944
rect 14978 5888 14983 5944
rect 11329 5886 14983 5888
rect 11329 5883 11395 5886
rect 14917 5883 14983 5886
rect 10961 5810 11027 5813
rect 9857 5808 10426 5810
rect 9857 5752 9862 5808
rect 9918 5752 10426 5808
rect 9857 5750 10426 5752
rect 10596 5808 11027 5810
rect 10596 5752 10966 5808
rect 11022 5752 11027 5808
rect 10596 5750 11027 5752
rect 9857 5747 9923 5750
rect 10041 5674 10107 5677
rect 3880 5672 10107 5674
rect 3880 5616 10046 5672
rect 10102 5616 10107 5672
rect 3880 5614 10107 5616
rect 3880 5541 3940 5614
rect 10041 5611 10107 5614
rect 3877 5536 3943 5541
rect 3877 5480 3882 5536
rect 3938 5480 3943 5536
rect 3877 5475 3943 5480
rect 5073 5538 5139 5541
rect 7833 5538 7899 5541
rect 5073 5536 7899 5538
rect 5073 5480 5078 5536
rect 5134 5480 7838 5536
rect 7894 5480 7899 5536
rect 5073 5478 7899 5480
rect 5073 5475 5139 5478
rect 7833 5475 7899 5478
rect 8886 5476 8892 5540
rect 8956 5538 8962 5540
rect 9305 5538 9371 5541
rect 8956 5536 9371 5538
rect 8956 5480 9310 5536
rect 9366 5480 9371 5536
rect 8956 5478 9371 5480
rect 10366 5538 10426 5750
rect 10961 5747 11027 5750
rect 10501 5674 10567 5677
rect 13118 5674 13124 5676
rect 10501 5672 13124 5674
rect 10501 5616 10506 5672
rect 10562 5616 13124 5672
rect 10501 5614 13124 5616
rect 10501 5611 10567 5614
rect 13118 5612 13124 5614
rect 13188 5612 13194 5676
rect 11329 5538 11395 5541
rect 10366 5536 11395 5538
rect 10366 5480 11334 5536
rect 11390 5480 11395 5536
rect 10366 5478 11395 5480
rect 8956 5476 8962 5478
rect 9305 5475 9371 5478
rect 11329 5475 11395 5478
rect 3409 5472 3729 5473
rect 0 5402 480 5432
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 2957 5402 3023 5405
rect 7741 5402 7807 5405
rect 0 5400 3023 5402
rect 0 5344 2962 5400
rect 3018 5344 3023 5400
rect 0 5342 3023 5344
rect 0 5312 480 5342
rect 2957 5339 3023 5342
rect 4110 5400 7807 5402
rect 4110 5344 7746 5400
rect 7802 5344 7807 5400
rect 4110 5342 7807 5344
rect 3417 5130 3483 5133
rect 4110 5130 4170 5342
rect 7741 5339 7807 5342
rect 8886 5340 8892 5404
rect 8956 5402 8962 5404
rect 9029 5402 9095 5405
rect 8956 5400 9095 5402
rect 8956 5344 9034 5400
rect 9090 5344 9095 5400
rect 8956 5342 9095 5344
rect 8956 5340 8962 5342
rect 9029 5339 9095 5342
rect 9213 5402 9279 5405
rect 10501 5402 10567 5405
rect 9213 5400 10567 5402
rect 9213 5344 9218 5400
rect 9274 5344 10506 5400
rect 10562 5344 10567 5400
rect 9213 5342 10567 5344
rect 9213 5339 9279 5342
rect 10501 5339 10567 5342
rect 4286 5204 4292 5268
rect 4356 5266 4362 5268
rect 13445 5266 13511 5269
rect 4356 5264 13511 5266
rect 4356 5208 13450 5264
rect 13506 5208 13511 5264
rect 4356 5206 13511 5208
rect 4356 5204 4362 5206
rect 13445 5203 13511 5206
rect 3417 5128 4170 5130
rect 3417 5072 3422 5128
rect 3478 5072 4170 5128
rect 3417 5070 4170 5072
rect 4245 5130 4311 5133
rect 11513 5130 11579 5133
rect 13629 5130 13695 5133
rect 14406 5130 14412 5132
rect 4245 5128 11579 5130
rect 4245 5072 4250 5128
rect 4306 5072 11518 5128
rect 11574 5072 11579 5128
rect 4245 5070 11579 5072
rect 3417 5067 3483 5070
rect 4245 5067 4311 5070
rect 11513 5067 11579 5070
rect 11792 5128 14412 5130
rect 11792 5072 13634 5128
rect 13690 5072 14412 5128
rect 11792 5070 14412 5072
rect 11792 4997 11852 5070
rect 13629 5067 13695 5070
rect 14406 5068 14412 5070
rect 14476 5068 14482 5132
rect 9029 4994 9095 4997
rect 11237 4996 11303 4997
rect 10174 4994 10180 4996
rect 6318 4992 9095 4994
rect 6318 4936 9034 4992
rect 9090 4936 9095 4992
rect 6318 4934 9095 4936
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 1853 4722 1919 4725
rect 6318 4722 6378 4934
rect 9029 4931 9095 4934
rect 9262 4934 10180 4994
rect 6637 4858 6703 4861
rect 6821 4858 6887 4861
rect 8477 4858 8543 4861
rect 9262 4858 9322 4934
rect 10174 4932 10180 4934
rect 10244 4932 10250 4996
rect 11237 4992 11284 4996
rect 11348 4994 11354 4996
rect 11237 4936 11242 4992
rect 11237 4932 11284 4936
rect 11348 4934 11394 4994
rect 11789 4992 11855 4997
rect 15193 4994 15259 4997
rect 11789 4936 11794 4992
rect 11850 4936 11855 4992
rect 11348 4932 11354 4934
rect 11237 4931 11303 4932
rect 11789 4931 11855 4936
rect 12206 4992 15259 4994
rect 12206 4936 15198 4992
rect 15254 4936 15259 4992
rect 12206 4934 15259 4936
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 6637 4856 6887 4858
rect 6637 4800 6642 4856
rect 6698 4800 6826 4856
rect 6882 4800 6887 4856
rect 6637 4798 6887 4800
rect 6637 4795 6703 4798
rect 6821 4795 6887 4798
rect 7836 4856 9322 4858
rect 7836 4800 8482 4856
rect 8538 4800 9322 4856
rect 7836 4798 9322 4800
rect 9397 4860 9463 4861
rect 9397 4856 9444 4860
rect 9508 4858 9514 4860
rect 9673 4858 9739 4861
rect 9857 4858 9923 4861
rect 9397 4800 9402 4856
rect 1853 4720 6378 4722
rect 1853 4664 1858 4720
rect 1914 4664 6378 4720
rect 1853 4662 6378 4664
rect 6913 4722 6979 4725
rect 7836 4722 7896 4798
rect 8477 4795 8543 4798
rect 9397 4796 9444 4800
rect 9508 4798 9554 4858
rect 9673 4856 9923 4858
rect 9673 4800 9678 4856
rect 9734 4800 9862 4856
rect 9918 4800 9923 4856
rect 9673 4798 9923 4800
rect 9508 4796 9514 4798
rect 9397 4795 9463 4796
rect 9673 4795 9739 4798
rect 9857 4795 9923 4798
rect 6913 4720 7896 4722
rect 6913 4664 6918 4720
rect 6974 4664 7896 4720
rect 6913 4662 7896 4664
rect 8017 4722 8083 4725
rect 12206 4722 12266 4934
rect 15193 4931 15259 4934
rect 12341 4858 12407 4861
rect 14089 4858 14155 4861
rect 12341 4856 14155 4858
rect 12341 4800 12346 4856
rect 12402 4800 14094 4856
rect 14150 4800 14155 4856
rect 12341 4798 14155 4800
rect 12341 4795 12407 4798
rect 14089 4795 14155 4798
rect 8017 4720 12266 4722
rect 8017 4664 8022 4720
rect 8078 4664 12266 4720
rect 8017 4662 12266 4664
rect 1853 4659 1919 4662
rect 6913 4659 6979 4662
rect 8017 4659 8083 4662
rect 2129 4586 2195 4589
rect 14641 4586 14707 4589
rect 2129 4584 14707 4586
rect 2129 4528 2134 4584
rect 2190 4528 14646 4584
rect 14702 4528 14707 4584
rect 2129 4526 14707 4528
rect 2129 4523 2195 4526
rect 14641 4523 14707 4526
rect 0 4450 480 4480
rect 2957 4450 3023 4453
rect 0 4448 3023 4450
rect 0 4392 2962 4448
rect 3018 4392 3023 4448
rect 0 4390 3023 4392
rect 0 4360 480 4390
rect 2957 4387 3023 4390
rect 4613 4450 4679 4453
rect 7465 4450 7531 4453
rect 4613 4448 7531 4450
rect 4613 4392 4618 4448
rect 4674 4392 7470 4448
rect 7526 4392 7531 4448
rect 4613 4390 7531 4392
rect 4613 4387 4679 4390
rect 7465 4387 7531 4390
rect 9121 4450 9187 4453
rect 11830 4450 11836 4452
rect 9121 4448 11836 4450
rect 9121 4392 9126 4448
rect 9182 4392 11836 4448
rect 9121 4390 11836 4392
rect 9121 4387 9187 4390
rect 11830 4388 11836 4390
rect 11900 4388 11906 4452
rect 3409 4384 3729 4385
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 4319 13590 4320
rect 4337 4314 4403 4317
rect 4981 4314 5047 4317
rect 4337 4312 5047 4314
rect 4337 4256 4342 4312
rect 4398 4256 4986 4312
rect 5042 4256 5047 4312
rect 4337 4254 5047 4256
rect 4337 4251 4403 4254
rect 4981 4251 5047 4254
rect 5349 4314 5415 4317
rect 7741 4314 7807 4317
rect 9622 4314 9628 4316
rect 5349 4312 8264 4314
rect 5349 4256 5354 4312
rect 5410 4256 7746 4312
rect 7802 4256 8264 4312
rect 5349 4254 8264 4256
rect 5349 4251 5415 4254
rect 7741 4251 7807 4254
rect 5073 4178 5139 4181
rect 7557 4178 7623 4181
rect 5073 4176 7623 4178
rect 5073 4120 5078 4176
rect 5134 4120 7562 4176
rect 7618 4120 7623 4176
rect 5073 4118 7623 4120
rect 8204 4178 8264 4254
rect 8848 4254 9628 4314
rect 8848 4178 8908 4254
rect 9622 4252 9628 4254
rect 9692 4314 9698 4316
rect 11329 4314 11395 4317
rect 9692 4312 11395 4314
rect 9692 4256 11334 4312
rect 11390 4256 11395 4312
rect 9692 4254 11395 4256
rect 9692 4252 9698 4254
rect 11329 4251 11395 4254
rect 8204 4118 8908 4178
rect 9581 4178 9647 4181
rect 12157 4178 12223 4181
rect 12750 4178 12756 4180
rect 9581 4176 12756 4178
rect 9581 4120 9586 4176
rect 9642 4120 12162 4176
rect 12218 4120 12756 4176
rect 9581 4118 12756 4120
rect 5073 4115 5139 4118
rect 7557 4115 7623 4118
rect 9581 4115 9647 4118
rect 12157 4115 12223 4118
rect 12750 4116 12756 4118
rect 12820 4116 12826 4180
rect 12934 4116 12940 4180
rect 13004 4178 13010 4180
rect 13261 4178 13327 4181
rect 14917 4178 14983 4181
rect 13004 4176 14983 4178
rect 13004 4120 13266 4176
rect 13322 4120 14922 4176
rect 14978 4120 14983 4176
rect 13004 4118 14983 4120
rect 13004 4116 13010 4118
rect 13261 4115 13327 4118
rect 14917 4115 14983 4118
rect 2497 4042 2563 4045
rect 16757 4042 16823 4045
rect 2497 4040 16823 4042
rect 2497 3984 2502 4040
rect 2558 3984 16762 4040
rect 16818 3984 16823 4040
rect 2497 3982 16823 3984
rect 2497 3979 2563 3982
rect 16757 3979 16823 3982
rect 7925 3906 7991 3909
rect 10041 3906 10107 3909
rect 7925 3904 10107 3906
rect 7925 3848 7930 3904
rect 7986 3848 10046 3904
rect 10102 3848 10107 3904
rect 7925 3846 10107 3848
rect 7925 3843 7991 3846
rect 10041 3843 10107 3846
rect 10225 3906 10291 3909
rect 10358 3906 10364 3908
rect 10225 3904 10364 3906
rect 10225 3848 10230 3904
rect 10286 3848 10364 3904
rect 10225 3846 10364 3848
rect 10225 3843 10291 3846
rect 10358 3844 10364 3846
rect 10428 3844 10434 3908
rect 11421 3906 11487 3909
rect 11646 3906 11652 3908
rect 11421 3904 11652 3906
rect 11421 3848 11426 3904
rect 11482 3848 11652 3904
rect 11421 3846 11652 3848
rect 11421 3843 11487 3846
rect 11646 3844 11652 3846
rect 11716 3844 11722 3908
rect 12157 3906 12223 3909
rect 13629 3906 13695 3909
rect 14089 3908 14155 3909
rect 14038 3906 14044 3908
rect 12157 3904 14044 3906
rect 14108 3906 14155 3908
rect 14108 3904 14236 3906
rect 12157 3848 12162 3904
rect 12218 3848 13634 3904
rect 13690 3848 14044 3904
rect 14150 3848 14236 3904
rect 12157 3846 14044 3848
rect 12157 3843 12223 3846
rect 13629 3843 13695 3846
rect 14038 3844 14044 3846
rect 14108 3846 14236 3848
rect 14108 3844 14155 3846
rect 14089 3843 14155 3844
rect 5874 3840 6194 3841
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 7557 3770 7623 3773
rect 10225 3770 10291 3773
rect 10409 3770 10475 3773
rect 14641 3770 14707 3773
rect 7557 3768 10475 3770
rect 7557 3712 7562 3768
rect 7618 3712 10230 3768
rect 10286 3712 10414 3768
rect 10470 3712 10475 3768
rect 7557 3710 10475 3712
rect 7557 3707 7623 3710
rect 10225 3707 10291 3710
rect 10409 3707 10475 3710
rect 11286 3768 14707 3770
rect 11286 3712 14646 3768
rect 14702 3712 14707 3768
rect 11286 3710 14707 3712
rect 1761 3634 1827 3637
rect 11286 3634 11346 3710
rect 14641 3707 14707 3710
rect 1761 3632 11346 3634
rect 1761 3576 1766 3632
rect 1822 3576 11346 3632
rect 1761 3574 11346 3576
rect 1761 3571 1827 3574
rect 0 3498 480 3528
rect 2589 3498 2655 3501
rect 12617 3498 12683 3501
rect 0 3496 2655 3498
rect 0 3440 2594 3496
rect 2650 3440 2655 3496
rect 0 3438 2655 3440
rect 0 3408 480 3438
rect 2589 3435 2655 3438
rect 2776 3438 9736 3498
rect 1485 3226 1551 3229
rect 2776 3226 2836 3438
rect 9676 3365 9736 3438
rect 9952 3496 12683 3498
rect 9952 3440 12622 3496
rect 12678 3440 12683 3496
rect 9952 3438 12683 3440
rect 8845 3364 8911 3365
rect 8845 3362 8892 3364
rect 8800 3360 8892 3362
rect 8800 3304 8850 3360
rect 8800 3302 8892 3304
rect 8845 3300 8892 3302
rect 8956 3300 8962 3364
rect 9029 3362 9095 3365
rect 9489 3362 9555 3365
rect 9029 3360 9555 3362
rect 9029 3304 9034 3360
rect 9090 3304 9494 3360
rect 9550 3304 9555 3360
rect 9029 3302 9555 3304
rect 8845 3299 8911 3300
rect 9029 3299 9095 3302
rect 9489 3299 9555 3302
rect 9673 3360 9739 3365
rect 9673 3304 9678 3360
rect 9734 3304 9739 3360
rect 9673 3299 9739 3304
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 1485 3224 2836 3226
rect 1485 3168 1490 3224
rect 1546 3168 2836 3224
rect 1485 3166 2836 3168
rect 4429 3226 4495 3229
rect 5625 3226 5691 3229
rect 8201 3228 8267 3229
rect 8150 3226 8156 3228
rect 4429 3224 5691 3226
rect 4429 3168 4434 3224
rect 4490 3168 5630 3224
rect 5686 3168 5691 3224
rect 4429 3166 5691 3168
rect 8110 3166 8156 3226
rect 8220 3224 8267 3228
rect 9952 3226 10012 3438
rect 12617 3435 12683 3438
rect 13261 3498 13327 3501
rect 14089 3498 14155 3501
rect 13261 3496 14155 3498
rect 13261 3440 13266 3496
rect 13322 3440 14094 3496
rect 14150 3440 14155 3496
rect 13261 3438 14155 3440
rect 13261 3435 13327 3438
rect 14089 3435 14155 3438
rect 10542 3300 10548 3364
rect 10612 3362 10618 3364
rect 10777 3362 10843 3365
rect 12617 3364 12683 3365
rect 10612 3360 10843 3362
rect 10612 3304 10782 3360
rect 10838 3304 10843 3360
rect 10612 3302 10843 3304
rect 10612 3300 10618 3302
rect 10777 3299 10843 3302
rect 12566 3300 12572 3364
rect 12636 3362 12683 3364
rect 15561 3362 15627 3365
rect 16520 3362 17000 3392
rect 12636 3360 12728 3362
rect 12678 3304 12728 3360
rect 12636 3302 12728 3304
rect 15561 3360 17000 3362
rect 15561 3304 15566 3360
rect 15622 3304 17000 3360
rect 15561 3302 17000 3304
rect 12636 3300 12683 3302
rect 12617 3299 12683 3300
rect 15561 3299 15627 3302
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 16520 3272 17000 3302
rect 13270 3231 13590 3232
rect 8262 3168 8267 3224
rect 1485 3163 1551 3166
rect 4429 3163 4495 3166
rect 5625 3163 5691 3166
rect 8150 3164 8156 3166
rect 8220 3164 8267 3168
rect 8201 3163 8267 3164
rect 8848 3166 10012 3226
rect 2773 3090 2839 3093
rect 8848 3090 8908 3166
rect 10174 3164 10180 3228
rect 10244 3226 10250 3228
rect 10777 3226 10843 3229
rect 10244 3224 10843 3226
rect 10244 3168 10782 3224
rect 10838 3168 10843 3224
rect 10244 3166 10843 3168
rect 10244 3164 10250 3166
rect 10777 3163 10843 3166
rect 12206 3166 13186 3226
rect 9765 3092 9831 3093
rect 9765 3090 9812 3092
rect 2773 3088 8908 3090
rect 2773 3032 2778 3088
rect 2834 3032 8908 3088
rect 2773 3030 8908 3032
rect 9720 3088 9812 3090
rect 9720 3032 9770 3088
rect 9720 3030 9812 3032
rect 2773 3027 2839 3030
rect 9765 3028 9812 3030
rect 9876 3028 9882 3092
rect 11237 3090 11303 3093
rect 11421 3090 11487 3093
rect 12206 3092 12266 3166
rect 12893 3092 12959 3093
rect 12198 3090 12204 3092
rect 11237 3088 12204 3090
rect 11237 3032 11242 3088
rect 11298 3032 11426 3088
rect 11482 3032 12204 3088
rect 11237 3030 12204 3032
rect 9765 3027 9831 3028
rect 11237 3027 11303 3030
rect 11421 3027 11487 3030
rect 12198 3028 12204 3030
rect 12268 3028 12274 3092
rect 12893 3088 12940 3092
rect 13004 3090 13010 3092
rect 13126 3090 13186 3166
rect 14457 3090 14523 3093
rect 12893 3032 12898 3088
rect 12893 3028 12940 3032
rect 13004 3030 13050 3090
rect 13126 3088 14523 3090
rect 13126 3032 14462 3088
rect 14518 3032 14523 3088
rect 13126 3030 14523 3032
rect 13004 3028 13010 3030
rect 12893 3027 12959 3028
rect 14457 3027 14523 3030
rect 1117 2954 1183 2957
rect 14089 2954 14155 2957
rect 1117 2952 14155 2954
rect 1117 2896 1122 2952
rect 1178 2896 14094 2952
rect 14150 2896 14155 2952
rect 1117 2894 14155 2896
rect 1117 2891 1183 2894
rect 14089 2891 14155 2894
rect 4613 2818 4679 2821
rect 4981 2818 5047 2821
rect 4613 2816 5047 2818
rect 4613 2760 4618 2816
rect 4674 2760 4986 2816
rect 5042 2760 5047 2816
rect 4613 2758 5047 2760
rect 4613 2755 4679 2758
rect 4981 2755 5047 2758
rect 7005 2818 7071 2821
rect 10041 2818 10107 2821
rect 7005 2816 10107 2818
rect 7005 2760 7010 2816
rect 7066 2760 10046 2816
rect 10102 2760 10107 2816
rect 7005 2758 10107 2760
rect 7005 2755 7071 2758
rect 10041 2755 10107 2758
rect 13629 2820 13695 2821
rect 13629 2816 13676 2820
rect 13740 2818 13746 2820
rect 13629 2760 13634 2816
rect 13629 2756 13676 2760
rect 13740 2758 13786 2818
rect 13740 2756 13746 2758
rect 13629 2755 13695 2756
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 9213 2682 9279 2685
rect 9949 2684 10015 2685
rect 11421 2684 11487 2685
rect 9438 2682 9444 2684
rect 9213 2680 9444 2682
rect 9213 2624 9218 2680
rect 9274 2624 9444 2680
rect 9213 2622 9444 2624
rect 9213 2619 9279 2622
rect 9438 2620 9444 2622
rect 9508 2620 9514 2684
rect 9949 2682 9996 2684
rect 9904 2680 9996 2682
rect 9904 2624 9954 2680
rect 9904 2622 9996 2624
rect 9949 2620 9996 2622
rect 10060 2620 10066 2684
rect 11421 2680 11468 2684
rect 11532 2682 11538 2684
rect 11421 2624 11426 2680
rect 11421 2620 11468 2624
rect 11532 2622 11578 2682
rect 11532 2620 11538 2622
rect 9949 2619 10015 2620
rect 11421 2619 11487 2620
rect 3049 2546 3115 2549
rect 4470 2546 4476 2548
rect 3049 2544 4476 2546
rect 3049 2488 3054 2544
rect 3110 2488 4476 2544
rect 3049 2486 4476 2488
rect 3049 2483 3115 2486
rect 4470 2484 4476 2486
rect 4540 2546 4546 2548
rect 7557 2546 7623 2549
rect 4540 2544 7623 2546
rect 4540 2488 7562 2544
rect 7618 2488 7623 2544
rect 4540 2486 7623 2488
rect 4540 2484 4546 2486
rect 7557 2483 7623 2486
rect 8569 2546 8635 2549
rect 12893 2548 12959 2549
rect 9254 2546 9260 2548
rect 8569 2544 9260 2546
rect 8569 2488 8574 2544
rect 8630 2488 9260 2544
rect 8569 2486 9260 2488
rect 8569 2483 8635 2486
rect 9254 2484 9260 2486
rect 9324 2546 9330 2548
rect 12893 2546 12940 2548
rect 9324 2544 12940 2546
rect 13004 2546 13010 2548
rect 9324 2488 12898 2544
rect 9324 2486 12940 2488
rect 9324 2484 9330 2486
rect 12893 2484 12940 2486
rect 13004 2486 13086 2546
rect 13004 2484 13010 2486
rect 12893 2483 12959 2484
rect 0 2410 480 2440
rect 8661 2410 8727 2413
rect 0 2408 8727 2410
rect 0 2352 8666 2408
rect 8722 2352 8727 2408
rect 0 2350 8727 2352
rect 0 2320 480 2350
rect 8661 2347 8727 2350
rect 8845 2410 8911 2413
rect 12433 2410 12499 2413
rect 8845 2408 12499 2410
rect 8845 2352 8850 2408
rect 8906 2352 12438 2408
rect 12494 2352 12499 2408
rect 8845 2350 12499 2352
rect 8845 2347 8911 2350
rect 12433 2347 12499 2350
rect 10961 2274 11027 2277
rect 12014 2274 12020 2276
rect 10961 2272 12020 2274
rect 10961 2216 10966 2272
rect 11022 2216 12020 2272
rect 10961 2214 12020 2216
rect 10961 2211 11027 2214
rect 12014 2212 12020 2214
rect 12084 2212 12090 2276
rect 3409 2208 3729 2209
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
rect 9029 2138 9095 2141
rect 11789 2138 11855 2141
rect 9029 2136 11855 2138
rect 9029 2080 9034 2136
rect 9090 2080 11794 2136
rect 11850 2080 11855 2136
rect 9029 2078 11855 2080
rect 9029 2075 9095 2078
rect 11789 2075 11855 2078
rect 4153 2002 4219 2005
rect 9070 2002 9076 2004
rect 4153 2000 9076 2002
rect 4153 1944 4158 2000
rect 4214 1944 9076 2000
rect 4153 1942 9076 1944
rect 4153 1939 4219 1942
rect 9070 1940 9076 1942
rect 9140 1940 9146 2004
rect 0 1458 480 1488
rect 2037 1458 2103 1461
rect 0 1456 2103 1458
rect 0 1400 2042 1456
rect 2098 1400 2103 1456
rect 0 1398 2103 1400
rect 0 1368 480 1398
rect 2037 1395 2103 1398
rect 0 506 480 536
rect 2865 506 2931 509
rect 0 504 2931 506
rect 0 448 2870 504
rect 2926 448 2931 504
rect 0 446 2931 448
rect 0 416 480 446
rect 2865 443 2931 446
<< via3 >>
rect 13124 17580 13188 17644
rect 3417 17436 3481 17440
rect 3417 17380 3421 17436
rect 3421 17380 3477 17436
rect 3477 17380 3481 17436
rect 3417 17376 3481 17380
rect 3497 17436 3561 17440
rect 3497 17380 3501 17436
rect 3501 17380 3557 17436
rect 3557 17380 3561 17436
rect 3497 17376 3561 17380
rect 3577 17436 3641 17440
rect 3577 17380 3581 17436
rect 3581 17380 3637 17436
rect 3637 17380 3641 17436
rect 3577 17376 3641 17380
rect 3657 17436 3721 17440
rect 3657 17380 3661 17436
rect 3661 17380 3717 17436
rect 3717 17380 3721 17436
rect 3657 17376 3721 17380
rect 8348 17436 8412 17440
rect 8348 17380 8352 17436
rect 8352 17380 8408 17436
rect 8408 17380 8412 17436
rect 8348 17376 8412 17380
rect 8428 17436 8492 17440
rect 8428 17380 8432 17436
rect 8432 17380 8488 17436
rect 8488 17380 8492 17436
rect 8428 17376 8492 17380
rect 8508 17436 8572 17440
rect 8508 17380 8512 17436
rect 8512 17380 8568 17436
rect 8568 17380 8572 17436
rect 8508 17376 8572 17380
rect 8588 17436 8652 17440
rect 8588 17380 8592 17436
rect 8592 17380 8648 17436
rect 8648 17380 8652 17436
rect 8588 17376 8652 17380
rect 13278 17436 13342 17440
rect 13278 17380 13282 17436
rect 13282 17380 13338 17436
rect 13338 17380 13342 17436
rect 13278 17376 13342 17380
rect 13358 17436 13422 17440
rect 13358 17380 13362 17436
rect 13362 17380 13418 17436
rect 13418 17380 13422 17436
rect 13358 17376 13422 17380
rect 13438 17436 13502 17440
rect 13438 17380 13442 17436
rect 13442 17380 13498 17436
rect 13498 17380 13502 17436
rect 13438 17376 13502 17380
rect 13518 17436 13582 17440
rect 13518 17380 13522 17436
rect 13522 17380 13578 17436
rect 13578 17380 13582 17436
rect 13518 17376 13582 17380
rect 9812 17172 9876 17236
rect 11284 17036 11348 17100
rect 5882 16892 5946 16896
rect 5882 16836 5886 16892
rect 5886 16836 5942 16892
rect 5942 16836 5946 16892
rect 5882 16832 5946 16836
rect 5962 16892 6026 16896
rect 5962 16836 5966 16892
rect 5966 16836 6022 16892
rect 6022 16836 6026 16892
rect 5962 16832 6026 16836
rect 6042 16892 6106 16896
rect 6042 16836 6046 16892
rect 6046 16836 6102 16892
rect 6102 16836 6106 16892
rect 6042 16832 6106 16836
rect 6122 16892 6186 16896
rect 6122 16836 6126 16892
rect 6126 16836 6182 16892
rect 6182 16836 6186 16892
rect 6122 16832 6186 16836
rect 10813 16892 10877 16896
rect 10813 16836 10817 16892
rect 10817 16836 10873 16892
rect 10873 16836 10877 16892
rect 10813 16832 10877 16836
rect 10893 16892 10957 16896
rect 10893 16836 10897 16892
rect 10897 16836 10953 16892
rect 10953 16836 10957 16892
rect 10893 16832 10957 16836
rect 10973 16892 11037 16896
rect 10973 16836 10977 16892
rect 10977 16836 11033 16892
rect 11033 16836 11037 16892
rect 10973 16832 11037 16836
rect 11053 16892 11117 16896
rect 11053 16836 11057 16892
rect 11057 16836 11113 16892
rect 11113 16836 11117 16892
rect 11053 16832 11117 16836
rect 4292 16764 4356 16828
rect 9996 16764 10060 16828
rect 14044 16764 14108 16828
rect 13860 16688 13924 16692
rect 13860 16632 13910 16688
rect 13910 16632 13924 16688
rect 13860 16628 13924 16632
rect 13676 16492 13740 16556
rect 3417 16348 3481 16352
rect 3417 16292 3421 16348
rect 3421 16292 3477 16348
rect 3477 16292 3481 16348
rect 3417 16288 3481 16292
rect 3497 16348 3561 16352
rect 3497 16292 3501 16348
rect 3501 16292 3557 16348
rect 3557 16292 3561 16348
rect 3497 16288 3561 16292
rect 3577 16348 3641 16352
rect 3577 16292 3581 16348
rect 3581 16292 3637 16348
rect 3637 16292 3641 16348
rect 3577 16288 3641 16292
rect 3657 16348 3721 16352
rect 3657 16292 3661 16348
rect 3661 16292 3717 16348
rect 3717 16292 3721 16348
rect 3657 16288 3721 16292
rect 8348 16348 8412 16352
rect 8348 16292 8352 16348
rect 8352 16292 8408 16348
rect 8408 16292 8412 16348
rect 8348 16288 8412 16292
rect 8428 16348 8492 16352
rect 8428 16292 8432 16348
rect 8432 16292 8488 16348
rect 8488 16292 8492 16348
rect 8428 16288 8492 16292
rect 8508 16348 8572 16352
rect 8508 16292 8512 16348
rect 8512 16292 8568 16348
rect 8568 16292 8572 16348
rect 8508 16288 8572 16292
rect 8588 16348 8652 16352
rect 8588 16292 8592 16348
rect 8592 16292 8648 16348
rect 8648 16292 8652 16348
rect 8588 16288 8652 16292
rect 13278 16348 13342 16352
rect 13278 16292 13282 16348
rect 13282 16292 13338 16348
rect 13338 16292 13342 16348
rect 13278 16288 13342 16292
rect 13358 16348 13422 16352
rect 13358 16292 13362 16348
rect 13362 16292 13418 16348
rect 13418 16292 13422 16348
rect 13358 16288 13422 16292
rect 13438 16348 13502 16352
rect 13438 16292 13442 16348
rect 13442 16292 13498 16348
rect 13498 16292 13502 16348
rect 13438 16288 13502 16292
rect 13518 16348 13582 16352
rect 13518 16292 13522 16348
rect 13522 16292 13578 16348
rect 13578 16292 13582 16348
rect 13518 16288 13582 16292
rect 7972 16220 8036 16284
rect 9260 16220 9324 16284
rect 9996 16220 10060 16284
rect 8156 16084 8220 16148
rect 5882 15804 5946 15808
rect 5882 15748 5886 15804
rect 5886 15748 5942 15804
rect 5942 15748 5946 15804
rect 5882 15744 5946 15748
rect 5962 15804 6026 15808
rect 5962 15748 5966 15804
rect 5966 15748 6022 15804
rect 6022 15748 6026 15804
rect 5962 15744 6026 15748
rect 6042 15804 6106 15808
rect 6042 15748 6046 15804
rect 6046 15748 6102 15804
rect 6102 15748 6106 15804
rect 6042 15744 6106 15748
rect 6122 15804 6186 15808
rect 6122 15748 6126 15804
rect 6126 15748 6182 15804
rect 6182 15748 6186 15804
rect 6122 15744 6186 15748
rect 10813 15804 10877 15808
rect 10813 15748 10817 15804
rect 10817 15748 10873 15804
rect 10873 15748 10877 15804
rect 10813 15744 10877 15748
rect 10893 15804 10957 15808
rect 10893 15748 10897 15804
rect 10897 15748 10953 15804
rect 10953 15748 10957 15804
rect 10893 15744 10957 15748
rect 10973 15804 11037 15808
rect 10973 15748 10977 15804
rect 10977 15748 11033 15804
rect 11033 15748 11037 15804
rect 10973 15744 11037 15748
rect 11053 15804 11117 15808
rect 11053 15748 11057 15804
rect 11057 15748 11113 15804
rect 11113 15748 11117 15804
rect 11053 15744 11117 15748
rect 8156 15736 8220 15740
rect 8156 15680 8170 15736
rect 8170 15680 8220 15736
rect 8156 15676 8220 15680
rect 9628 15676 9692 15740
rect 9996 15676 10060 15740
rect 3417 15260 3481 15264
rect 3417 15204 3421 15260
rect 3421 15204 3477 15260
rect 3477 15204 3481 15260
rect 3417 15200 3481 15204
rect 3497 15260 3561 15264
rect 3497 15204 3501 15260
rect 3501 15204 3557 15260
rect 3557 15204 3561 15260
rect 3497 15200 3561 15204
rect 3577 15260 3641 15264
rect 3577 15204 3581 15260
rect 3581 15204 3637 15260
rect 3637 15204 3641 15260
rect 3577 15200 3641 15204
rect 3657 15260 3721 15264
rect 3657 15204 3661 15260
rect 3661 15204 3717 15260
rect 3717 15204 3721 15260
rect 3657 15200 3721 15204
rect 8348 15260 8412 15264
rect 8348 15204 8352 15260
rect 8352 15204 8408 15260
rect 8408 15204 8412 15260
rect 8348 15200 8412 15204
rect 8428 15260 8492 15264
rect 8428 15204 8432 15260
rect 8432 15204 8488 15260
rect 8488 15204 8492 15260
rect 8428 15200 8492 15204
rect 8508 15260 8572 15264
rect 8508 15204 8512 15260
rect 8512 15204 8568 15260
rect 8568 15204 8572 15260
rect 8508 15200 8572 15204
rect 8588 15260 8652 15264
rect 8588 15204 8592 15260
rect 8592 15204 8648 15260
rect 8648 15204 8652 15260
rect 8588 15200 8652 15204
rect 11836 15268 11900 15332
rect 13278 15260 13342 15264
rect 13278 15204 13282 15260
rect 13282 15204 13338 15260
rect 13338 15204 13342 15260
rect 13278 15200 13342 15204
rect 13358 15260 13422 15264
rect 13358 15204 13362 15260
rect 13362 15204 13418 15260
rect 13418 15204 13422 15260
rect 13358 15200 13422 15204
rect 13438 15260 13502 15264
rect 13438 15204 13442 15260
rect 13442 15204 13498 15260
rect 13498 15204 13502 15260
rect 13438 15200 13502 15204
rect 13518 15260 13582 15264
rect 13518 15204 13522 15260
rect 13522 15204 13578 15260
rect 13578 15204 13582 15260
rect 13518 15200 13582 15204
rect 13676 14860 13740 14924
rect 7972 14724 8036 14788
rect 10548 14724 10612 14788
rect 12940 14724 13004 14788
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 6122 14716 6186 14720
rect 6122 14660 6126 14716
rect 6126 14660 6182 14716
rect 6182 14660 6186 14716
rect 6122 14656 6186 14660
rect 10813 14716 10877 14720
rect 10813 14660 10817 14716
rect 10817 14660 10873 14716
rect 10873 14660 10877 14716
rect 10813 14656 10877 14660
rect 10893 14716 10957 14720
rect 10893 14660 10897 14716
rect 10897 14660 10953 14716
rect 10953 14660 10957 14716
rect 10893 14656 10957 14660
rect 10973 14716 11037 14720
rect 10973 14660 10977 14716
rect 10977 14660 11033 14716
rect 11033 14660 11037 14716
rect 10973 14656 11037 14660
rect 11053 14716 11117 14720
rect 11053 14660 11057 14716
rect 11057 14660 11113 14716
rect 11113 14660 11117 14716
rect 11053 14656 11117 14660
rect 11284 14452 11348 14516
rect 12204 14452 12268 14516
rect 11652 14316 11716 14380
rect 11468 14180 11532 14244
rect 3417 14172 3481 14176
rect 3417 14116 3421 14172
rect 3421 14116 3477 14172
rect 3477 14116 3481 14172
rect 3417 14112 3481 14116
rect 3497 14172 3561 14176
rect 3497 14116 3501 14172
rect 3501 14116 3557 14172
rect 3557 14116 3561 14172
rect 3497 14112 3561 14116
rect 3577 14172 3641 14176
rect 3577 14116 3581 14172
rect 3581 14116 3637 14172
rect 3637 14116 3641 14172
rect 3577 14112 3641 14116
rect 3657 14172 3721 14176
rect 3657 14116 3661 14172
rect 3661 14116 3717 14172
rect 3717 14116 3721 14172
rect 3657 14112 3721 14116
rect 8348 14172 8412 14176
rect 8348 14116 8352 14172
rect 8352 14116 8408 14172
rect 8408 14116 8412 14172
rect 8348 14112 8412 14116
rect 8428 14172 8492 14176
rect 8428 14116 8432 14172
rect 8432 14116 8488 14172
rect 8488 14116 8492 14172
rect 8428 14112 8492 14116
rect 8508 14172 8572 14176
rect 8508 14116 8512 14172
rect 8512 14116 8568 14172
rect 8568 14116 8572 14172
rect 8508 14112 8572 14116
rect 8588 14172 8652 14176
rect 8588 14116 8592 14172
rect 8592 14116 8648 14172
rect 8648 14116 8652 14172
rect 8588 14112 8652 14116
rect 13278 14172 13342 14176
rect 13278 14116 13282 14172
rect 13282 14116 13338 14172
rect 13338 14116 13342 14172
rect 13278 14112 13342 14116
rect 13358 14172 13422 14176
rect 13358 14116 13362 14172
rect 13362 14116 13418 14172
rect 13418 14116 13422 14172
rect 13358 14112 13422 14116
rect 13438 14172 13502 14176
rect 13438 14116 13442 14172
rect 13442 14116 13498 14172
rect 13498 14116 13502 14172
rect 13438 14112 13502 14116
rect 13518 14172 13582 14176
rect 13518 14116 13522 14172
rect 13522 14116 13578 14172
rect 13578 14116 13582 14172
rect 13518 14112 13582 14116
rect 9444 14044 9508 14108
rect 12388 13908 12452 13972
rect 9076 13772 9140 13836
rect 10364 13772 10428 13836
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 6122 13628 6186 13632
rect 6122 13572 6126 13628
rect 6126 13572 6182 13628
rect 6182 13572 6186 13628
rect 6122 13568 6186 13572
rect 10813 13628 10877 13632
rect 10813 13572 10817 13628
rect 10817 13572 10873 13628
rect 10873 13572 10877 13628
rect 10813 13568 10877 13572
rect 10893 13628 10957 13632
rect 10893 13572 10897 13628
rect 10897 13572 10953 13628
rect 10953 13572 10957 13628
rect 10893 13568 10957 13572
rect 10973 13628 11037 13632
rect 10973 13572 10977 13628
rect 10977 13572 11033 13628
rect 11033 13572 11037 13628
rect 10973 13568 11037 13572
rect 11053 13628 11117 13632
rect 11053 13572 11057 13628
rect 11057 13572 11113 13628
rect 11113 13572 11117 13628
rect 11053 13568 11117 13572
rect 13124 13228 13188 13292
rect 8892 13092 8956 13156
rect 3417 13084 3481 13088
rect 3417 13028 3421 13084
rect 3421 13028 3477 13084
rect 3477 13028 3481 13084
rect 3417 13024 3481 13028
rect 3497 13084 3561 13088
rect 3497 13028 3501 13084
rect 3501 13028 3557 13084
rect 3557 13028 3561 13084
rect 3497 13024 3561 13028
rect 3577 13084 3641 13088
rect 3577 13028 3581 13084
rect 3581 13028 3637 13084
rect 3637 13028 3641 13084
rect 3577 13024 3641 13028
rect 3657 13084 3721 13088
rect 3657 13028 3661 13084
rect 3661 13028 3717 13084
rect 3717 13028 3721 13084
rect 3657 13024 3721 13028
rect 8348 13084 8412 13088
rect 8348 13028 8352 13084
rect 8352 13028 8408 13084
rect 8408 13028 8412 13084
rect 8348 13024 8412 13028
rect 8428 13084 8492 13088
rect 8428 13028 8432 13084
rect 8432 13028 8488 13084
rect 8488 13028 8492 13084
rect 8428 13024 8492 13028
rect 8508 13084 8572 13088
rect 8508 13028 8512 13084
rect 8512 13028 8568 13084
rect 8568 13028 8572 13084
rect 8508 13024 8572 13028
rect 8588 13084 8652 13088
rect 8588 13028 8592 13084
rect 8592 13028 8648 13084
rect 8648 13028 8652 13084
rect 8588 13024 8652 13028
rect 9260 12956 9324 13020
rect 13278 13084 13342 13088
rect 13278 13028 13282 13084
rect 13282 13028 13338 13084
rect 13338 13028 13342 13084
rect 13278 13024 13342 13028
rect 13358 13084 13422 13088
rect 13358 13028 13362 13084
rect 13362 13028 13418 13084
rect 13418 13028 13422 13084
rect 13358 13024 13422 13028
rect 13438 13084 13502 13088
rect 13438 13028 13442 13084
rect 13442 13028 13498 13084
rect 13498 13028 13502 13084
rect 13438 13024 13502 13028
rect 13518 13084 13582 13088
rect 13518 13028 13522 13084
rect 13522 13028 13578 13084
rect 13578 13028 13582 13084
rect 13518 13024 13582 13028
rect 11284 12956 11348 13020
rect 10180 12684 10244 12748
rect 11468 12684 11532 12748
rect 14044 12684 14108 12748
rect 8892 12548 8956 12612
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 6122 12540 6186 12544
rect 6122 12484 6126 12540
rect 6126 12484 6182 12540
rect 6182 12484 6186 12540
rect 6122 12480 6186 12484
rect 11468 12548 11532 12612
rect 10813 12540 10877 12544
rect 10813 12484 10817 12540
rect 10817 12484 10873 12540
rect 10873 12484 10877 12540
rect 10813 12480 10877 12484
rect 10893 12540 10957 12544
rect 10893 12484 10897 12540
rect 10897 12484 10953 12540
rect 10953 12484 10957 12540
rect 10893 12480 10957 12484
rect 10973 12540 11037 12544
rect 10973 12484 10977 12540
rect 10977 12484 11033 12540
rect 11033 12484 11037 12540
rect 10973 12480 11037 12484
rect 11053 12540 11117 12544
rect 11053 12484 11057 12540
rect 11057 12484 11113 12540
rect 11113 12484 11117 12540
rect 11053 12480 11117 12484
rect 9260 12472 9324 12476
rect 9260 12416 9310 12472
rect 9310 12416 9324 12472
rect 9260 12412 9324 12416
rect 12020 12608 12084 12612
rect 12020 12552 12034 12608
rect 12034 12552 12084 12608
rect 12020 12548 12084 12552
rect 11652 12276 11716 12340
rect 9996 12140 10060 12204
rect 11284 12140 11348 12204
rect 12756 12140 12820 12204
rect 3417 11996 3481 12000
rect 3417 11940 3421 11996
rect 3421 11940 3477 11996
rect 3477 11940 3481 11996
rect 3417 11936 3481 11940
rect 3497 11996 3561 12000
rect 3497 11940 3501 11996
rect 3501 11940 3557 11996
rect 3557 11940 3561 11996
rect 3497 11936 3561 11940
rect 3577 11996 3641 12000
rect 3577 11940 3581 11996
rect 3581 11940 3637 11996
rect 3637 11940 3641 11996
rect 3577 11936 3641 11940
rect 3657 11996 3721 12000
rect 3657 11940 3661 11996
rect 3661 11940 3717 11996
rect 3717 11940 3721 11996
rect 3657 11936 3721 11940
rect 8348 11996 8412 12000
rect 8348 11940 8352 11996
rect 8352 11940 8408 11996
rect 8408 11940 8412 11996
rect 8348 11936 8412 11940
rect 8428 11996 8492 12000
rect 8428 11940 8432 11996
rect 8432 11940 8488 11996
rect 8488 11940 8492 11996
rect 8428 11936 8492 11940
rect 8508 11996 8572 12000
rect 8508 11940 8512 11996
rect 8512 11940 8568 11996
rect 8568 11940 8572 11996
rect 8508 11936 8572 11940
rect 8588 11996 8652 12000
rect 8588 11940 8592 11996
rect 8592 11940 8648 11996
rect 8648 11940 8652 11996
rect 8588 11936 8652 11940
rect 13278 11996 13342 12000
rect 13278 11940 13282 11996
rect 13282 11940 13338 11996
rect 13338 11940 13342 11996
rect 13278 11936 13342 11940
rect 13358 11996 13422 12000
rect 13358 11940 13362 11996
rect 13362 11940 13418 11996
rect 13418 11940 13422 11996
rect 13358 11936 13422 11940
rect 13438 11996 13502 12000
rect 13438 11940 13442 11996
rect 13442 11940 13498 11996
rect 13498 11940 13502 11996
rect 13438 11936 13502 11940
rect 13518 11996 13582 12000
rect 13518 11940 13522 11996
rect 13522 11940 13578 11996
rect 13578 11940 13582 11996
rect 13518 11936 13582 11940
rect 9996 11928 10060 11932
rect 9996 11872 10010 11928
rect 10010 11872 10060 11928
rect 9996 11868 10060 11872
rect 10548 11868 10612 11932
rect 12572 11868 12636 11932
rect 9628 11596 9692 11660
rect 11468 11596 11532 11660
rect 13860 11732 13924 11796
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 6122 11452 6186 11456
rect 6122 11396 6126 11452
rect 6126 11396 6182 11452
rect 6182 11396 6186 11452
rect 6122 11392 6186 11396
rect 10813 11452 10877 11456
rect 10813 11396 10817 11452
rect 10817 11396 10873 11452
rect 10873 11396 10877 11452
rect 10813 11392 10877 11396
rect 10893 11452 10957 11456
rect 10893 11396 10897 11452
rect 10897 11396 10953 11452
rect 10953 11396 10957 11452
rect 10893 11392 10957 11396
rect 10973 11452 11037 11456
rect 10973 11396 10977 11452
rect 10977 11396 11033 11452
rect 11033 11396 11037 11452
rect 10973 11392 11037 11396
rect 11053 11452 11117 11456
rect 11053 11396 11057 11452
rect 11057 11396 11113 11452
rect 11113 11396 11117 11452
rect 11053 11392 11117 11396
rect 10180 11384 10244 11388
rect 10180 11328 10230 11384
rect 10230 11328 10244 11384
rect 10180 11324 10244 11328
rect 12940 11324 13004 11388
rect 13860 11188 13924 11252
rect 9076 10976 9140 10980
rect 9076 10920 9090 10976
rect 9090 10920 9140 10976
rect 9076 10916 9140 10920
rect 10180 10916 10244 10980
rect 3417 10908 3481 10912
rect 3417 10852 3421 10908
rect 3421 10852 3477 10908
rect 3477 10852 3481 10908
rect 3417 10848 3481 10852
rect 3497 10908 3561 10912
rect 3497 10852 3501 10908
rect 3501 10852 3557 10908
rect 3557 10852 3561 10908
rect 3497 10848 3561 10852
rect 3577 10908 3641 10912
rect 3577 10852 3581 10908
rect 3581 10852 3637 10908
rect 3637 10852 3641 10908
rect 3577 10848 3641 10852
rect 3657 10908 3721 10912
rect 3657 10852 3661 10908
rect 3661 10852 3717 10908
rect 3717 10852 3721 10908
rect 3657 10848 3721 10852
rect 8348 10908 8412 10912
rect 8348 10852 8352 10908
rect 8352 10852 8408 10908
rect 8408 10852 8412 10908
rect 8348 10848 8412 10852
rect 8428 10908 8492 10912
rect 8428 10852 8432 10908
rect 8432 10852 8488 10908
rect 8488 10852 8492 10908
rect 8428 10848 8492 10852
rect 8508 10908 8572 10912
rect 8508 10852 8512 10908
rect 8512 10852 8568 10908
rect 8568 10852 8572 10908
rect 8508 10848 8572 10852
rect 8588 10908 8652 10912
rect 8588 10852 8592 10908
rect 8592 10852 8648 10908
rect 8648 10852 8652 10908
rect 8588 10848 8652 10852
rect 13278 10908 13342 10912
rect 13278 10852 13282 10908
rect 13282 10852 13338 10908
rect 13338 10852 13342 10908
rect 13278 10848 13342 10852
rect 13358 10908 13422 10912
rect 13358 10852 13362 10908
rect 13362 10852 13418 10908
rect 13418 10852 13422 10908
rect 13358 10848 13422 10852
rect 13438 10908 13502 10912
rect 13438 10852 13442 10908
rect 13442 10852 13498 10908
rect 13498 10852 13502 10908
rect 13438 10848 13502 10852
rect 13518 10908 13582 10912
rect 13518 10852 13522 10908
rect 13522 10852 13578 10908
rect 13578 10852 13582 10908
rect 13518 10848 13582 10852
rect 12388 10780 12452 10844
rect 14412 10644 14476 10708
rect 9444 10568 9508 10572
rect 9444 10512 9458 10568
rect 9458 10512 9508 10568
rect 9444 10508 9508 10512
rect 11652 10568 11716 10572
rect 11652 10512 11702 10568
rect 11702 10512 11716 10568
rect 11652 10508 11716 10512
rect 12020 10372 12084 10436
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 6122 10364 6186 10368
rect 6122 10308 6126 10364
rect 6126 10308 6182 10364
rect 6182 10308 6186 10364
rect 6122 10304 6186 10308
rect 10813 10364 10877 10368
rect 10813 10308 10817 10364
rect 10817 10308 10873 10364
rect 10873 10308 10877 10364
rect 10813 10304 10877 10308
rect 10893 10364 10957 10368
rect 10893 10308 10897 10364
rect 10897 10308 10953 10364
rect 10953 10308 10957 10364
rect 10893 10304 10957 10308
rect 10973 10364 11037 10368
rect 10973 10308 10977 10364
rect 10977 10308 11033 10364
rect 11033 10308 11037 10364
rect 10973 10304 11037 10308
rect 11053 10364 11117 10368
rect 11053 10308 11057 10364
rect 11057 10308 11113 10364
rect 11113 10308 11117 10364
rect 11053 10304 11117 10308
rect 12204 10100 12268 10164
rect 13676 10100 13740 10164
rect 3417 9820 3481 9824
rect 3417 9764 3421 9820
rect 3421 9764 3477 9820
rect 3477 9764 3481 9820
rect 3417 9760 3481 9764
rect 3497 9820 3561 9824
rect 3497 9764 3501 9820
rect 3501 9764 3557 9820
rect 3557 9764 3561 9820
rect 3497 9760 3561 9764
rect 3577 9820 3641 9824
rect 3577 9764 3581 9820
rect 3581 9764 3637 9820
rect 3637 9764 3641 9820
rect 3577 9760 3641 9764
rect 3657 9820 3721 9824
rect 3657 9764 3661 9820
rect 3661 9764 3717 9820
rect 3717 9764 3721 9820
rect 3657 9760 3721 9764
rect 8348 9820 8412 9824
rect 8348 9764 8352 9820
rect 8352 9764 8408 9820
rect 8408 9764 8412 9820
rect 8348 9760 8412 9764
rect 8428 9820 8492 9824
rect 8428 9764 8432 9820
rect 8432 9764 8488 9820
rect 8488 9764 8492 9820
rect 8428 9760 8492 9764
rect 8508 9820 8572 9824
rect 8508 9764 8512 9820
rect 8512 9764 8568 9820
rect 8568 9764 8572 9820
rect 8508 9760 8572 9764
rect 8588 9820 8652 9824
rect 8588 9764 8592 9820
rect 8592 9764 8648 9820
rect 8648 9764 8652 9820
rect 8588 9760 8652 9764
rect 13278 9820 13342 9824
rect 13278 9764 13282 9820
rect 13282 9764 13338 9820
rect 13338 9764 13342 9820
rect 13278 9760 13342 9764
rect 13358 9820 13422 9824
rect 13358 9764 13362 9820
rect 13362 9764 13418 9820
rect 13418 9764 13422 9820
rect 13358 9760 13422 9764
rect 13438 9820 13502 9824
rect 13438 9764 13442 9820
rect 13442 9764 13498 9820
rect 13498 9764 13502 9820
rect 13438 9760 13502 9764
rect 13518 9820 13582 9824
rect 13518 9764 13522 9820
rect 13522 9764 13578 9820
rect 13578 9764 13582 9820
rect 13518 9760 13582 9764
rect 12572 9752 12636 9756
rect 12572 9696 12622 9752
rect 12622 9696 12636 9752
rect 12572 9692 12636 9696
rect 9996 9556 10060 9620
rect 13124 9556 13188 9620
rect 8892 9284 8956 9348
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 6122 9276 6186 9280
rect 6122 9220 6126 9276
rect 6126 9220 6182 9276
rect 6182 9220 6186 9276
rect 6122 9216 6186 9220
rect 11284 9284 11348 9348
rect 13124 9344 13188 9348
rect 13124 9288 13138 9344
rect 13138 9288 13188 9344
rect 13124 9284 13188 9288
rect 10813 9276 10877 9280
rect 10813 9220 10817 9276
rect 10817 9220 10873 9276
rect 10873 9220 10877 9276
rect 10813 9216 10877 9220
rect 10893 9276 10957 9280
rect 10893 9220 10897 9276
rect 10897 9220 10953 9276
rect 10953 9220 10957 9276
rect 10893 9216 10957 9220
rect 10973 9276 11037 9280
rect 10973 9220 10977 9276
rect 10977 9220 11033 9276
rect 11033 9220 11037 9276
rect 10973 9216 11037 9220
rect 11053 9276 11117 9280
rect 11053 9220 11057 9276
rect 11057 9220 11113 9276
rect 11113 9220 11117 9276
rect 11053 9216 11117 9220
rect 12940 9148 13004 9212
rect 4476 8936 4540 8940
rect 4476 8880 4526 8936
rect 4526 8880 4540 8936
rect 4476 8876 4540 8880
rect 10548 8876 10612 8940
rect 11284 8876 11348 8940
rect 11652 8876 11716 8940
rect 12388 8876 12452 8940
rect 14044 8876 14108 8940
rect 12388 8740 12452 8804
rect 3417 8732 3481 8736
rect 3417 8676 3421 8732
rect 3421 8676 3477 8732
rect 3477 8676 3481 8732
rect 3417 8672 3481 8676
rect 3497 8732 3561 8736
rect 3497 8676 3501 8732
rect 3501 8676 3557 8732
rect 3557 8676 3561 8732
rect 3497 8672 3561 8676
rect 3577 8732 3641 8736
rect 3577 8676 3581 8732
rect 3581 8676 3637 8732
rect 3637 8676 3641 8732
rect 3577 8672 3641 8676
rect 3657 8732 3721 8736
rect 3657 8676 3661 8732
rect 3661 8676 3717 8732
rect 3717 8676 3721 8732
rect 3657 8672 3721 8676
rect 8348 8732 8412 8736
rect 8348 8676 8352 8732
rect 8352 8676 8408 8732
rect 8408 8676 8412 8732
rect 8348 8672 8412 8676
rect 8428 8732 8492 8736
rect 8428 8676 8432 8732
rect 8432 8676 8488 8732
rect 8488 8676 8492 8732
rect 8428 8672 8492 8676
rect 8508 8732 8572 8736
rect 8508 8676 8512 8732
rect 8512 8676 8568 8732
rect 8568 8676 8572 8732
rect 8508 8672 8572 8676
rect 8588 8732 8652 8736
rect 8588 8676 8592 8732
rect 8592 8676 8648 8732
rect 8648 8676 8652 8732
rect 8588 8672 8652 8676
rect 13278 8732 13342 8736
rect 13278 8676 13282 8732
rect 13282 8676 13338 8732
rect 13338 8676 13342 8732
rect 13278 8672 13342 8676
rect 13358 8732 13422 8736
rect 13358 8676 13362 8732
rect 13362 8676 13418 8732
rect 13418 8676 13422 8732
rect 13358 8672 13422 8676
rect 13438 8732 13502 8736
rect 13438 8676 13442 8732
rect 13442 8676 13498 8732
rect 13498 8676 13502 8732
rect 13438 8672 13502 8676
rect 13518 8732 13582 8736
rect 13518 8676 13522 8732
rect 13522 8676 13578 8732
rect 13578 8676 13582 8732
rect 13518 8672 13582 8676
rect 9628 8604 9692 8668
rect 9444 8468 9508 8532
rect 12756 8604 12820 8668
rect 12388 8392 12452 8396
rect 12388 8336 12438 8392
rect 12438 8336 12452 8392
rect 12388 8332 12452 8336
rect 9260 8256 9324 8260
rect 9260 8200 9274 8256
rect 9274 8200 9324 8256
rect 9260 8196 9324 8200
rect 9444 8196 9508 8260
rect 12388 8256 12452 8260
rect 12388 8200 12402 8256
rect 12402 8200 12452 8256
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 6122 8188 6186 8192
rect 6122 8132 6126 8188
rect 6126 8132 6182 8188
rect 6182 8132 6186 8188
rect 6122 8128 6186 8132
rect 12388 8196 12452 8200
rect 10813 8188 10877 8192
rect 10813 8132 10817 8188
rect 10817 8132 10873 8188
rect 10873 8132 10877 8188
rect 10813 8128 10877 8132
rect 10893 8188 10957 8192
rect 10893 8132 10897 8188
rect 10897 8132 10953 8188
rect 10953 8132 10957 8188
rect 10893 8128 10957 8132
rect 10973 8188 11037 8192
rect 10973 8132 10977 8188
rect 10977 8132 11033 8188
rect 11033 8132 11037 8188
rect 10973 8128 11037 8132
rect 11053 8188 11117 8192
rect 11053 8132 11057 8188
rect 11057 8132 11113 8188
rect 11113 8132 11117 8188
rect 11053 8128 11117 8132
rect 14044 8060 14108 8124
rect 7972 7924 8036 7988
rect 8156 7924 8220 7988
rect 12020 7788 12084 7852
rect 13860 7788 13924 7852
rect 3417 7644 3481 7648
rect 3417 7588 3421 7644
rect 3421 7588 3477 7644
rect 3477 7588 3481 7644
rect 3417 7584 3481 7588
rect 3497 7644 3561 7648
rect 3497 7588 3501 7644
rect 3501 7588 3557 7644
rect 3557 7588 3561 7644
rect 3497 7584 3561 7588
rect 3577 7644 3641 7648
rect 3577 7588 3581 7644
rect 3581 7588 3637 7644
rect 3637 7588 3641 7644
rect 3577 7584 3641 7588
rect 3657 7644 3721 7648
rect 3657 7588 3661 7644
rect 3661 7588 3717 7644
rect 3717 7588 3721 7644
rect 3657 7584 3721 7588
rect 8348 7644 8412 7648
rect 8348 7588 8352 7644
rect 8352 7588 8408 7644
rect 8408 7588 8412 7644
rect 8348 7584 8412 7588
rect 8428 7644 8492 7648
rect 8428 7588 8432 7644
rect 8432 7588 8488 7644
rect 8488 7588 8492 7644
rect 8428 7584 8492 7588
rect 8508 7644 8572 7648
rect 8508 7588 8512 7644
rect 8512 7588 8568 7644
rect 8568 7588 8572 7644
rect 8508 7584 8572 7588
rect 8588 7644 8652 7648
rect 8588 7588 8592 7644
rect 8592 7588 8648 7644
rect 8648 7588 8652 7644
rect 8588 7584 8652 7588
rect 13278 7644 13342 7648
rect 13278 7588 13282 7644
rect 13282 7588 13338 7644
rect 13338 7588 13342 7644
rect 13278 7584 13342 7588
rect 13358 7644 13422 7648
rect 13358 7588 13362 7644
rect 13362 7588 13418 7644
rect 13418 7588 13422 7644
rect 13358 7584 13422 7588
rect 13438 7644 13502 7648
rect 13438 7588 13442 7644
rect 13442 7588 13498 7644
rect 13498 7588 13502 7644
rect 13438 7584 13502 7588
rect 13518 7644 13582 7648
rect 13518 7588 13522 7644
rect 13522 7588 13578 7644
rect 13578 7588 13582 7644
rect 13518 7584 13582 7588
rect 9076 7516 9140 7580
rect 11284 7108 11348 7172
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 6122 7100 6186 7104
rect 6122 7044 6126 7100
rect 6126 7044 6182 7100
rect 6182 7044 6186 7100
rect 6122 7040 6186 7044
rect 10813 7100 10877 7104
rect 10813 7044 10817 7100
rect 10817 7044 10873 7100
rect 10873 7044 10877 7100
rect 10813 7040 10877 7044
rect 10893 7100 10957 7104
rect 10893 7044 10897 7100
rect 10897 7044 10953 7100
rect 10953 7044 10957 7100
rect 10893 7040 10957 7044
rect 10973 7100 11037 7104
rect 10973 7044 10977 7100
rect 10977 7044 11033 7100
rect 11033 7044 11037 7100
rect 10973 7040 11037 7044
rect 11053 7100 11117 7104
rect 11053 7044 11057 7100
rect 11057 7044 11113 7100
rect 11113 7044 11117 7100
rect 11053 7040 11117 7044
rect 10180 6972 10244 7036
rect 11836 6836 11900 6900
rect 12388 6700 12452 6764
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 8156 6080 8220 6084
rect 8156 6024 8206 6080
rect 8206 6024 8220 6080
rect 8156 6020 8220 6024
rect 11836 6020 11900 6084
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 8892 5476 8956 5540
rect 13124 5612 13188 5676
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 8892 5340 8956 5404
rect 4292 5204 4356 5268
rect 14412 5068 14476 5132
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 10180 4932 10244 4996
rect 11284 4992 11348 4996
rect 11284 4936 11298 4992
rect 11298 4936 11348 4992
rect 11284 4932 11348 4936
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 9444 4856 9508 4860
rect 9444 4800 9458 4856
rect 9458 4800 9508 4856
rect 9444 4796 9508 4800
rect 11836 4388 11900 4452
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 9628 4252 9692 4316
rect 12756 4116 12820 4180
rect 12940 4116 13004 4180
rect 10364 3844 10428 3908
rect 11652 3844 11716 3908
rect 14044 3904 14108 3908
rect 14044 3848 14094 3904
rect 14094 3848 14108 3904
rect 14044 3844 14108 3848
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 8892 3360 8956 3364
rect 8892 3304 8906 3360
rect 8906 3304 8956 3360
rect 8892 3300 8956 3304
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 8156 3224 8220 3228
rect 10548 3300 10612 3364
rect 12572 3360 12636 3364
rect 12572 3304 12622 3360
rect 12622 3304 12636 3360
rect 12572 3300 12636 3304
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 8156 3168 8206 3224
rect 8206 3168 8220 3224
rect 8156 3164 8220 3168
rect 10180 3164 10244 3228
rect 9812 3088 9876 3092
rect 9812 3032 9826 3088
rect 9826 3032 9876 3088
rect 9812 3028 9876 3032
rect 12204 3028 12268 3092
rect 12940 3088 13004 3092
rect 12940 3032 12954 3088
rect 12954 3032 13004 3088
rect 12940 3028 13004 3032
rect 13676 2816 13740 2820
rect 13676 2760 13690 2816
rect 13690 2760 13740 2816
rect 13676 2756 13740 2760
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 9444 2620 9508 2684
rect 9996 2680 10060 2684
rect 9996 2624 10010 2680
rect 10010 2624 10060 2680
rect 9996 2620 10060 2624
rect 11468 2680 11532 2684
rect 11468 2624 11482 2680
rect 11482 2624 11532 2680
rect 11468 2620 11532 2624
rect 4476 2484 4540 2548
rect 9260 2484 9324 2548
rect 12940 2544 13004 2548
rect 12940 2488 12954 2544
rect 12954 2488 13004 2544
rect 12940 2484 13004 2488
rect 12020 2212 12084 2276
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
rect 9076 1940 9140 2004
<< metal4 >>
rect 13123 17644 13189 17645
rect 13123 17580 13124 17644
rect 13188 17580 13189 17644
rect 13123 17579 13189 17580
rect 3409 17440 3729 17456
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 16352 3729 17376
rect 5874 16896 6195 17456
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6195 16896
rect 4291 16828 4357 16829
rect 4291 16764 4292 16828
rect 4356 16764 4357 16828
rect 4291 16763 4357 16764
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 15264 3729 16288
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 14176 3729 15200
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 13088 3729 14112
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 12000 3729 13024
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 10912 3729 11936
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 9824 3729 10848
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 8736 3729 9760
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 7648 3729 8672
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 6560 3729 7584
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 5472 3729 6496
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 4294 5269 4354 16763
rect 5874 15808 6195 16832
rect 8340 17440 8660 17456
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 16352 8660 17376
rect 9811 17236 9877 17237
rect 9811 17172 9812 17236
rect 9876 17172 9877 17236
rect 9811 17171 9877 17172
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 7971 16284 8037 16285
rect 7971 16220 7972 16284
rect 8036 16220 8037 16284
rect 7971 16219 8037 16220
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6195 15808
rect 5874 14720 6195 15744
rect 7974 14789 8034 16219
rect 8155 16148 8221 16149
rect 8155 16084 8156 16148
rect 8220 16084 8221 16148
rect 8155 16083 8221 16084
rect 8158 15741 8218 16083
rect 8155 15740 8221 15741
rect 8155 15676 8156 15740
rect 8220 15676 8221 15740
rect 8155 15675 8221 15676
rect 8340 15264 8660 16288
rect 9259 16284 9325 16285
rect 9259 16220 9260 16284
rect 9324 16220 9325 16284
rect 9259 16219 9325 16220
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 7971 14788 8037 14789
rect 7971 14724 7972 14788
rect 8036 14724 8037 14788
rect 7971 14723 8037 14724
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6195 14720
rect 5874 13632 6195 14656
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6195 13632
rect 5874 12544 6195 13568
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6195 12544
rect 5874 11456 6195 12480
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6195 11456
rect 5874 10368 6195 11392
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6195 10368
rect 5874 9280 6195 10304
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6195 9280
rect 4475 8940 4541 8941
rect 4475 8876 4476 8940
rect 4540 8876 4541 8940
rect 4475 8875 4541 8876
rect 4291 5268 4357 5269
rect 4291 5204 4292 5268
rect 4356 5204 4357 5268
rect 4291 5203 4357 5204
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 3296 3729 4320
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 2208 3729 3232
rect 4478 2549 4538 8875
rect 5874 8192 6195 9216
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6195 8192
rect 5874 7104 6195 8128
rect 8340 14176 8660 15200
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 13088 8660 14112
rect 9075 13836 9141 13837
rect 9075 13772 9076 13836
rect 9140 13772 9141 13836
rect 9075 13771 9141 13772
rect 8891 13156 8957 13157
rect 8891 13092 8892 13156
rect 8956 13092 8957 13156
rect 8891 13091 8957 13092
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 12000 8660 13024
rect 8894 12613 8954 13091
rect 8891 12612 8957 12613
rect 8891 12548 8892 12612
rect 8956 12548 8957 12612
rect 8891 12547 8957 12548
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 10912 8660 11936
rect 9078 10981 9138 13771
rect 9262 13021 9322 16219
rect 9627 15740 9693 15741
rect 9627 15676 9628 15740
rect 9692 15676 9693 15740
rect 9627 15675 9693 15676
rect 9443 14108 9509 14109
rect 9443 14044 9444 14108
rect 9508 14044 9509 14108
rect 9443 14043 9509 14044
rect 9259 13020 9325 13021
rect 9259 12956 9260 13020
rect 9324 12956 9325 13020
rect 9259 12955 9325 12956
rect 9262 12477 9322 12955
rect 9259 12476 9325 12477
rect 9259 12412 9260 12476
rect 9324 12412 9325 12476
rect 9259 12411 9325 12412
rect 9075 10980 9141 10981
rect 9075 10916 9076 10980
rect 9140 10916 9141 10980
rect 9075 10915 9141 10916
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 9824 8660 10848
rect 9446 10573 9506 14043
rect 9630 11661 9690 15675
rect 9627 11660 9693 11661
rect 9627 11596 9628 11660
rect 9692 11596 9693 11660
rect 9627 11595 9693 11596
rect 9443 10572 9509 10573
rect 9443 10508 9444 10572
rect 9508 10508 9509 10572
rect 9443 10507 9509 10508
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 8736 8660 9760
rect 8891 9348 8957 9349
rect 8891 9284 8892 9348
rect 8956 9284 8957 9348
rect 8891 9283 8957 9284
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 7971 7988 8037 7989
rect 7971 7924 7972 7988
rect 8036 7924 8037 7988
rect 7971 7923 8037 7924
rect 8155 7988 8221 7989
rect 8155 7924 8156 7988
rect 8220 7924 8221 7988
rect 8155 7923 8221 7924
rect 7974 7850 8034 7923
rect 8158 7850 8218 7923
rect 7974 7790 8218 7850
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6195 7104
rect 5874 6016 6195 7040
rect 8340 7648 8660 8672
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 6560 8660 7584
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8155 6084 8221 6085
rect 8155 6020 8156 6084
rect 8220 6020 8221 6084
rect 8155 6019 8221 6020
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5874 3840 6195 4864
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5874 2752 6195 3776
rect 8158 3229 8218 6019
rect 8340 5472 8660 6496
rect 8894 5541 8954 9283
rect 9630 8669 9690 11595
rect 9627 8668 9693 8669
rect 9627 8604 9628 8668
rect 9692 8604 9693 8668
rect 9627 8603 9693 8604
rect 9443 8532 9509 8533
rect 9443 8468 9444 8532
rect 9508 8468 9509 8532
rect 9443 8467 9509 8468
rect 9446 8261 9506 8467
rect 9259 8260 9325 8261
rect 9259 8196 9260 8260
rect 9324 8196 9325 8260
rect 9259 8195 9325 8196
rect 9443 8260 9509 8261
rect 9443 8196 9444 8260
rect 9508 8196 9509 8260
rect 9443 8195 9509 8196
rect 9075 7580 9141 7581
rect 9075 7516 9076 7580
rect 9140 7516 9141 7580
rect 9075 7515 9141 7516
rect 8891 5540 8957 5541
rect 8891 5476 8892 5540
rect 8956 5476 8957 5540
rect 8891 5475 8957 5476
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8891 5404 8957 5405
rect 8891 5340 8892 5404
rect 8956 5340 8957 5404
rect 8891 5339 8957 5340
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 3296 8660 4320
rect 8894 3365 8954 5339
rect 8891 3364 8957 3365
rect 8891 3300 8892 3364
rect 8956 3300 8957 3364
rect 8891 3299 8957 3300
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8155 3228 8221 3229
rect 8155 3164 8156 3228
rect 8220 3164 8221 3228
rect 8155 3163 8221 3164
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 4475 2548 4541 2549
rect 4475 2484 4476 2548
rect 4540 2484 4541 2548
rect 4475 2483 4541 2484
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 5874 2128 6195 2688
rect 8340 2208 8660 3232
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 9078 2005 9138 7515
rect 9262 2549 9322 8195
rect 9443 4860 9509 4861
rect 9443 4796 9444 4860
rect 9508 4796 9509 4860
rect 9443 4795 9509 4796
rect 9446 2685 9506 4795
rect 9630 4317 9690 8603
rect 9627 4316 9693 4317
rect 9627 4252 9628 4316
rect 9692 4252 9693 4316
rect 9627 4251 9693 4252
rect 9814 3093 9874 17171
rect 10805 16896 11125 17456
rect 11283 17100 11349 17101
rect 11283 17036 11284 17100
rect 11348 17036 11349 17100
rect 11283 17035 11349 17036
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 9995 16828 10061 16829
rect 9995 16764 9996 16828
rect 10060 16764 10061 16828
rect 9995 16763 10061 16764
rect 9998 16285 10058 16763
rect 9995 16284 10061 16285
rect 9995 16220 9996 16284
rect 10060 16220 10061 16284
rect 9995 16219 10061 16220
rect 10805 15808 11125 16832
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 9995 15740 10061 15741
rect 9995 15676 9996 15740
rect 10060 15676 10061 15740
rect 9995 15675 10061 15676
rect 9998 12205 10058 15675
rect 10547 14788 10613 14789
rect 10547 14724 10548 14788
rect 10612 14724 10613 14788
rect 10547 14723 10613 14724
rect 10363 13836 10429 13837
rect 10363 13772 10364 13836
rect 10428 13772 10429 13836
rect 10363 13771 10429 13772
rect 10179 12748 10245 12749
rect 10179 12684 10180 12748
rect 10244 12684 10245 12748
rect 10179 12683 10245 12684
rect 9995 12204 10061 12205
rect 9995 12140 9996 12204
rect 10060 12140 10061 12204
rect 9995 12139 10061 12140
rect 9995 11932 10061 11933
rect 9995 11868 9996 11932
rect 10060 11868 10061 11932
rect 9995 11867 10061 11868
rect 9998 9621 10058 11867
rect 10182 11389 10242 12683
rect 10179 11388 10245 11389
rect 10179 11324 10180 11388
rect 10244 11324 10245 11388
rect 10179 11323 10245 11324
rect 10179 10980 10245 10981
rect 10179 10916 10180 10980
rect 10244 10916 10245 10980
rect 10179 10915 10245 10916
rect 9995 9620 10061 9621
rect 9995 9556 9996 9620
rect 10060 9556 10061 9620
rect 9995 9555 10061 9556
rect 9811 3092 9877 3093
rect 9811 3028 9812 3092
rect 9876 3028 9877 3092
rect 9811 3027 9877 3028
rect 9998 2685 10058 9555
rect 10182 7037 10242 10915
rect 10179 7036 10245 7037
rect 10179 6972 10180 7036
rect 10244 6972 10245 7036
rect 10179 6971 10245 6972
rect 10179 4996 10245 4997
rect 10179 4932 10180 4996
rect 10244 4932 10245 4996
rect 10179 4931 10245 4932
rect 10182 3229 10242 4931
rect 10366 3909 10426 13771
rect 10550 11933 10610 14723
rect 10805 14720 11125 15744
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 13632 11125 14656
rect 11286 14517 11346 17035
rect 11835 15332 11901 15333
rect 11835 15268 11836 15332
rect 11900 15268 11901 15332
rect 11835 15267 11901 15268
rect 11283 14516 11349 14517
rect 11283 14452 11284 14516
rect 11348 14452 11349 14516
rect 11283 14451 11349 14452
rect 11651 14380 11717 14381
rect 11651 14316 11652 14380
rect 11716 14316 11717 14380
rect 11651 14315 11717 14316
rect 11467 14244 11533 14245
rect 11467 14180 11468 14244
rect 11532 14180 11533 14244
rect 11467 14179 11533 14180
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 12544 11125 13568
rect 11283 13020 11349 13021
rect 11283 12956 11284 13020
rect 11348 12956 11349 13020
rect 11283 12955 11349 12956
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10547 11932 10613 11933
rect 10547 11868 10548 11932
rect 10612 11868 10613 11932
rect 10547 11867 10613 11868
rect 10805 11456 11125 12480
rect 11286 12205 11346 12955
rect 11470 12749 11530 14179
rect 11467 12748 11533 12749
rect 11467 12684 11468 12748
rect 11532 12684 11533 12748
rect 11467 12683 11533 12684
rect 11467 12612 11533 12613
rect 11467 12548 11468 12612
rect 11532 12548 11533 12612
rect 11467 12547 11533 12548
rect 11283 12204 11349 12205
rect 11283 12140 11284 12204
rect 11348 12140 11349 12204
rect 11283 12139 11349 12140
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 10368 11125 11392
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 9280 11125 10304
rect 11286 9349 11346 12139
rect 11470 11930 11530 12547
rect 11654 12341 11714 14315
rect 11651 12340 11717 12341
rect 11651 12276 11652 12340
rect 11716 12276 11717 12340
rect 11651 12275 11717 12276
rect 11470 11870 11714 11930
rect 11467 11660 11533 11661
rect 11467 11596 11468 11660
rect 11532 11596 11533 11660
rect 11467 11595 11533 11596
rect 11283 9348 11349 9349
rect 11283 9284 11284 9348
rect 11348 9284 11349 9348
rect 11283 9283 11349 9284
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10547 8940 10613 8941
rect 10547 8876 10548 8940
rect 10612 8876 10613 8940
rect 10547 8875 10613 8876
rect 10363 3908 10429 3909
rect 10363 3844 10364 3908
rect 10428 3844 10429 3908
rect 10363 3843 10429 3844
rect 10550 3365 10610 8875
rect 10805 8192 11125 9216
rect 11286 8941 11346 9283
rect 11283 8940 11349 8941
rect 11283 8876 11284 8940
rect 11348 8876 11349 8940
rect 11283 8875 11349 8876
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 7104 11125 8128
rect 11283 7172 11349 7173
rect 11283 7108 11284 7172
rect 11348 7108 11349 7172
rect 11283 7107 11349 7108
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 6016 11125 7040
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 11286 4997 11346 7107
rect 11283 4996 11349 4997
rect 11283 4932 11284 4996
rect 11348 4932 11349 4996
rect 11283 4931 11349 4932
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 3840 11125 4864
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10547 3364 10613 3365
rect 10547 3300 10548 3364
rect 10612 3300 10613 3364
rect 10547 3299 10613 3300
rect 10179 3228 10245 3229
rect 10179 3164 10180 3228
rect 10244 3164 10245 3228
rect 10179 3163 10245 3164
rect 10805 2752 11125 3776
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 9443 2684 9509 2685
rect 9443 2620 9444 2684
rect 9508 2620 9509 2684
rect 9443 2619 9509 2620
rect 9995 2684 10061 2685
rect 9995 2620 9996 2684
rect 10060 2620 10061 2684
rect 9995 2619 10061 2620
rect 9259 2548 9325 2549
rect 9259 2484 9260 2548
rect 9324 2484 9325 2548
rect 9259 2483 9325 2484
rect 10805 2128 11125 2688
rect 11470 2685 11530 11595
rect 11654 10573 11714 11870
rect 11651 10572 11717 10573
rect 11651 10508 11652 10572
rect 11716 10508 11717 10572
rect 11651 10507 11717 10508
rect 11651 8940 11717 8941
rect 11651 8876 11652 8940
rect 11716 8876 11717 8940
rect 11651 8875 11717 8876
rect 11654 3909 11714 8875
rect 11838 6901 11898 15267
rect 12939 14788 13005 14789
rect 12939 14724 12940 14788
rect 13004 14724 13005 14788
rect 12939 14723 13005 14724
rect 12203 14516 12269 14517
rect 12203 14452 12204 14516
rect 12268 14452 12269 14516
rect 12203 14451 12269 14452
rect 12019 12612 12085 12613
rect 12019 12548 12020 12612
rect 12084 12548 12085 12612
rect 12019 12547 12085 12548
rect 12022 10437 12082 12547
rect 12019 10436 12085 10437
rect 12019 10372 12020 10436
rect 12084 10372 12085 10436
rect 12019 10371 12085 10372
rect 12206 10165 12266 14451
rect 12387 13972 12453 13973
rect 12387 13908 12388 13972
rect 12452 13908 12453 13972
rect 12387 13907 12453 13908
rect 12390 10845 12450 13907
rect 12942 13154 13002 14723
rect 13126 13293 13186 17579
rect 13270 17440 13590 17456
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 13270 16352 13590 17376
rect 14043 16828 14109 16829
rect 14043 16764 14044 16828
rect 14108 16764 14109 16828
rect 14043 16763 14109 16764
rect 13859 16692 13925 16693
rect 13859 16628 13860 16692
rect 13924 16628 13925 16692
rect 13859 16627 13925 16628
rect 13675 16556 13741 16557
rect 13675 16492 13676 16556
rect 13740 16492 13741 16556
rect 13675 16491 13741 16492
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 15264 13590 16288
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 14176 13590 15200
rect 13678 14925 13738 16491
rect 13675 14924 13741 14925
rect 13675 14860 13676 14924
rect 13740 14860 13741 14924
rect 13675 14859 13741 14860
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13123 13292 13189 13293
rect 13123 13228 13124 13292
rect 13188 13228 13189 13292
rect 13123 13227 13189 13228
rect 12942 13094 13186 13154
rect 12755 12204 12821 12205
rect 12755 12140 12756 12204
rect 12820 12140 12821 12204
rect 12755 12139 12821 12140
rect 12571 11932 12637 11933
rect 12571 11868 12572 11932
rect 12636 11868 12637 11932
rect 12571 11867 12637 11868
rect 12387 10844 12453 10845
rect 12387 10780 12388 10844
rect 12452 10780 12453 10844
rect 12387 10779 12453 10780
rect 12574 10570 12634 11867
rect 12390 10510 12634 10570
rect 12203 10164 12269 10165
rect 12203 10100 12204 10164
rect 12268 10100 12269 10164
rect 12203 10099 12269 10100
rect 12019 7852 12085 7853
rect 12019 7788 12020 7852
rect 12084 7788 12085 7852
rect 12019 7787 12085 7788
rect 11835 6900 11901 6901
rect 11835 6836 11836 6900
rect 11900 6836 11901 6900
rect 11835 6835 11901 6836
rect 11835 6084 11901 6085
rect 11835 6020 11836 6084
rect 11900 6020 11901 6084
rect 11835 6019 11901 6020
rect 11838 4453 11898 6019
rect 11835 4452 11901 4453
rect 11835 4388 11836 4452
rect 11900 4388 11901 4452
rect 11835 4387 11901 4388
rect 11651 3908 11717 3909
rect 11651 3844 11652 3908
rect 11716 3844 11717 3908
rect 11651 3843 11717 3844
rect 11467 2684 11533 2685
rect 11467 2620 11468 2684
rect 11532 2620 11533 2684
rect 11467 2619 11533 2620
rect 12022 2277 12082 7787
rect 12206 3093 12266 10099
rect 12390 8941 12450 10510
rect 12571 9756 12637 9757
rect 12571 9692 12572 9756
rect 12636 9692 12637 9756
rect 12571 9691 12637 9692
rect 12387 8940 12453 8941
rect 12387 8876 12388 8940
rect 12452 8876 12453 8940
rect 12387 8875 12453 8876
rect 12387 8804 12453 8805
rect 12387 8740 12388 8804
rect 12452 8740 12453 8804
rect 12387 8739 12453 8740
rect 12390 8397 12450 8739
rect 12387 8396 12453 8397
rect 12387 8332 12388 8396
rect 12452 8332 12453 8396
rect 12387 8331 12453 8332
rect 12387 8260 12453 8261
rect 12387 8196 12388 8260
rect 12452 8196 12453 8260
rect 12387 8195 12453 8196
rect 12390 6765 12450 8195
rect 12387 6764 12453 6765
rect 12387 6700 12388 6764
rect 12452 6700 12453 6764
rect 12387 6699 12453 6700
rect 12574 3365 12634 9691
rect 12758 8669 12818 12139
rect 12939 11388 13005 11389
rect 12939 11324 12940 11388
rect 13004 11324 13005 11388
rect 12939 11323 13005 11324
rect 12942 9213 13002 11323
rect 13126 9621 13186 13094
rect 13270 13088 13590 14112
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 12000 13590 13024
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 10912 13590 11936
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 9824 13590 10848
rect 13678 10165 13738 14859
rect 13862 11797 13922 16627
rect 14046 12749 14106 16763
rect 14043 12748 14109 12749
rect 14043 12684 14044 12748
rect 14108 12684 14109 12748
rect 14043 12683 14109 12684
rect 13859 11796 13925 11797
rect 13859 11732 13860 11796
rect 13924 11732 13925 11796
rect 13859 11731 13925 11732
rect 13859 11252 13925 11253
rect 13859 11188 13860 11252
rect 13924 11188 13925 11252
rect 13859 11187 13925 11188
rect 13675 10164 13741 10165
rect 13675 10100 13676 10164
rect 13740 10100 13741 10164
rect 13675 10099 13741 10100
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13123 9620 13189 9621
rect 13123 9556 13124 9620
rect 13188 9556 13189 9620
rect 13123 9555 13189 9556
rect 13123 9348 13189 9349
rect 13123 9284 13124 9348
rect 13188 9284 13189 9348
rect 13123 9283 13189 9284
rect 12939 9212 13005 9213
rect 12939 9148 12940 9212
rect 13004 9148 13005 9212
rect 12939 9147 13005 9148
rect 12755 8668 12821 8669
rect 12755 8604 12756 8668
rect 12820 8604 12821 8668
rect 12755 8603 12821 8604
rect 12758 4181 12818 8603
rect 12942 4181 13002 9147
rect 13126 5677 13186 9283
rect 13270 8736 13590 9760
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 7648 13590 8672
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 6560 13590 7584
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13123 5676 13189 5677
rect 13123 5612 13124 5676
rect 13188 5612 13189 5676
rect 13123 5611 13189 5612
rect 13270 5472 13590 6496
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 12755 4180 12821 4181
rect 12755 4116 12756 4180
rect 12820 4116 12821 4180
rect 12755 4115 12821 4116
rect 12939 4180 13005 4181
rect 12939 4116 12940 4180
rect 13004 4116 13005 4180
rect 12939 4115 13005 4116
rect 12571 3364 12637 3365
rect 12571 3300 12572 3364
rect 12636 3300 12637 3364
rect 12571 3299 12637 3300
rect 13270 3296 13590 4320
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 12203 3092 12269 3093
rect 12203 3028 12204 3092
rect 12268 3028 12269 3092
rect 12203 3027 12269 3028
rect 12939 3092 13005 3093
rect 12939 3028 12940 3092
rect 13004 3028 13005 3092
rect 12939 3027 13005 3028
rect 12942 2549 13002 3027
rect 12939 2548 13005 2549
rect 12939 2484 12940 2548
rect 13004 2484 13005 2548
rect 12939 2483 13005 2484
rect 12019 2276 12085 2277
rect 12019 2212 12020 2276
rect 12084 2212 12085 2276
rect 12019 2211 12085 2212
rect 13270 2208 13590 3232
rect 13678 2821 13738 10099
rect 13862 7853 13922 11187
rect 14046 8941 14106 12683
rect 14411 10708 14477 10709
rect 14411 10644 14412 10708
rect 14476 10644 14477 10708
rect 14411 10643 14477 10644
rect 14043 8940 14109 8941
rect 14043 8876 14044 8940
rect 14108 8876 14109 8940
rect 14043 8875 14109 8876
rect 14043 8124 14109 8125
rect 14043 8060 14044 8124
rect 14108 8060 14109 8124
rect 14043 8059 14109 8060
rect 13859 7852 13925 7853
rect 13859 7788 13860 7852
rect 13924 7788 13925 7852
rect 13859 7787 13925 7788
rect 14046 3909 14106 8059
rect 14414 5133 14474 10643
rect 14411 5132 14477 5133
rect 14411 5068 14412 5132
rect 14476 5068 14477 5132
rect 14411 5067 14477 5068
rect 14043 3908 14109 3909
rect 14043 3844 14044 3908
rect 14108 3844 14109 3908
rect 14043 3843 14109 3844
rect 13675 2820 13741 2821
rect 13675 2756 13676 2820
rect 13740 2756 13741 2820
rect 13675 2755 13741 2756
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2128 13590 2144
rect 9075 2004 9141 2005
rect 9075 1940 9076 2004
rect 9140 1940 9141 2004
rect 9075 1939 9141 1940
use sky130_fd_sc_hd__buf_2  _53_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2116 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2484 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_S_FTB01 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1564 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1606821651
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4876 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1606821651
transform 1 0 3680 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1606821651
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1606821651
transform 1 0 4600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 1606821651
transform 1 0 3312 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1606821651
transform 1 0 4508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4968 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58
timestamp 1606821651
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1606821651
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1606821651
transform 1 0 8648 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1606821651
transform 1 0 7728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1606821651
transform 1 0 8280 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1606821651
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1606821651
transform 1 0 8924 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_right_ipin_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 9292 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1606821651
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1606821651
transform 1 0 9844 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_104
timestamp 1606821651
transform 1 0 10672 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11040 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1606821651
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1606821651
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1606821651
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116
timestamp 1606821651
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 12144 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13616 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_134
timestamp 1606821651
transform 1 0 13432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1606821651
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1606821651
transform 1 0 14444 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606821651
transform 1 0 14812 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 14996 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_147
timestamp 1606821651
transform 1 0 14628 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1606821651
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_153
timestamp 1606821651
transform 1 0 15180 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 1564 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2760 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1606821651
transform 1 0 2392 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4508 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606821651
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_36
timestamp 1606821651
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5704 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_46
timestamp 1606821651
transform 1 0 5336 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7544 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1606821651
transform 1 0 7176 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 9016 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1606821651
transform 1 0 10488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10856 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12052 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1606821651
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1606821651
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 13248 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1606821651
transform 1 0 12880 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1606821651
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1606821651
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1840 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1606821651
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_17
timestamp 1606821651
transform 1 0 2668 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 3036 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4876 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1606821651
transform 1 0 4508 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1606821651
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8648 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1606821651
transform 1 0 8280 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1606821651
transform 1 0 9844 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_91
timestamp 1606821651
transform 1 0 9476 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_104
timestamp 1606821651
transform 1 0 10672 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11040 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1606821651
transform 1 0 11868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1606821651
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13616 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1606821651
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1606821651
transform 1 0 14444 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606821651
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_153
timestamp 1606821651
transform 1 0 15180 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2116 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1606821651
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606821651
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1606821651
transform 1 0 4876 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5244 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_61
timestamp 1606821651
transform 1 0 6716 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7084 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_81
timestamp 1606821651
transform 1 0 8556 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _16_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8924 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1606821651
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1606821651
transform 1 0 10488 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10856 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_115
timestamp 1606821651
transform 1 0 11684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1606821651
transform 1 0 14444 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13248 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp 1606821651
transform 1 0 12880 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1606821651
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1606821651
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1840 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1606821651
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_17
timestamp 1606821651
transform 1 0 2668 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4876 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 3036 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1606821651
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1606821651
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8648 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1606821651
transform 1 0 8280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10488 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_98
timestamp 1606821651
transform 1 0 10120 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1606821651
transform 1 0 11684 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_111
timestamp 1606821651
transform 1 0 11316 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1606821651
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1606821651
transform 1 0 13616 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1606821651
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_132
timestamp 1606821651
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1606821651
transform 1 0 14444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1606821651
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_153
timestamp 1606821651
transform 1 0 15180 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2116 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1606821651
transform 1 0 1840 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1606821651
transform 1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1606821651
transform 1 0 1748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1606821651
transform 1 0 2668 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 3036 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4876 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1606821651
transform 1 0 4232 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606821651
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1606821651
transform 1 0 4508 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 5428 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_43
timestamp 1606821651
transform 1 0 5060 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1606821651
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7268 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 8648 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_63
timestamp 1606821651
transform 1 0 6900 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_83
timestamp 1606821651
transform 1 0 8740 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1606821651
transform 1 0 8280 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1606821651
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1606821651
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1606821651
transform 1 0 10120 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1606821651
transform 1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1606821651
transform 1 0 11500 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1606821651
transform 1 0 11132 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_122
timestamp 1606821651
transform 1 0 12328 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_111
timestamp 1606821651
transform 1 0 11316 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1606821651
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 13616 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13892 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1606821651
transform 1 0 12696 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1606821651
transform 1 0 13524 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1606821651
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1606821651
transform 1 0 14444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1606821651
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_148
timestamp 1606821651
transform 1 0 14720 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1606821651
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1606821651
transform 1 0 15180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2116 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1606821651
transform 1 0 1748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 4232 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606821651
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 5704 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_46
timestamp 1606821651
transform 1 0 5336 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7544 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_66
timestamp 1606821651
transform 1 0 7176 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_86
timestamp 1606821651
transform 1 0 9016 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_102
timestamp 1606821651
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1606821651
transform 1 0 10856 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1606821651
transform 1 0 12052 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_115
timestamp 1606821651
transform 1 0 11684 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1606821651
transform 1 0 14444 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13248 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1606821651
transform 1 0 12880 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1606821651
transform 1 0 14076 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1606821651
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1606821651
transform 1 0 1840 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1606821651
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_17
timestamp 1606821651
transform 1 0 2668 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 3036 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4876 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_37
timestamp 1606821651
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1606821651
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8648 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_78
timestamp 1606821651
transform 1 0 8280 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1606821651
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1606821651
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1606821651
transform 1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_111
timestamp 1606821651
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1606821651
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1606821651
transform 1 0 13616 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1606821651
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_145
timestamp 1606821651
transform 1 0 14444 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1606821651
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1606821651
transform 1 0 15180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2760 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 1564 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1606821651
transform 1 0 2392 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606821651
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 5888 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1606821651
transform 1 0 5520 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7728 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 1606821651
transform 1 0 7360 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1606821651
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_102
timestamp 1606821651
transform 1 0 10488 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10856 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12052 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_115
timestamp 1606821651
transform 1 0 11684 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1606821651
transform 1 0 14444 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13248 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_128
timestamp 1606821651
transform 1 0 12880 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1606821651
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1606821651
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2484 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1606821651
transform 1 0 2116 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4876 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1606821651
transform 1 0 3680 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1606821651
transform 1 0 3312 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_37
timestamp 1606821651
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1606821651
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8648 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_78
timestamp 1606821651
transform 1 0 8280 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1606821651
transform 1 0 9844 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1606821651
transform 1 0 9476 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_104
timestamp 1606821651
transform 1 0 10672 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11040 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1606821651
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1606821651
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1606821651
transform 1 0 13616 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp 1606821651
transform 1 0 13248 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_145
timestamp 1606821651
transform 1 0 14444 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1606821651
transform 1 0 14812 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1606821651
transform 1 0 15180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1564 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 2760 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_14
timestamp 1606821651
transform 1 0 2392 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4232 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1606821651
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_right_ipin_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5888 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_12_43 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5060 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_51
timestamp 1606821651
transform 1 0 5796 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1606821651
transform 1 0 7728 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 8556 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1606821651
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1606821651
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1606821651
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1606821651
transform 1 0 12052 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1606821651
transform 1 0 10856 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_115
timestamp 1606821651
transform 1 0 11684 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1606821651
transform 1 0 14444 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13248 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_128
timestamp 1606821651
transform 1 0 12880 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1606821651
transform 1 0 14076 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1606821651
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1606821651
transform 1 0 2392 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1606821651
transform 1 0 2760 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2116 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2944 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 3772 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4232 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606821651
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 5428 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 5244 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_43
timestamp 1606821651
transform 1 0 5060 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7268 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8648 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1606821651
transform 1 0 8280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_63
timestamp 1606821651
transform 1 0 6900 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_83
timestamp 1606821651
transform 1 0 8740 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1606821651
transform 1 0 9844 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 1606821651
transform 1 0 9476 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_104
timestamp 1606821651
transform 1 0 10672 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606821651
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1606821651
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12052 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1606821651
transform 1 0 11040 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10856 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_117
timestamp 1606821651
transform 1 0 11868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1606821651
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_115
timestamp 1606821651
transform 1 0 11684 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1606821651
transform 1 0 14444 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13616 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1606821651
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1606821651
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1606821651
transform 1 0 14444 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_128
timestamp 1606821651
transform 1 0 12880 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1606821651
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1606821651
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1606821651
transform 1 0 15180 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1606821651
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2484 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_11
timestamp 1606821651
transform 1 0 2116 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4876 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1606821651
transform 1 0 3680 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1606821651
transform 1 0 3312 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_37
timestamp 1606821651
transform 1 0 4508 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1606821651
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 8464 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 8004 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_71
timestamp 1606821651
transform 1 0 7636 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1606821651
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1606821651
transform 1 0 10304 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1606821651
transform 1 0 9936 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1606821651
transform 1 0 11500 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_109
timestamp 1606821651
transform 1 0 11132 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_117
timestamp 1606821651
transform 1 0 11868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1606821651
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1606821651
transform 1 0 13616 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1606821651
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_145
timestamp 1606821651
transform 1 0 14444 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1606821651
transform 1 0 14812 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1606821651
transform 1 0 15180 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1606821651
transform 1 0 2760 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1606821651
transform 1 0 1564 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_14
timestamp 1606821651
transform 1 0 2392 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4600 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606821651
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_32
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5796 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_47
timestamp 1606821651
transform 1 0 5428 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7636 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1606821651
transform 1 0 7268 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1606821651
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1606821651
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_102
timestamp 1606821651
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1606821651
transform 1 0 10856 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12052 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_115
timestamp 1606821651
transform 1 0 11684 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1606821651
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1606821651
transform 1 0 13248 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_128
timestamp 1606821651
transform 1 0 12880 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1606821651
transform 1 0 14076 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1606821651
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2484 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_11
timestamp 1606821651
transform 1 0 2116 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4876 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1606821651
transform 1 0 3680 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_24
timestamp 1606821651
transform 1 0 3312 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_37
timestamp 1606821651
transform 1 0 4508 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1606821651
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_62
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7360 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1606821651
transform 1 0 9200 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1606821651
transform 1 0 10396 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_84
timestamp 1606821651
transform 1 0 8832 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_97
timestamp 1606821651
transform 1 0 10028 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1606821651
transform 1 0 11592 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_110
timestamp 1606821651
transform 1 0 11224 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1606821651
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  Test_en_E_FTB01
timestamp 1606821651
transform 1 0 13616 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1606821651
transform 1 0 13248 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp 1606821651
transform 1 0 14168 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1606821651
transform 1 0 14536 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_152
timestamp 1606821651
transform 1 0 15088 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_156
timestamp 1606821651
transform 1 0 15456 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1564 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2760 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1606821651
transform 1 0 2392 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4324 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606821651
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_32
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5520 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_44
timestamp 1606821651
transform 1 0 5152 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7360 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_64
timestamp 1606821651
transform 1 0 6992 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 9200 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_84
timestamp 1606821651
transform 1 0 8832 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1606821651
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 1606821651
transform 1 0 10488 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10856 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12052 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_115
timestamp 1606821651
transform 1 0 11684 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606821651
transform 1 0 14444 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_2_S_FTB01
timestamp 1606821651
transform 1 0 13524 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 13248 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_128
timestamp 1606821651
transform 1 0 12880 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1606821651
transform 1 0 14076 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1606821651
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1606821651
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1606821651
transform 1 0 1564 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1606821651
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_14
timestamp 1606821651
transform 1 0 2392 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_17
timestamp 1606821651
transform 1 0 2668 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2760 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3036 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4324 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4876 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_37
timestamp 1606821651
transform 1 0 4508 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1606821651
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6164 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1606821651
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_51
timestamp 1606821651
transform 1 0 5796 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8648 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1606821651
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_78
timestamp 1606821651
transform 1 0 8280 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_71
timestamp 1606821651
transform 1 0 7636 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1606821651
transform 1 0 10488 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 9200 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1606821651
transform 1 0 10120 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_84
timestamp 1606821651
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606821651
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1606821651
transform 1 0 11684 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1606821651
transform 1 0 11500 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_111
timestamp 1606821651
transform 1 0 11316 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1606821651
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_109
timestamp 1606821651
transform 1 0 11132 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_122
timestamp 1606821651
transform 1 0 12328 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_3_S_FTB01
timestamp 1606821651
transform 1 0 13892 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12696 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13892 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 13616 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1606821651
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1606821651
transform 1 0 14444 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1606821651
transform 1 0 13524 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1606821651
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1606821651
transform 1 0 14812 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1606821651
transform 1 0 15180 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2484 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_11
timestamp 1606821651
transform 1 0 2116 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4876 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1606821651
transform 1 0 3680 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_24
timestamp 1606821651
transform 1 0 3312 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_37
timestamp 1606821651
transform 1 0 4508 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1606821651
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8648 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_78
timestamp 1606821651
transform 1 0 8280 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10488 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1606821651
transform 1 0 10120 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1606821651
transform 1 0 11684 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_111
timestamp 1606821651
transform 1 0 11316 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1606821651
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606821651
transform 1 0 13800 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_132
timestamp 1606821651
transform 1 0 13248 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_142
timestamp 1606821651
transform 1 0 14168 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1606821651
transform 1 0 14536 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1606821651
transform 1 0 14812 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1606821651
transform 1 0 2760 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1840 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1606821651
transform 1 0 1748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_14
timestamp 1606821651
transform 1 0 2392 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4416 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606821651
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5612 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_45
timestamp 1606821651
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7452 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_65
timestamp 1606821651
transform 1 0 7084 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1606821651
transform 1 0 8924 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1606821651
transform 1 0 10488 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12052 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10856 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_115
timestamp 1606821651
transform 1 0 11684 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_125
timestamp 1606821651
transform 1 0 12604 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1606821651
transform 1 0 14076 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606821651
transform 1 0 13340 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_137
timestamp 1606821651
transform 1 0 13708 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_144
timestamp 1606821651
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1606821651
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1606821651
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1748 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2668 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1606821651
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_13
timestamp 1606821651
transform 1 0 2300 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4876 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1606821651
transform 1 0 3680 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_23
timestamp 1606821651
transform 1 0 3220 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_27
timestamp 1606821651
transform 1 0 3588 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_37
timestamp 1606821651
transform 1 0 4508 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1606821651
transform 1 0 6348 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8648 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_78
timestamp 1606821651
transform 1 0 8280 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9844 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1606821651
transform 1 0 9476 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_104
timestamp 1606821651
transform 1 0 10672 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1606821651
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1606821651
transform 1 0 11040 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1606821651
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1606821651
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1606821651
transform 1 0 13064 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1606821651
transform 1 0 13708 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1606821651
transform 1 0 14352 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_126
timestamp 1606821651
transform 1 0 12696 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_133
timestamp 1606821651
transform 1 0 13340 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 1606821651
transform 1 0 13984 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp 1606821651
transform 1 0 14628 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1606821651
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2300 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1380 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_9
timestamp 1606821651
transform 1 0 1932 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_19
timestamp 1606821651
transform 1 0 2852 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1606821651
transform 1 0 3220 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4600 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1606821651
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_32
timestamp 1606821651
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 5796 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_47
timestamp 1606821651
transform 1 0 5428 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1606821651
transform 1 0 7636 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_67
timestamp 1606821651
transform 1 0 7268 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1606821651
transform 1 0 8464 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606821651
transform 1 0 8832 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1606821651
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1606821651
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1606821651
transform 1 0 10488 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606821651
transform 1 0 10856 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606821651
transform 1 0 11592 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606821651
transform 1 0 12328 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1606821651
transform 1 0 11224 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_118
timestamp 1606821651
transform 1 0 11960 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1606821651
transform 1 0 13064 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1606821651
transform 1 0 13708 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_126
timestamp 1606821651
transform 1 0 12696 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_133
timestamp 1606821651
transform 1 0 13340 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_140 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 13984 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1606821651
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1606821651
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  clk_2_N_FTB01
timestamp 1606821651
transform 1 0 1472 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1606821651
transform 1 0 2392 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1606821651
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_10
timestamp 1606821651
transform 1 0 2024 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_20
timestamp 1606821651
transform 1 0 2944 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4324 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 3312 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 1606821651
transform 1 0 3864 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_34
timestamp 1606821651
transform 1 0 4232 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1606821651
transform 1 0 5520 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_44
timestamp 1606821651
transform 1 0 5152 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1606821651
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8004 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_71
timestamp 1606821651
transform 1 0 7636 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606821651
transform 1 0 10396 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1606821651
transform 1 0 9200 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_84
timestamp 1606821651
transform 1 0 8832 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1606821651
transform 1 0 10028 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606821651
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1606821651
transform 1 0 11132 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_105
timestamp 1606821651
transform 1 0 10764 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1606821651
transform 1 0 11500 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1606821651
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606821651
transform 1 0 13156 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_127
timestamp 1606821651
transform 1 0 12788 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1606821651
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_147
timestamp 1606821651
transform 1 0 14628 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1606821651
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1606821651
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1606821651
transform 1 0 1472 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  Test_en_W_FTB01
timestamp 1606821651
transform 1 0 1380 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_10
timestamp 1606821651
transform 1 0 2024 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_9
timestamp 1606821651
transform 1 0 1932 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_20
timestamp 1606821651
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 2484 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1606821651
transform 1 0 2760 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1606821651
transform 1 0 2392 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1606821651
transform 1 0 3588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1606821651
transform 1 0 3312 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606821651
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1606821651
transform 1 0 3312 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 4048 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01
timestamp 1606821651
transform 1 0 4048 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1606821651
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_38
timestamp 1606821651
transform 1 0 4600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606821651
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1606821651
transform 1 0 4968 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5612 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1606821651
transform 1 0 6256 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4968 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_51
timestamp 1606821651
transform 1 0 5796 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_55
timestamp 1606821651
transform 1 0 6164 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1606821651
transform 1 0 5244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_58
timestamp 1606821651
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 8648 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6900 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1606821651
transform 1 0 8096 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1606821651
transform 1 0 7452 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_65
timestamp 1606821651
transform 1 0 7084 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_78
timestamp 1606821651
transform 1 0 8280 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_72
timestamp 1606821651
transform 1 0 7728 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1606821651
transform 1 0 8924 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1606821651
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_92
timestamp 1606821651
transform 1 0 9568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_right_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 9292 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606821651
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp 1606821651
transform 1 0 10028 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606821651
transform 1 0 9752 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_98
timestamp 1606821651
transform 1 0 10120 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606821651
transform 1 0 10396 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606821651
transform 1 0 10488 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_106
timestamp 1606821651
transform 1 0 10856 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_113
timestamp 1606821651
transform 1 0 11500 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_105
timestamp 1606821651
transform 1 0 10764 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606821651
transform 1 0 11132 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606821651
transform 1 0 11224 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_114
timestamp 1606821651
transform 1 0 11592 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_121
timestamp 1606821651
transform 1 0 12236 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606821651
transform 1 0 11868 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_122
timestamp 1606821651
transform 1 0 12328 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606821651
transform 1 0 12604 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606821651
transform 1 0 12604 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606821651
transform 1 0 13340 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606821651
transform 1 0 14076 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606821651
transform 1 0 13340 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1606821651
transform 1 0 12972 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_137
timestamp 1606821651
transform 1 0 13708 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_145
timestamp 1606821651
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_129
timestamp 1606821651
transform 1 0 12972 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1606821651
transform 1 0 13708 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 15824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 15824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1606821651
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_149
timestamp 1606821651
transform 1 0 14812 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1606821651
transform 1 0 15456 0 1 16864
box -38 -48 130 592
<< labels >>
rlabel metal3 s 16520 16600 17000 16720 6 Test_en_E_in
port 0 nsew default input
rlabel metal3 s 16520 9936 17000 10056 6 Test_en_E_out
port 1 nsew default tristate
rlabel metal2 s 3146 19520 3202 20000 6 Test_en_N_out
port 2 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 Test_en_S_in
port 3 nsew default input
rlabel metal3 s 0 17280 480 17400 6 Test_en_W_in
port 4 nsew default input
rlabel metal3 s 0 18368 480 18488 6 Test_en_W_out
port 5 nsew default tristate
rlabel metal3 s 0 416 480 536 6 ccff_head
port 6 nsew default input
rlabel metal3 s 16520 3272 17000 3392 6 ccff_tail
port 7 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[0]
port 8 nsew default input
rlabel metal2 s 10322 0 10378 480 6 chany_bottom_in[10]
port 9 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[11]
port 10 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[12]
port 11 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[13]
port 12 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_in[14]
port 13 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[15]
port 14 nsew default input
rlabel metal2 s 12346 0 12402 480 6 chany_bottom_in[16]
port 15 nsew default input
rlabel metal2 s 12622 0 12678 480 6 chany_bottom_in[17]
port 16 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[18]
port 17 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[19]
port 18 nsew default input
rlabel metal2 s 7194 0 7250 480 6 chany_bottom_in[1]
port 19 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[2]
port 20 nsew default input
rlabel metal2 s 7930 0 7986 480 6 chany_bottom_in[3]
port 21 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[4]
port 22 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[5]
port 23 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[6]
port 24 nsew default input
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_in[7]
port 25 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_in[8]
port 26 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[9]
port 27 nsew default input
rlabel metal2 s 110 0 166 480 6 chany_bottom_out[0]
port 28 nsew default tristate
rlabel metal2 s 3514 0 3570 480 6 chany_bottom_out[10]
port 29 nsew default tristate
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_out[11]
port 30 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_out[12]
port 31 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_out[13]
port 32 nsew default tristate
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_out[14]
port 33 nsew default tristate
rlabel metal2 s 5170 0 5226 480 6 chany_bottom_out[15]
port 34 nsew default tristate
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_out[16]
port 35 nsew default tristate
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_out[17]
port 36 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_out[18]
port 37 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[19]
port 38 nsew default tristate
rlabel metal2 s 386 0 442 480 6 chany_bottom_out[1]
port 39 nsew default tristate
rlabel metal2 s 754 0 810 480 6 chany_bottom_out[2]
port 40 nsew default tristate
rlabel metal2 s 1122 0 1178 480 6 chany_bottom_out[3]
port 41 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[4]
port 42 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_out[5]
port 43 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_out[6]
port 44 nsew default tristate
rlabel metal2 s 2410 0 2466 480 6 chany_bottom_out[7]
port 45 nsew default tristate
rlabel metal2 s 2778 0 2834 480 6 chany_bottom_out[8]
port 46 nsew default tristate
rlabel metal2 s 3146 0 3202 480 6 chany_bottom_out[9]
port 47 nsew default tristate
rlabel metal2 s 10322 19520 10378 20000 6 chany_top_in[0]
port 48 nsew default input
rlabel metal2 s 13726 19520 13782 20000 6 chany_top_in[10]
port 49 nsew default input
rlabel metal2 s 14002 19520 14058 20000 6 chany_top_in[11]
port 50 nsew default input
rlabel metal2 s 14370 19520 14426 20000 6 chany_top_in[12]
port 51 nsew default input
rlabel metal2 s 14738 19520 14794 20000 6 chany_top_in[13]
port 52 nsew default input
rlabel metal2 s 15014 19520 15070 20000 6 chany_top_in[14]
port 53 nsew default input
rlabel metal2 s 15382 19520 15438 20000 6 chany_top_in[15]
port 54 nsew default input
rlabel metal2 s 15750 19520 15806 20000 6 chany_top_in[16]
port 55 nsew default input
rlabel metal2 s 16026 19520 16082 20000 6 chany_top_in[17]
port 56 nsew default input
rlabel metal2 s 16394 19520 16450 20000 6 chany_top_in[18]
port 57 nsew default input
rlabel metal2 s 16762 19520 16818 20000 6 chany_top_in[19]
port 58 nsew default input
rlabel metal2 s 10598 19520 10654 20000 6 chany_top_in[1]
port 59 nsew default input
rlabel metal2 s 10966 19520 11022 20000 6 chany_top_in[2]
port 60 nsew default input
rlabel metal2 s 11334 19520 11390 20000 6 chany_top_in[3]
port 61 nsew default input
rlabel metal2 s 11610 19520 11666 20000 6 chany_top_in[4]
port 62 nsew default input
rlabel metal2 s 11978 19520 12034 20000 6 chany_top_in[5]
port 63 nsew default input
rlabel metal2 s 12346 19520 12402 20000 6 chany_top_in[6]
port 64 nsew default input
rlabel metal2 s 12622 19520 12678 20000 6 chany_top_in[7]
port 65 nsew default input
rlabel metal2 s 12990 19520 13046 20000 6 chany_top_in[8]
port 66 nsew default input
rlabel metal2 s 13358 19520 13414 20000 6 chany_top_in[9]
port 67 nsew default input
rlabel metal2 s 3514 19520 3570 20000 6 chany_top_out[0]
port 68 nsew default tristate
rlabel metal2 s 6918 19520 6974 20000 6 chany_top_out[10]
port 69 nsew default tristate
rlabel metal2 s 7194 19520 7250 20000 6 chany_top_out[11]
port 70 nsew default tristate
rlabel metal2 s 7562 19520 7618 20000 6 chany_top_out[12]
port 71 nsew default tristate
rlabel metal2 s 7930 19520 7986 20000 6 chany_top_out[13]
port 72 nsew default tristate
rlabel metal2 s 8206 19520 8262 20000 6 chany_top_out[14]
port 73 nsew default tristate
rlabel metal2 s 8574 19520 8630 20000 6 chany_top_out[15]
port 74 nsew default tristate
rlabel metal2 s 8942 19520 8998 20000 6 chany_top_out[16]
port 75 nsew default tristate
rlabel metal2 s 9218 19520 9274 20000 6 chany_top_out[17]
port 76 nsew default tristate
rlabel metal2 s 9586 19520 9642 20000 6 chany_top_out[18]
port 77 nsew default tristate
rlabel metal2 s 9954 19520 10010 20000 6 chany_top_out[19]
port 78 nsew default tristate
rlabel metal2 s 3790 19520 3846 20000 6 chany_top_out[1]
port 79 nsew default tristate
rlabel metal2 s 4158 19520 4214 20000 6 chany_top_out[2]
port 80 nsew default tristate
rlabel metal2 s 4526 19520 4582 20000 6 chany_top_out[3]
port 81 nsew default tristate
rlabel metal2 s 4802 19520 4858 20000 6 chany_top_out[4]
port 82 nsew default tristate
rlabel metal2 s 5170 19520 5226 20000 6 chany_top_out[5]
port 83 nsew default tristate
rlabel metal2 s 5538 19520 5594 20000 6 chany_top_out[6]
port 84 nsew default tristate
rlabel metal2 s 5814 19520 5870 20000 6 chany_top_out[7]
port 85 nsew default tristate
rlabel metal2 s 6182 19520 6238 20000 6 chany_top_out[8]
port 86 nsew default tristate
rlabel metal2 s 6550 19520 6606 20000 6 chany_top_out[9]
port 87 nsew default tristate
rlabel metal2 s 110 19520 166 20000 6 clk_2_N_in
port 88 nsew default input
rlabel metal2 s 1398 19520 1454 20000 6 clk_2_N_out
port 89 nsew default tristate
rlabel metal2 s 14002 0 14058 480 6 clk_2_S_in
port 90 nsew default input
rlabel metal2 s 15382 0 15438 480 6 clk_2_S_out
port 91 nsew default tristate
rlabel metal2 s 386 19520 442 20000 6 clk_3_N_in
port 92 nsew default input
rlabel metal2 s 1766 19520 1822 20000 6 clk_3_N_out
port 93 nsew default tristate
rlabel metal2 s 14370 0 14426 480 6 clk_3_S_in
port 94 nsew default input
rlabel metal2 s 15750 0 15806 480 6 clk_3_S_out
port 95 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 left_grid_pin_16_
port 96 nsew default tristate
rlabel metal3 s 0 2320 480 2440 6 left_grid_pin_17_
port 97 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 left_grid_pin_18_
port 98 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 left_grid_pin_19_
port 99 nsew default tristate
rlabel metal3 s 0 5312 480 5432 6 left_grid_pin_20_
port 100 nsew default tristate
rlabel metal3 s 0 6400 480 6520 6 left_grid_pin_21_
port 101 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 left_grid_pin_22_
port 102 nsew default tristate
rlabel metal3 s 0 8304 480 8424 6 left_grid_pin_23_
port 103 nsew default tristate
rlabel metal3 s 0 9392 480 9512 6 left_grid_pin_24_
port 104 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 left_grid_pin_25_
port 105 nsew default tristate
rlabel metal3 s 0 11296 480 11416 6 left_grid_pin_26_
port 106 nsew default tristate
rlabel metal3 s 0 12384 480 12504 6 left_grid_pin_27_
port 107 nsew default tristate
rlabel metal3 s 0 13336 480 13456 6 left_grid_pin_28_
port 108 nsew default tristate
rlabel metal3 s 0 14288 480 14408 6 left_grid_pin_29_
port 109 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 left_grid_pin_30_
port 110 nsew default tristate
rlabel metal3 s 0 16328 480 16448 6 left_grid_pin_31_
port 111 nsew default tristate
rlabel metal2 s 2134 19520 2190 20000 6 prog_clk_0_N_out
port 112 nsew default tristate
rlabel metal2 s 16026 0 16082 480 6 prog_clk_0_S_out
port 113 nsew default tristate
rlabel metal3 s 0 19320 480 19440 6 prog_clk_0_W_in
port 114 nsew default input
rlabel metal2 s 754 19520 810 20000 6 prog_clk_2_N_in
port 115 nsew default input
rlabel metal2 s 2410 19520 2466 20000 6 prog_clk_2_N_out
port 116 nsew default tristate
rlabel metal2 s 14738 0 14794 480 6 prog_clk_2_S_in
port 117 nsew default input
rlabel metal2 s 16394 0 16450 480 6 prog_clk_2_S_out
port 118 nsew default tristate
rlabel metal2 s 1122 19520 1178 20000 6 prog_clk_3_N_in
port 119 nsew default input
rlabel metal2 s 2778 19520 2834 20000 6 prog_clk_3_N_out
port 120 nsew default tristate
rlabel metal2 s 15014 0 15070 480 6 prog_clk_3_S_in
port 121 nsew default input
rlabel metal2 s 16762 0 16818 480 6 prog_clk_3_S_out
port 122 nsew default tristate
rlabel metal4 s 3409 2128 3729 17456 6 VPWR
port 123 nsew default input
rlabel metal4 s 5875 2128 6195 17456 6 VGND
port 124 nsew default input
<< properties >>
string FIXED_BBOX 0 0 17000 20000
<< end >>
